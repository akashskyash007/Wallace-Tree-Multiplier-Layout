magic
tech scmos
timestamp 1199203224
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 68
rect 36 63 38 68
rect 46 59 48 64
rect 53 59 55 64
rect 9 39 11 43
rect 19 39 21 43
rect 9 37 21 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 29 34 31 43
rect 36 40 38 43
rect 46 40 48 43
rect 36 38 48 40
rect 53 40 55 43
rect 53 38 62 40
rect 38 36 48 38
rect 38 34 42 36
rect 44 34 48 36
rect 56 36 58 38
rect 60 36 62 38
rect 56 34 62 36
rect 9 30 11 33
rect 28 32 34 34
rect 28 30 30 32
rect 32 30 34 32
rect 28 28 34 30
rect 38 32 48 34
rect 28 25 30 28
rect 38 25 40 32
rect 28 10 30 15
rect 38 10 40 15
rect 9 6 11 10
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 25 26 30
rect 11 22 28 25
rect 11 20 14 22
rect 16 20 28 22
rect 11 15 28 20
rect 30 23 38 25
rect 30 21 33 23
rect 35 21 38 23
rect 30 15 38 21
rect 40 19 48 25
rect 40 17 43 19
rect 45 17 48 19
rect 40 15 48 17
rect 11 14 26 15
rect 11 12 14 14
rect 16 12 22 14
rect 24 12 26 14
rect 11 10 26 12
<< pdif >>
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 43 9 52
rect 11 54 19 63
rect 11 52 14 54
rect 16 52 19 54
rect 11 47 19 52
rect 11 45 14 47
rect 16 45 19 47
rect 11 43 19 45
rect 21 61 29 63
rect 21 59 24 61
rect 26 59 29 61
rect 21 43 29 59
rect 31 43 36 63
rect 38 59 43 63
rect 38 53 46 59
rect 38 51 41 53
rect 43 51 46 53
rect 38 43 46 51
rect 48 43 53 59
rect 55 57 62 59
rect 55 55 58 57
rect 60 55 62 57
rect 55 43 62 55
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 13 54 17 56
rect 13 52 14 54
rect 16 52 17 54
rect 13 47 17 52
rect 2 45 14 47
rect 16 45 17 47
rect 2 42 17 45
rect 2 30 6 42
rect 58 46 62 47
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 29 42 62 46
rect 29 32 33 42
rect 29 30 30 32
rect 32 30 33 32
rect 29 28 33 30
rect 41 36 47 38
rect 41 34 42 36
rect 44 34 47 36
rect 58 38 62 42
rect 60 36 62 38
rect 41 31 47 34
rect 58 33 62 36
rect 41 25 54 31
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 10 11 30
rect 28 15 30 25
rect 38 15 40 25
<< pmos >>
rect 9 43 11 63
rect 19 43 21 63
rect 29 43 31 63
rect 36 43 38 63
rect 46 43 48 59
rect 53 43 55 59
<< polyct0 >>
rect 17 35 19 37
<< polyct1 >>
rect 42 34 44 36
rect 58 36 60 38
rect 30 30 32 32
<< ndifct0 >>
rect 14 20 16 22
rect 33 21 35 23
rect 43 17 45 19
rect 14 12 16 14
rect 22 12 24 14
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 59 6 61
rect 4 52 6 54
rect 24 59 26 61
rect 41 51 43 53
rect 58 55 60 57
<< pdifct1 >>
rect 14 52 16 54
rect 14 45 16 47
<< alu0 >>
rect 2 61 8 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 54 8 59
rect 22 61 28 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 57 57 61 68
rect 2 52 4 54
rect 6 52 8 54
rect 2 51 8 52
rect 57 55 58 57
rect 60 55 61 57
rect 21 53 45 54
rect 57 53 61 55
rect 21 51 41 53
rect 43 51 45 53
rect 21 50 45 51
rect 21 38 25 50
rect 15 37 25 38
rect 15 35 17 37
rect 19 35 25 37
rect 15 34 25 35
rect 21 24 25 34
rect 56 35 58 42
rect 13 22 17 24
rect 13 20 14 22
rect 16 20 17 22
rect 21 23 37 24
rect 21 21 33 23
rect 35 21 37 23
rect 21 20 37 21
rect 13 14 17 20
rect 42 19 46 21
rect 42 17 43 19
rect 45 17 46 19
rect 13 12 14 14
rect 16 12 17 14
rect 21 14 25 16
rect 21 12 22 14
rect 24 12 25 14
rect 42 12 46 17
<< labels >>
rlabel alu0 20 36 20 36 6 zn
rlabel alu0 29 22 29 22 6 zn
rlabel alu0 33 52 33 52 6 zn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 32 44 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 b
rlabel alu1 60 40 60 40 6 a
rlabel alu1 52 44 52 44 6 a
<< end >>
