magic
tech scmos
timestamp 1199203040
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 26 70 28 74
rect 12 39 14 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 33 21 42
rect 26 39 28 42
rect 26 37 38 39
rect 29 35 34 37
rect 36 35 38 37
rect 29 33 38 35
rect 9 29 11 33
rect 19 31 25 33
rect 19 29 21 31
rect 23 29 25 31
rect 19 27 25 29
rect 19 24 21 27
rect 29 24 31 33
rect 9 15 11 19
rect 19 9 21 14
rect 29 9 31 14
<< ndif >>
rect 4 25 9 29
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 24 17 29
rect 11 19 19 24
rect 13 14 19 19
rect 21 21 29 24
rect 21 19 24 21
rect 26 19 29 21
rect 21 14 29 19
rect 31 18 38 24
rect 31 16 34 18
rect 36 16 38 18
rect 31 14 38 16
rect 13 13 17 14
rect 11 11 17 13
rect 11 9 13 11
rect 15 9 17 11
rect 11 7 17 9
<< pdif >>
rect 7 63 12 70
rect 5 61 12 63
rect 5 59 7 61
rect 9 59 12 61
rect 5 54 12 59
rect 5 52 7 54
rect 9 52 12 54
rect 5 50 12 52
rect 7 42 12 50
rect 14 42 19 70
rect 21 42 26 70
rect 28 68 38 70
rect 28 66 34 68
rect 36 66 38 68
rect 28 61 38 66
rect 28 59 34 61
rect 36 59 38 61
rect 28 42 38 59
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 5 61 11 62
rect 5 59 7 61
rect 9 59 11 61
rect 5 55 11 59
rect 2 54 11 55
rect 2 52 7 54
rect 9 52 11 54
rect 2 51 11 52
rect 2 25 6 51
rect 18 47 22 55
rect 34 47 38 55
rect 10 43 22 47
rect 10 37 14 43
rect 26 41 38 47
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 18 34 22 39
rect 18 31 24 34
rect 18 30 21 31
rect 20 29 21 30
rect 23 30 24 31
rect 23 29 31 30
rect 20 26 31 29
rect 2 23 7 25
rect 2 21 4 23
rect 6 22 7 23
rect 6 21 28 22
rect 2 19 24 21
rect 26 19 28 21
rect 2 18 28 19
rect -2 11 42 12
rect -2 9 13 11
rect 15 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 19 11 29
rect 19 14 21 24
rect 29 14 31 24
<< pmos >>
rect 12 42 14 70
rect 19 42 21 70
rect 26 42 28 70
<< polyct0 >>
rect 34 35 36 37
<< polyct1 >>
rect 11 35 13 37
rect 21 29 23 31
<< ndifct0 >>
rect 34 16 36 18
<< ndifct1 >>
rect 4 21 6 23
rect 24 19 26 21
rect 13 9 15 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 34 66 36 68
rect 34 59 36 61
<< pdifct1 >>
rect 7 59 9 61
rect 7 52 9 54
<< alu0 >>
rect 32 66 34 68
rect 36 66 38 68
rect 32 61 38 66
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 33 37 37 41
rect 33 35 34 37
rect 36 35 37 37
rect 33 33 37 35
rect 33 18 37 20
rect 33 16 34 18
rect 36 16 37 18
rect 33 12 37 16
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 40 12 40 6 c
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 36 20 36 6 b
rlabel alu1 28 28 28 28 6 b
rlabel alu1 28 44 28 44 6 a
rlabel alu1 20 52 20 52 6 c
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 48 36 48 6 a
<< end >>
