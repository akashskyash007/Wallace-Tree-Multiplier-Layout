magic
tech scmos
timestamp 1199203211
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 22 70 24 74
rect 29 70 31 74
rect 9 60 11 65
rect 9 39 11 42
rect 22 39 24 49
rect 29 46 31 49
rect 29 44 35 46
rect 29 42 31 44
rect 33 42 35 44
rect 29 40 35 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 40
rect 9 16 11 21
rect 19 19 21 24
rect 29 19 31 24
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 21 9 24
rect 11 24 19 30
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 24 29 26
rect 31 24 38 30
rect 11 21 17 24
rect 13 17 17 21
rect 33 17 38 24
rect 13 15 19 17
rect 13 13 15 15
rect 17 13 19 15
rect 13 11 19 13
rect 32 15 38 17
rect 32 13 34 15
rect 36 13 38 15
rect 32 11 38 13
<< pdif >>
rect 13 68 22 70
rect 13 66 15 68
rect 17 66 22 68
rect 13 60 22 66
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 51 9 56
rect 2 49 4 51
rect 6 49 9 51
rect 2 47 9 49
rect 4 42 9 47
rect 11 49 22 60
rect 24 49 29 70
rect 31 63 36 70
rect 31 61 38 63
rect 31 59 34 61
rect 36 59 38 61
rect 31 57 38 59
rect 31 49 36 57
rect 11 42 19 49
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 62 6 63
rect 2 58 15 62
rect 2 56 4 58
rect 2 51 6 56
rect 2 49 4 51
rect 2 30 6 49
rect 34 46 38 55
rect 17 44 38 46
rect 17 42 31 44
rect 33 42 38 44
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 24 7 26
rect 17 37 38 38
rect 17 35 21 37
rect 23 35 38 37
rect 17 34 38 35
rect 34 25 38 34
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 21 11 30
rect 19 24 21 30
rect 29 24 31 30
<< pmos >>
rect 9 42 11 60
rect 22 49 24 70
rect 29 49 31 70
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 42 33 44
rect 21 35 23 37
<< ndifct0 >>
rect 24 26 26 28
rect 15 13 17 15
rect 34 13 36 15
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 15 66 17 68
rect 34 59 36 61
<< pdifct1 >>
rect 4 56 6 58
rect 4 49 6 51
<< alu0 >>
rect 13 66 15 68
rect 17 66 19 68
rect 13 65 19 66
rect 21 61 38 62
rect 21 59 34 61
rect 36 59 38 61
rect 21 58 38 59
rect 6 47 7 58
rect 21 54 25 58
rect 10 50 25 54
rect 10 37 14 50
rect 29 41 35 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 10 28 28 29
rect 10 26 24 28
rect 26 26 28 28
rect 10 25 28 26
rect 13 15 19 16
rect 13 13 15 15
rect 17 13 19 15
rect 13 12 19 13
rect 32 15 38 16
rect 32 13 34 15
rect 36 13 38 15
rect 32 12 38 13
<< labels >>
rlabel alu0 12 39 12 39 6 zn
rlabel alu0 19 27 19 27 6 zn
rlabel alu0 29 60 29 60 6 zn
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 36 28 36 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 44 20 44 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 52 36 52 6 b
<< end >>
