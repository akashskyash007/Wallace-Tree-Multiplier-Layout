magic
tech scmos
timestamp 1199202386
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 10 62 12 67
rect 20 54 22 59
rect 10 35 12 38
rect 20 35 22 38
rect 9 33 23 35
rect 9 31 19 33
rect 21 31 23 33
rect 9 29 23 31
rect 9 26 11 29
rect 9 6 11 11
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 11 9 13
rect 11 23 19 26
rect 11 21 14 23
rect 16 21 19 23
rect 11 15 19 21
rect 11 13 14 15
rect 16 13 19 15
rect 11 11 19 13
<< pdif >>
rect 2 60 10 62
rect 2 58 5 60
rect 7 58 10 60
rect 2 52 10 58
rect 2 50 5 52
rect 7 50 10 52
rect 2 38 10 50
rect 12 54 17 62
rect 12 49 20 54
rect 12 47 15 49
rect 17 47 20 49
rect 12 42 20 47
rect 12 40 15 42
rect 17 40 20 42
rect 12 38 20 40
rect 22 52 30 54
rect 22 50 25 52
rect 27 50 30 52
rect 22 38 30 50
<< alu1 >>
rect -2 67 34 72
rect -2 65 24 67
rect 26 65 34 67
rect -2 64 34 65
rect 2 37 14 43
rect 2 26 6 37
rect 26 35 30 43
rect 18 33 30 35
rect 18 31 19 33
rect 21 31 30 33
rect 18 29 30 31
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 17 7 22
rect 2 15 4 17
rect 6 15 7 17
rect 2 13 7 15
rect -2 7 34 8
rect -2 5 25 7
rect 27 5 34 7
rect -2 0 34 5
<< ptie >>
rect 23 7 29 24
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< ntie >>
rect 22 67 28 69
rect 22 65 24 67
rect 26 65 28 67
rect 22 62 28 65
<< nmos >>
rect 9 11 11 26
<< pmos >>
rect 10 38 12 62
rect 20 38 22 54
<< polyct1 >>
rect 19 31 21 33
<< ndifct0 >>
rect 14 21 16 23
rect 14 13 16 15
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
<< ntiect1 >>
rect 24 65 26 67
<< ptiect1 >>
rect 25 5 27 7
<< pdifct0 >>
rect 5 58 7 60
rect 5 50 7 52
rect 15 47 17 49
rect 15 40 17 42
rect 25 50 27 52
<< alu0 >>
rect 4 60 8 64
rect 4 58 5 60
rect 7 58 8 60
rect 4 52 8 58
rect 4 50 5 52
rect 7 50 8 52
rect 24 52 28 64
rect 24 50 25 52
rect 27 50 28 52
rect 4 48 8 50
rect 13 49 19 50
rect 13 47 15 49
rect 17 47 19 49
rect 24 48 28 50
rect 13 43 19 47
rect 14 42 19 43
rect 14 40 15 42
rect 17 40 19 42
rect 14 39 19 40
rect 13 23 17 25
rect 13 21 14 23
rect 16 21 17 23
rect 13 15 17 21
rect 13 13 14 15
rect 16 13 17 15
rect 13 8 17 13
<< labels >>
rlabel alu1 4 28 4 28 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 12 40 12 40 6 z
rlabel alu1 16 68 16 68 6 vdd
rlabel polyct1 20 32 20 32 6 a
rlabel alu1 28 36 28 36 6 a
<< end >>
