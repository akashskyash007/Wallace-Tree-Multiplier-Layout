magic
tech scmos
timestamp 1199202935
<< ab >>
rect 0 0 152 72
<< nwell >>
rect -5 32 157 77
<< pwell >>
rect -5 -5 157 32
<< poly >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 50 66 52 70
rect 60 66 62 70
rect 67 66 69 70
rect 77 66 79 70
rect 84 66 86 70
rect 94 66 96 70
rect 101 66 103 70
rect 111 66 113 70
rect 118 66 120 70
rect 128 57 130 61
rect 135 57 137 61
rect 9 29 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 33 35 35 38
rect 43 35 45 38
rect 50 35 52 38
rect 60 35 62 38
rect 16 33 29 35
rect 33 33 45 35
rect 23 31 25 33
rect 27 31 29 33
rect 23 29 29 31
rect 9 27 15 29
rect 9 25 11 27
rect 13 25 15 27
rect 27 26 29 29
rect 37 31 39 33
rect 41 32 45 33
rect 49 33 62 35
rect 67 35 69 38
rect 77 35 79 38
rect 67 33 79 35
rect 41 31 43 32
rect 37 29 43 31
rect 49 31 51 33
rect 53 31 56 33
rect 49 29 56 31
rect 67 31 75 33
rect 77 31 79 33
rect 84 35 86 38
rect 94 35 96 38
rect 84 33 96 35
rect 84 32 91 33
rect 67 29 79 31
rect 86 31 91 32
rect 93 32 96 33
rect 93 31 95 32
rect 86 29 95 31
rect 37 26 39 29
rect 9 23 15 25
rect 54 24 56 29
rect 64 27 69 29
rect 64 24 66 27
rect 76 26 78 29
rect 86 26 88 29
rect 101 27 103 38
rect 111 27 113 38
rect 118 35 120 38
rect 128 35 130 38
rect 118 33 130 35
rect 118 31 120 33
rect 122 31 124 33
rect 118 29 124 31
rect 135 27 137 38
rect 101 25 113 27
rect 129 25 137 27
rect 104 23 106 25
rect 108 23 110 25
rect 104 21 110 23
rect 129 23 131 25
rect 133 23 137 25
rect 129 21 137 23
rect 27 2 29 6
rect 37 2 39 6
rect 54 2 56 6
rect 64 2 66 6
rect 76 2 78 6
rect 86 2 88 6
<< ndif >>
rect 19 10 27 26
rect 19 8 22 10
rect 24 8 27 10
rect 19 6 27 8
rect 29 17 37 26
rect 29 15 32 17
rect 34 15 37 17
rect 29 6 37 15
rect 39 24 51 26
rect 71 24 76 26
rect 39 10 54 24
rect 39 8 45 10
rect 47 8 54 10
rect 39 6 54 8
rect 56 17 64 24
rect 56 15 59 17
rect 61 15 64 17
rect 56 6 64 15
rect 66 10 76 24
rect 66 8 70 10
rect 72 8 76 10
rect 66 6 76 8
rect 78 17 86 26
rect 78 15 81 17
rect 83 15 86 17
rect 78 6 86 15
rect 88 17 96 26
rect 88 15 91 17
rect 93 15 96 17
rect 88 10 96 15
rect 88 8 91 10
rect 93 8 96 10
rect 88 6 96 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 38 16 66
rect 18 57 26 66
rect 18 55 21 57
rect 23 55 26 57
rect 18 49 26 55
rect 18 47 21 49
rect 23 47 26 49
rect 18 38 26 47
rect 28 38 33 66
rect 35 64 43 66
rect 35 62 38 64
rect 40 62 43 64
rect 35 57 43 62
rect 35 55 38 57
rect 40 55 43 57
rect 35 38 43 55
rect 45 38 50 66
rect 52 56 60 66
rect 52 54 55 56
rect 57 54 60 56
rect 52 49 60 54
rect 52 47 55 49
rect 57 47 60 49
rect 52 38 60 47
rect 62 38 67 66
rect 69 64 77 66
rect 69 62 72 64
rect 74 62 77 64
rect 69 57 77 62
rect 69 55 72 57
rect 74 55 77 57
rect 69 38 77 55
rect 79 38 84 66
rect 86 57 94 66
rect 86 55 89 57
rect 91 55 94 57
rect 86 49 94 55
rect 86 47 89 49
rect 91 47 94 49
rect 86 38 94 47
rect 96 38 101 66
rect 103 64 111 66
rect 103 62 106 64
rect 108 62 111 64
rect 103 57 111 62
rect 103 55 106 57
rect 108 55 111 57
rect 103 38 111 55
rect 113 38 118 66
rect 120 57 125 66
rect 120 49 128 57
rect 120 47 123 49
rect 125 47 128 49
rect 120 42 128 47
rect 120 40 123 42
rect 125 40 128 42
rect 120 38 128 40
rect 130 38 135 57
rect 137 55 145 57
rect 137 53 140 55
rect 142 53 145 55
rect 137 48 145 53
rect 137 46 140 48
rect 142 46 145 48
rect 137 38 145 46
<< alu1 >>
rect -2 67 154 72
rect -2 65 132 67
rect 134 65 141 67
rect 143 65 154 67
rect -2 64 154 65
rect 18 57 24 59
rect 18 55 21 57
rect 23 55 24 57
rect 18 50 24 55
rect 88 57 94 59
rect 88 55 89 57
rect 91 55 94 57
rect 88 50 94 55
rect 2 49 127 50
rect 2 47 21 49
rect 23 47 55 49
rect 57 47 89 49
rect 91 47 123 49
rect 125 47 127 49
rect 2 46 127 47
rect 2 18 6 46
rect 121 42 127 46
rect 25 38 95 42
rect 121 40 123 42
rect 125 40 127 42
rect 121 38 127 40
rect 25 34 31 38
rect 23 33 31 34
rect 23 31 25 33
rect 27 31 31 33
rect 23 30 31 31
rect 10 27 14 29
rect 10 25 11 27
rect 13 26 14 27
rect 49 33 55 38
rect 89 34 95 38
rect 49 31 51 33
rect 53 31 55 33
rect 49 30 55 31
rect 73 33 79 34
rect 73 31 75 33
rect 77 31 79 33
rect 73 26 79 31
rect 89 33 127 34
rect 89 31 91 33
rect 93 31 120 33
rect 122 31 127 33
rect 89 30 127 31
rect 13 25 135 26
rect 10 23 106 25
rect 108 23 131 25
rect 133 23 135 25
rect 10 22 135 23
rect 2 17 85 18
rect 2 15 32 17
rect 34 15 59 17
rect 61 15 81 17
rect 83 15 85 17
rect 2 14 85 15
rect -2 7 154 8
rect -2 5 5 7
rect 7 5 102 7
rect 104 5 133 7
rect 135 5 141 7
rect 143 5 154 7
rect -2 0 154 5
<< ptie >>
rect 3 7 9 20
rect 3 5 5 7
rect 7 5 9 7
rect 100 7 106 19
rect 3 3 9 5
rect 100 5 102 7
rect 104 5 106 7
rect 100 3 106 5
rect 131 7 145 18
rect 131 5 133 7
rect 135 5 141 7
rect 143 5 145 7
rect 131 3 145 5
<< ntie >>
rect 130 67 145 69
rect 130 65 132 67
rect 134 65 141 67
rect 143 65 145 67
rect 130 63 145 65
<< nmos >>
rect 27 6 29 26
rect 37 6 39 26
rect 54 6 56 24
rect 64 6 66 24
rect 76 6 78 26
rect 86 6 88 26
<< pmos >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 38 45 66
rect 50 38 52 66
rect 60 38 62 66
rect 67 38 69 66
rect 77 38 79 66
rect 84 38 86 66
rect 94 38 96 66
rect 101 38 103 66
rect 111 38 113 66
rect 118 38 120 66
rect 128 38 130 57
rect 135 38 137 57
<< polyct0 >>
rect 39 31 41 33
<< polyct1 >>
rect 25 31 27 33
rect 11 25 13 27
rect 51 31 53 33
rect 75 31 77 33
rect 91 31 93 33
rect 120 31 122 33
rect 106 23 108 25
rect 131 23 133 25
<< ndifct0 >>
rect 22 8 24 10
rect 45 8 47 10
rect 70 8 72 10
rect 91 15 93 17
rect 91 8 93 10
<< ndifct1 >>
rect 32 15 34 17
rect 59 15 61 17
rect 81 15 83 17
<< ntiect1 >>
rect 132 65 134 67
rect 141 65 143 67
<< ptiect1 >>
rect 5 5 7 7
rect 102 5 104 7
rect 133 5 135 7
rect 141 5 143 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 38 62 40 64
rect 38 55 40 57
rect 55 54 57 56
rect 72 62 74 64
rect 72 55 74 57
rect 106 62 108 64
rect 106 55 108 57
rect 140 53 142 55
rect 140 46 142 48
<< pdifct1 >>
rect 21 55 23 57
rect 21 47 23 49
rect 55 47 57 49
rect 89 55 91 57
rect 89 47 91 49
rect 123 47 125 49
rect 123 40 125 42
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 36 62 38 64
rect 40 62 42 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 36 57 42 62
rect 70 62 72 64
rect 74 62 76 64
rect 36 55 38 57
rect 40 55 42 57
rect 36 54 42 55
rect 54 56 58 58
rect 54 54 55 56
rect 57 54 58 56
rect 70 57 76 62
rect 104 62 106 64
rect 108 62 110 64
rect 70 55 72 57
rect 74 55 76 57
rect 70 54 76 55
rect 54 50 58 54
rect 104 57 110 62
rect 104 55 106 57
rect 108 55 110 57
rect 104 54 110 55
rect 138 55 144 64
rect 138 53 140 55
rect 142 53 144 55
rect 138 48 144 53
rect 138 46 140 48
rect 142 46 144 48
rect 138 45 144 46
rect 37 33 43 34
rect 37 31 39 33
rect 41 31 43 33
rect 37 26 43 31
rect 89 17 95 18
rect 89 15 91 17
rect 93 15 95 17
rect 20 10 26 11
rect 20 8 22 10
rect 24 8 26 10
rect 43 10 49 11
rect 43 8 45 10
rect 47 8 49 10
rect 68 10 74 11
rect 68 8 70 10
rect 72 8 74 10
rect 89 10 95 15
rect 89 8 91 10
rect 93 8 95 10
<< labels >>
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 24 20 24 6 a
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 28 24 28 24 6 a
rlabel alu1 52 24 52 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 36 24 36 24 6 a
rlabel alu1 28 32 28 32 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 52 36 52 36 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 76 4 76 4 6 vss
rlabel alu1 76 16 76 16 6 z
rlabel alu1 68 16 68 16 6 z
rlabel ndifct1 60 16 60 16 6 z
rlabel alu1 60 24 60 24 6 a
rlabel alu1 84 24 84 24 6 a
rlabel alu1 68 24 68 24 6 a
rlabel alu1 76 28 76 28 6 a
rlabel alu1 60 40 60 40 6 b
rlabel alu1 84 40 84 40 6 b
rlabel alu1 76 40 76 40 6 b
rlabel alu1 68 40 68 40 6 b
rlabel alu1 60 48 60 48 6 z
rlabel alu1 84 48 84 48 6 z
rlabel alu1 76 48 76 48 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 76 68 76 68 6 vdd
rlabel alu1 92 24 92 24 6 a
rlabel alu1 116 24 116 24 6 a
rlabel alu1 108 24 108 24 6 a
rlabel alu1 100 24 100 24 6 a
rlabel alu1 116 32 116 32 6 b
rlabel alu1 108 32 108 32 6 b
rlabel alu1 100 32 100 32 6 b
rlabel alu1 92 36 92 36 6 b
rlabel alu1 92 52 92 52 6 z
rlabel alu1 116 48 116 48 6 z
rlabel alu1 108 48 108 48 6 z
rlabel alu1 100 48 100 48 6 z
rlabel alu1 124 24 124 24 6 a
rlabel polyct1 132 24 132 24 6 a
rlabel alu1 124 32 124 32 6 b
rlabel alu1 124 44 124 44 6 z
<< end >>
