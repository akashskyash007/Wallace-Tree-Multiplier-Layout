magic
tech scmos
timestamp 1199202138
<< ab >>
rect 0 0 200 72
<< nwell >>
rect -5 32 205 77
<< pwell >>
rect -5 -5 205 32
<< poly >>
rect 21 66 23 70
rect 31 66 33 70
rect 41 66 43 70
rect 51 66 53 70
rect 61 66 63 70
rect 71 66 73 70
rect 81 66 83 70
rect 91 66 93 70
rect 101 66 103 70
rect 108 66 110 70
rect 121 66 123 70
rect 128 66 130 70
rect 138 66 140 70
rect 145 66 147 70
rect 157 66 159 70
rect 167 66 169 70
rect 177 66 179 70
rect 10 46 12 51
rect 10 35 12 38
rect 21 35 23 38
rect 31 35 33 38
rect 10 33 33 35
rect 10 31 12 33
rect 14 31 19 33
rect 21 31 23 33
rect 10 29 23 31
rect 21 26 23 29
rect 31 26 33 33
rect 41 35 43 38
rect 51 35 53 38
rect 41 33 54 35
rect 41 31 43 33
rect 45 31 50 33
rect 52 31 54 33
rect 61 31 63 38
rect 41 29 63 31
rect 41 26 43 29
rect 51 26 53 29
rect 61 26 63 29
rect 71 35 73 38
rect 81 35 83 38
rect 91 35 93 38
rect 101 35 103 38
rect 71 33 93 35
rect 71 31 73 33
rect 75 31 83 33
rect 71 29 83 31
rect 71 26 73 29
rect 81 26 83 29
rect 91 26 93 33
rect 97 33 103 35
rect 97 31 99 33
rect 101 31 103 33
rect 97 29 103 31
rect 101 26 103 29
rect 108 35 110 38
rect 121 35 123 38
rect 108 33 123 35
rect 108 31 115 33
rect 117 31 123 33
rect 108 29 123 31
rect 108 26 110 29
rect 121 26 123 29
rect 128 35 130 38
rect 138 35 140 38
rect 128 33 140 35
rect 128 31 130 33
rect 132 31 140 33
rect 128 29 140 31
rect 128 26 130 29
rect 138 26 140 29
rect 145 35 147 38
rect 157 35 159 38
rect 167 35 169 38
rect 177 35 179 38
rect 145 33 179 35
rect 145 31 147 33
rect 149 31 160 33
rect 145 29 160 31
rect 145 26 147 29
rect 158 26 160 29
rect 168 26 170 33
rect 21 5 23 10
rect 31 5 33 10
rect 41 7 43 12
rect 51 7 53 12
rect 61 4 63 12
rect 71 8 73 12
rect 81 8 83 12
rect 91 8 93 12
rect 101 4 103 12
rect 108 7 110 12
rect 121 7 123 12
rect 128 7 130 12
rect 138 7 140 12
rect 145 7 147 12
rect 61 2 103 4
rect 158 2 160 6
rect 168 2 170 6
<< ndif >>
rect 14 23 21 26
rect 14 21 16 23
rect 18 21 21 23
rect 14 16 21 21
rect 14 14 16 16
rect 18 14 21 16
rect 14 10 21 14
rect 23 24 31 26
rect 23 22 26 24
rect 28 22 31 24
rect 23 17 31 22
rect 23 15 26 17
rect 28 15 31 17
rect 23 10 31 15
rect 33 23 41 26
rect 33 21 36 23
rect 38 21 41 23
rect 33 16 41 21
rect 33 14 36 16
rect 38 14 41 16
rect 33 12 41 14
rect 43 24 51 26
rect 43 22 46 24
rect 48 22 51 24
rect 43 17 51 22
rect 43 15 46 17
rect 48 15 51 17
rect 43 12 51 15
rect 53 16 61 26
rect 53 14 56 16
rect 58 14 61 16
rect 53 12 61 14
rect 63 24 71 26
rect 63 22 66 24
rect 68 22 71 24
rect 63 17 71 22
rect 63 15 66 17
rect 68 15 71 17
rect 63 12 71 15
rect 73 24 81 26
rect 73 22 76 24
rect 78 22 81 24
rect 73 12 81 22
rect 83 17 91 26
rect 83 15 86 17
rect 88 15 91 17
rect 83 12 91 15
rect 93 24 101 26
rect 93 22 96 24
rect 98 22 101 24
rect 93 12 101 22
rect 103 12 108 26
rect 110 12 121 26
rect 123 12 128 26
rect 130 24 138 26
rect 130 22 133 24
rect 135 22 138 24
rect 130 12 138 22
rect 140 12 145 26
rect 147 12 158 26
rect 33 10 39 12
rect 112 7 119 12
rect 149 10 158 12
rect 149 8 151 10
rect 153 8 158 10
rect 112 5 114 7
rect 116 5 119 7
rect 149 6 158 8
rect 160 24 168 26
rect 160 22 163 24
rect 165 22 168 24
rect 160 17 168 22
rect 160 15 163 17
rect 165 15 168 17
rect 160 6 168 15
rect 170 18 178 26
rect 170 16 173 18
rect 175 16 178 18
rect 170 10 178 16
rect 170 8 173 10
rect 175 8 178 10
rect 170 6 178 8
rect 112 3 119 5
<< pdif >>
rect 14 64 21 66
rect 14 62 16 64
rect 18 62 21 64
rect 14 57 21 62
rect 14 55 16 57
rect 18 55 21 57
rect 14 50 21 55
rect 14 48 16 50
rect 18 48 21 50
rect 14 46 21 48
rect 5 44 10 46
rect 3 42 10 44
rect 3 40 5 42
rect 7 40 10 42
rect 3 38 10 40
rect 12 38 21 46
rect 23 49 31 66
rect 23 47 26 49
rect 28 47 31 49
rect 23 42 31 47
rect 23 40 26 42
rect 28 40 31 42
rect 23 38 31 40
rect 33 64 41 66
rect 33 62 36 64
rect 38 62 41 64
rect 33 57 41 62
rect 33 55 36 57
rect 38 55 41 57
rect 33 50 41 55
rect 33 48 36 50
rect 38 48 41 50
rect 33 38 41 48
rect 43 57 51 66
rect 43 55 46 57
rect 48 55 51 57
rect 43 50 51 55
rect 43 48 46 50
rect 48 48 51 50
rect 43 38 51 48
rect 53 64 61 66
rect 53 62 56 64
rect 58 62 61 64
rect 53 57 61 62
rect 53 55 56 57
rect 58 55 61 57
rect 53 38 61 55
rect 63 57 71 66
rect 63 55 66 57
rect 68 55 71 57
rect 63 50 71 55
rect 63 48 66 50
rect 68 48 71 50
rect 63 38 71 48
rect 73 49 81 66
rect 73 47 76 49
rect 78 47 81 49
rect 73 42 81 47
rect 73 40 76 42
rect 78 40 81 42
rect 73 38 81 40
rect 83 57 91 66
rect 83 55 86 57
rect 88 55 91 57
rect 83 50 91 55
rect 83 48 86 50
rect 88 48 91 50
rect 83 38 91 48
rect 93 49 101 66
rect 93 47 96 49
rect 98 47 101 49
rect 93 42 101 47
rect 93 40 96 42
rect 98 40 101 42
rect 93 38 101 40
rect 103 38 108 66
rect 110 64 121 66
rect 110 62 114 64
rect 116 62 121 64
rect 110 38 121 62
rect 123 38 128 66
rect 130 49 138 66
rect 130 47 133 49
rect 135 47 138 49
rect 130 38 138 47
rect 140 38 145 66
rect 147 64 157 66
rect 147 62 151 64
rect 153 62 157 64
rect 147 38 157 62
rect 159 57 167 66
rect 159 55 162 57
rect 164 55 167 57
rect 159 50 167 55
rect 159 48 162 50
rect 164 48 167 50
rect 159 38 167 48
rect 169 64 177 66
rect 169 62 172 64
rect 174 62 177 64
rect 169 57 177 62
rect 169 55 172 57
rect 174 55 177 57
rect 169 38 177 55
rect 179 51 184 66
rect 179 49 186 51
rect 179 47 182 49
rect 184 47 186 49
rect 179 42 186 47
rect 179 40 182 42
rect 184 40 186 42
rect 179 38 186 40
<< alu1 >>
rect -2 67 202 72
rect -2 65 5 67
rect 7 65 190 67
rect 192 65 202 67
rect -2 64 202 65
rect 74 49 79 51
rect 74 47 76 49
rect 78 47 79 49
rect 74 43 79 47
rect 94 49 158 50
rect 94 47 96 49
rect 98 47 133 49
rect 135 47 158 49
rect 94 46 158 47
rect 94 43 99 46
rect 2 33 22 35
rect 2 31 12 33
rect 14 31 19 33
rect 21 31 22 33
rect 2 29 22 31
rect 66 35 70 43
rect 74 42 99 43
rect 74 40 76 42
rect 78 40 96 42
rect 98 40 99 42
rect 74 39 99 40
rect 82 38 99 39
rect 113 38 150 42
rect 66 33 78 35
rect 66 31 73 33
rect 75 31 78 33
rect 2 21 6 29
rect 66 29 78 31
rect 82 25 86 38
rect 113 33 119 38
rect 113 31 115 33
rect 117 31 119 33
rect 113 30 119 31
rect 146 33 150 38
rect 146 31 147 33
rect 149 31 150 33
rect 146 29 150 31
rect 74 24 100 25
rect 74 22 76 24
rect 78 22 96 24
rect 98 22 100 24
rect 154 25 158 46
rect 131 24 158 25
rect 131 22 133 24
rect 135 22 158 24
rect 74 21 100 22
rect 131 21 158 22
rect -2 7 202 8
rect -2 5 5 7
rect 7 5 114 7
rect 116 5 187 7
rect 189 5 202 7
rect -2 0 202 5
<< ptie >>
rect 3 15 9 24
rect 3 13 5 15
rect 7 13 9 15
rect 3 7 9 13
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 185 15 191 24
rect 185 13 187 15
rect 189 13 191 15
rect 185 7 191 13
rect 185 5 187 7
rect 189 5 191 7
rect 185 3 191 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 188 67 194 69
rect 3 59 9 65
rect 3 57 5 59
rect 7 57 9 59
rect 3 55 9 57
rect 188 65 190 67
rect 192 65 194 67
rect 188 59 194 65
rect 188 57 190 59
rect 192 57 194 59
rect 188 55 194 57
<< nmos >>
rect 21 10 23 26
rect 31 10 33 26
rect 41 12 43 26
rect 51 12 53 26
rect 61 12 63 26
rect 71 12 73 26
rect 81 12 83 26
rect 91 12 93 26
rect 101 12 103 26
rect 108 12 110 26
rect 121 12 123 26
rect 128 12 130 26
rect 138 12 140 26
rect 145 12 147 26
rect 158 6 160 26
rect 168 6 170 26
<< pmos >>
rect 10 38 12 46
rect 21 38 23 66
rect 31 38 33 66
rect 41 38 43 66
rect 51 38 53 66
rect 61 38 63 66
rect 71 38 73 66
rect 81 38 83 66
rect 91 38 93 66
rect 101 38 103 66
rect 108 38 110 66
rect 121 38 123 66
rect 128 38 130 66
rect 138 38 140 66
rect 145 38 147 66
rect 157 38 159 66
rect 167 38 169 66
rect 177 38 179 66
<< polyct0 >>
rect 43 31 45 33
rect 50 31 52 33
rect 99 31 101 33
rect 130 31 132 33
<< polyct1 >>
rect 12 31 14 33
rect 19 31 21 33
rect 73 31 75 33
rect 115 31 117 33
rect 147 31 149 33
<< ndifct0 >>
rect 16 21 18 23
rect 16 14 18 16
rect 26 22 28 24
rect 26 15 28 17
rect 36 21 38 23
rect 36 14 38 16
rect 46 22 48 24
rect 46 15 48 17
rect 56 14 58 16
rect 66 22 68 24
rect 66 15 68 17
rect 86 15 88 17
rect 151 8 153 10
rect 163 22 165 24
rect 163 15 165 17
rect 173 16 175 18
rect 173 8 175 10
<< ndifct1 >>
rect 76 22 78 24
rect 96 22 98 24
rect 133 22 135 24
rect 114 5 116 7
<< ntiect0 >>
rect 5 57 7 59
rect 190 57 192 59
<< ntiect1 >>
rect 5 65 7 67
rect 190 65 192 67
<< ptiect0 >>
rect 5 13 7 15
rect 187 13 189 15
<< ptiect1 >>
rect 5 5 7 7
rect 187 5 189 7
<< pdifct0 >>
rect 16 62 18 64
rect 16 55 18 57
rect 16 48 18 50
rect 5 40 7 42
rect 26 47 28 49
rect 26 40 28 42
rect 36 62 38 64
rect 36 55 38 57
rect 36 48 38 50
rect 46 55 48 57
rect 46 48 48 50
rect 56 62 58 64
rect 56 55 58 57
rect 66 55 68 57
rect 66 48 68 50
rect 86 55 88 57
rect 86 48 88 50
rect 114 62 116 64
rect 151 62 153 64
rect 162 55 164 57
rect 162 48 164 50
rect 172 62 174 64
rect 172 55 174 57
rect 182 47 184 49
rect 182 40 184 42
<< pdifct1 >>
rect 76 47 78 49
rect 76 40 78 42
rect 96 47 98 49
rect 96 40 98 42
rect 133 47 135 49
<< alu0 >>
rect 4 59 8 64
rect 4 57 5 59
rect 7 57 8 59
rect 4 55 8 57
rect 15 62 16 64
rect 18 62 19 64
rect 15 57 19 62
rect 15 55 16 57
rect 18 55 19 57
rect 15 50 19 55
rect 35 62 36 64
rect 38 62 39 64
rect 35 57 39 62
rect 55 62 56 64
rect 58 62 59 64
rect 35 55 36 57
rect 38 55 39 57
rect 15 48 16 50
rect 18 48 19 50
rect 15 46 19 48
rect 25 49 29 51
rect 25 47 26 49
rect 28 47 29 49
rect 25 43 29 47
rect 35 50 39 55
rect 35 48 36 50
rect 38 48 39 50
rect 35 46 39 48
rect 45 57 49 59
rect 45 55 46 57
rect 48 55 49 57
rect 45 50 49 55
rect 55 57 59 62
rect 112 62 114 64
rect 116 62 118 64
rect 112 61 118 62
rect 149 62 151 64
rect 153 62 155 64
rect 149 61 155 62
rect 170 62 172 64
rect 174 62 176 64
rect 55 55 56 57
rect 58 55 59 57
rect 55 53 59 55
rect 64 57 166 58
rect 64 55 66 57
rect 68 55 86 57
rect 88 55 162 57
rect 164 55 166 57
rect 64 54 166 55
rect 170 57 176 62
rect 170 55 172 57
rect 174 55 176 57
rect 189 59 193 64
rect 189 57 190 59
rect 192 57 193 59
rect 189 55 193 57
rect 170 54 176 55
rect 64 50 69 54
rect 45 48 46 50
rect 48 48 66 50
rect 68 48 69 50
rect 45 46 69 48
rect 85 50 89 54
rect 161 50 166 54
rect 85 48 86 50
rect 88 48 89 50
rect 85 46 89 48
rect 161 48 162 50
rect 164 49 186 50
rect 164 48 182 49
rect 161 47 182 48
rect 184 47 186 49
rect 161 46 186 47
rect 3 42 29 43
rect 3 40 5 42
rect 7 40 26 42
rect 28 40 29 42
rect 3 39 29 40
rect 25 34 29 39
rect 25 33 54 34
rect 25 31 43 33
rect 45 31 50 33
rect 52 31 54 33
rect 25 30 54 31
rect 15 23 19 25
rect 15 21 16 23
rect 18 21 19 23
rect 4 15 8 17
rect 4 13 5 15
rect 7 13 8 15
rect 4 8 8 13
rect 15 16 19 21
rect 15 14 16 16
rect 18 14 19 16
rect 15 8 19 14
rect 25 24 29 30
rect 25 22 26 24
rect 28 22 29 24
rect 25 17 29 22
rect 25 15 26 17
rect 28 15 29 17
rect 25 13 29 15
rect 35 23 39 25
rect 35 21 36 23
rect 38 21 39 23
rect 35 16 39 21
rect 35 14 36 16
rect 38 14 39 16
rect 35 8 39 14
rect 45 24 69 26
rect 97 33 108 34
rect 97 31 99 33
rect 101 31 108 33
rect 97 30 108 31
rect 123 33 134 34
rect 123 31 130 33
rect 132 31 134 33
rect 123 30 134 31
rect 104 26 108 30
rect 123 26 127 30
rect 45 22 46 24
rect 48 22 66 24
rect 68 22 69 24
rect 45 17 49 22
rect 64 18 69 22
rect 104 22 127 26
rect 180 42 186 46
rect 180 40 182 42
rect 184 40 186 42
rect 180 39 186 40
rect 162 24 167 26
rect 162 22 163 24
rect 165 22 167 24
rect 162 18 167 22
rect 45 15 46 17
rect 48 15 49 17
rect 45 13 49 15
rect 55 16 59 18
rect 55 14 56 16
rect 58 14 59 16
rect 64 17 167 18
rect 64 15 66 17
rect 68 15 86 17
rect 88 15 163 17
rect 165 15 167 17
rect 64 14 167 15
rect 172 18 176 20
rect 172 16 173 18
rect 175 16 176 18
rect 55 8 59 14
rect 149 10 155 11
rect 149 8 151 10
rect 153 8 155 10
rect 172 10 176 16
rect 172 8 173 10
rect 175 8 176 10
rect 186 15 190 17
rect 186 13 187 15
rect 189 13 190 15
rect 186 8 190 13
<< labels >>
rlabel alu0 47 19 47 19 6 n3
rlabel alu0 16 41 16 41 6 bn
rlabel alu0 47 52 47 52 6 n1
rlabel alu0 66 20 66 20 6 n3
rlabel alu0 39 32 39 32 6 bn
rlabel alu0 87 52 87 52 6 n1
rlabel alu0 66 52 66 52 6 n1
rlabel alu0 102 32 102 32 6 bn
rlabel alu0 128 32 128 32 6 bn
rlabel alu0 115 16 115 16 6 n3
rlabel alu0 164 20 164 20 6 n3
rlabel alu0 183 44 183 44 6 n1
rlabel alu0 163 52 163 52 6 n1
rlabel alu0 115 56 115 56 6 n1
rlabel polyct1 20 32 20 32 6 b
rlabel alu1 12 32 12 32 6 b
rlabel alu1 4 28 4 28 6 b
rlabel alu1 76 32 76 32 6 c
rlabel alu1 68 36 68 36 6 c
rlabel alu1 76 48 76 48 6 z
rlabel alu1 100 4 100 4 6 vss
rlabel alu1 84 32 84 32 6 z
rlabel alu1 92 40 92 40 6 z
rlabel alu1 116 36 116 36 6 a
rlabel alu1 108 48 108 48 6 z
rlabel alu1 100 48 100 48 6 z
rlabel alu1 116 48 116 48 6 z
rlabel alu1 100 68 100 68 6 vdd
rlabel alu1 156 32 156 32 6 z
rlabel polyct1 148 32 148 32 6 a
rlabel alu1 124 40 124 40 6 a
rlabel alu1 140 40 140 40 6 a
rlabel alu1 132 40 132 40 6 a
rlabel alu1 124 48 124 48 6 z
rlabel alu1 132 48 132 48 6 z
rlabel alu1 148 48 148 48 6 z
rlabel alu1 140 48 140 48 6 z
<< end >>
