magic
tech scmos
timestamp 1199470180
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -5 48 55 105
<< pwell >>
rect -5 -5 55 48
<< poly >>
rect 25 84 27 89
rect 33 84 35 89
rect 13 73 15 78
rect 13 53 15 61
rect 13 51 21 53
rect 13 49 17 51
rect 19 49 21 51
rect 13 47 21 49
rect 13 27 15 47
rect 25 43 27 61
rect 33 53 35 61
rect 33 51 43 53
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 25 41 33 43
rect 25 39 29 41
rect 31 39 33 41
rect 25 37 33 39
rect 25 27 27 37
rect 37 27 39 47
rect 13 12 15 17
rect 25 12 27 17
rect 37 12 39 17
<< ndif >>
rect 8 23 13 27
rect 5 21 13 23
rect 5 19 7 21
rect 9 19 13 21
rect 5 17 13 19
rect 15 21 25 27
rect 15 19 19 21
rect 21 19 25 21
rect 15 17 25 19
rect 27 17 37 27
rect 39 23 44 27
rect 39 21 47 23
rect 39 19 43 21
rect 45 19 47 21
rect 39 17 47 19
rect 29 11 35 17
rect 29 9 31 11
rect 33 9 35 11
rect 29 7 35 9
<< pdif >>
rect 20 73 25 84
rect 5 71 13 73
rect 5 69 7 71
rect 9 69 13 71
rect 5 61 13 69
rect 15 71 25 73
rect 15 69 19 71
rect 21 69 25 71
rect 15 61 25 69
rect 27 61 33 84
rect 35 81 43 84
rect 35 79 39 81
rect 41 79 43 81
rect 35 61 43 79
<< alu1 >>
rect -2 95 52 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 52 95
rect -2 88 52 93
rect 6 71 10 88
rect 38 81 42 88
rect 38 79 39 81
rect 41 79 42 81
rect 38 77 42 79
rect 6 69 7 71
rect 9 69 10 71
rect 6 67 10 69
rect 18 71 22 73
rect 18 69 19 71
rect 21 69 22 71
rect 18 63 22 69
rect 27 68 42 73
rect 8 57 22 63
rect 8 23 12 57
rect 16 51 22 53
rect 16 49 17 51
rect 19 49 22 51
rect 16 47 22 49
rect 18 32 22 47
rect 28 42 32 63
rect 38 51 42 68
rect 38 49 39 51
rect 41 49 42 51
rect 38 47 42 49
rect 28 41 43 42
rect 28 39 29 41
rect 31 39 43 41
rect 28 37 43 39
rect 18 27 33 32
rect 5 21 12 23
rect 5 19 7 21
rect 9 19 12 21
rect 5 17 12 19
rect 17 21 47 22
rect 17 19 19 21
rect 21 19 43 21
rect 45 19 47 21
rect 17 18 47 19
rect -2 11 52 12
rect -2 9 31 11
rect 33 9 52 11
rect -2 7 52 9
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 52 7
rect -2 0 52 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 13 17 15 27
rect 25 17 27 27
rect 37 17 39 27
<< pmos >>
rect 13 61 15 73
rect 25 61 27 84
rect 33 61 35 84
<< polyct1 >>
rect 17 49 19 51
rect 39 49 41 51
rect 29 39 31 41
<< ndifct1 >>
rect 7 19 9 21
rect 19 19 21 21
rect 43 19 45 21
rect 31 9 33 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 7 69 9 71
rect 19 69 21 71
rect 39 79 41 81
<< labels >>
rlabel ndifct1 20 20 20 20 6 n2
rlabel ndifct1 44 20 44 20 6 n2
rlabel alu1 10 40 10 40 6 z
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 65 20 65 6 z
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 30 30 30 6 b
rlabel alu1 30 50 30 50 6 a2
rlabel alu1 30 70 30 70 6 a1
rlabel alu1 25 94 25 94 6 vdd
rlabel alu1 40 40 40 40 6 a2
rlabel alu1 40 60 40 60 6 a1
<< end >>
