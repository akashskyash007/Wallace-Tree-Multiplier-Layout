magic
tech scmos
timestamp 1199201696
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 61 31 66
rect 39 61 41 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 46
rect 39 43 41 46
rect 39 41 47 43
rect 39 39 43 41
rect 45 39 47 41
rect 9 37 22 39
rect 9 35 18 37
rect 20 35 22 37
rect 9 33 22 35
rect 28 37 34 39
rect 28 35 30 37
rect 32 35 34 37
rect 28 33 34 35
rect 10 30 12 33
rect 20 30 22 33
rect 32 30 34 33
rect 39 37 47 39
rect 39 30 41 37
rect 10 11 12 16
rect 20 11 22 16
rect 32 13 34 18
rect 39 13 41 18
<< ndif >>
rect 2 16 10 30
rect 12 21 20 30
rect 12 19 15 21
rect 17 19 20 21
rect 12 16 20 19
rect 22 18 32 30
rect 34 18 39 30
rect 41 24 46 30
rect 41 22 48 24
rect 41 20 44 22
rect 46 20 48 22
rect 41 18 48 20
rect 22 16 30 18
rect 2 11 8 16
rect 24 11 30 16
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
rect 24 9 26 11
rect 28 9 30 11
rect 24 7 30 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 61 27 70
rect 21 59 29 61
rect 21 57 24 59
rect 26 57 29 59
rect 21 46 29 57
rect 31 59 39 61
rect 31 57 34 59
rect 36 57 39 59
rect 31 52 39 57
rect 31 50 34 52
rect 36 50 39 52
rect 31 46 39 50
rect 41 59 48 61
rect 41 57 44 59
rect 46 57 48 59
rect 41 52 48 57
rect 41 50 44 52
rect 46 50 48 52
rect 41 46 48 50
rect 21 42 27 46
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 22 6 50
rect 33 42 46 46
rect 42 41 46 42
rect 42 39 43 41
rect 45 39 46 41
rect 25 37 38 38
rect 25 35 30 37
rect 32 35 38 37
rect 25 34 38 35
rect 2 21 19 22
rect 2 19 15 21
rect 17 19 19 21
rect 2 17 19 19
rect 34 25 38 34
rect 42 33 46 39
rect -2 11 58 12
rect -2 9 4 11
rect 6 9 26 11
rect 28 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 10 16 12 30
rect 20 16 22 30
rect 32 18 34 30
rect 39 18 41 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 46 31 61
rect 39 46 41 61
<< polyct0 >>
rect 18 35 20 37
<< polyct1 >>
rect 43 39 45 41
rect 30 35 32 37
<< ndifct0 >>
rect 44 20 46 22
<< ndifct1 >>
rect 15 19 17 21
rect 4 9 6 11
rect 26 9 28 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 57 26 59
rect 34 57 36 59
rect 34 50 36 52
rect 44 57 46 59
rect 44 50 46 52
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 59 28 68
rect 22 57 24 59
rect 26 57 28 59
rect 22 56 28 57
rect 32 59 38 60
rect 32 57 34 59
rect 36 57 38 59
rect 32 53 38 57
rect 23 52 38 53
rect 23 50 34 52
rect 36 50 38 52
rect 23 49 38 50
rect 42 59 48 68
rect 42 57 44 59
rect 46 57 48 59
rect 42 52 48 57
rect 42 50 44 52
rect 46 50 48 52
rect 42 49 48 50
rect 23 46 27 49
rect 17 42 27 46
rect 17 37 21 42
rect 17 35 18 37
rect 20 35 21 37
rect 17 30 21 35
rect 17 26 28 30
rect 24 21 28 26
rect 43 22 47 24
rect 43 21 44 22
rect 24 20 44 21
rect 46 20 47 22
rect 24 17 47 20
<< labels >>
rlabel polyct0 19 36 19 36 6 zn
rlabel alu0 30 51 30 51 6 zn
rlabel alu0 35 54 35 54 6 zn
rlabel alu0 35 19 35 19 6 zn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 36 28 36 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 36 44 36 6 b
<< end >>
