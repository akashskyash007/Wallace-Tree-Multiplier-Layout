magic
tech scmos
timestamp 1199542433
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -5 48 105 105
<< pwell >>
rect -5 -5 105 48
<< poly >>
rect 23 94 25 98
rect 35 94 37 98
rect 11 76 13 80
rect 11 53 13 56
rect 51 85 53 89
rect 63 86 65 90
rect 75 85 77 89
rect 87 85 89 89
rect 11 51 19 53
rect 11 49 15 51
rect 17 49 19 51
rect 11 47 19 49
rect 23 43 25 55
rect 35 43 37 55
rect 9 41 37 43
rect 9 39 11 41
rect 13 39 37 41
rect 9 37 37 39
rect 11 31 19 33
rect 11 29 15 31
rect 17 29 19 31
rect 11 27 19 29
rect 11 24 13 27
rect 23 25 25 37
rect 35 25 37 37
rect 51 33 53 65
rect 63 63 65 66
rect 59 61 65 63
rect 59 43 61 61
rect 75 53 77 65
rect 67 51 77 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 47 31 53 33
rect 47 29 49 31
rect 51 29 53 31
rect 47 27 53 29
rect 11 10 13 14
rect 51 24 53 27
rect 59 24 61 37
rect 67 24 69 47
rect 77 41 83 43
rect 77 39 79 41
rect 81 39 83 41
rect 87 39 89 65
rect 75 37 89 39
rect 75 24 77 37
rect 23 2 25 6
rect 35 2 37 6
rect 51 2 53 6
rect 59 2 61 6
rect 67 2 69 6
rect 75 2 77 6
<< ndif >>
rect 18 24 23 25
rect 3 21 11 24
rect 3 19 5 21
rect 7 19 11 21
rect 3 14 11 19
rect 13 14 23 24
rect 15 11 23 14
rect 15 9 17 11
rect 19 9 23 11
rect 15 6 23 9
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 6 35 19
rect 37 24 45 25
rect 79 24 93 25
rect 37 11 51 24
rect 37 9 43 11
rect 45 9 51 11
rect 37 6 51 9
rect 53 6 59 24
rect 61 6 67 24
rect 69 6 75 24
rect 77 21 93 24
rect 77 19 89 21
rect 91 19 93 21
rect 77 15 93 19
rect 77 6 85 15
<< pdif >>
rect 15 91 23 94
rect 15 89 17 91
rect 19 89 23 91
rect 15 76 23 89
rect 3 71 11 76
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 56 11 59
rect 13 56 23 76
rect 18 55 23 56
rect 25 71 35 94
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 91 49 94
rect 37 89 43 91
rect 45 89 49 91
rect 67 91 73 93
rect 37 85 49 89
rect 67 89 69 91
rect 71 89 73 91
rect 91 91 97 93
rect 91 89 93 91
rect 95 89 97 91
rect 67 86 73 89
rect 55 85 63 86
rect 37 65 51 85
rect 53 81 63 85
rect 53 79 57 81
rect 59 79 63 81
rect 53 66 63 79
rect 65 85 73 86
rect 91 85 97 89
rect 65 66 75 85
rect 53 65 58 66
rect 37 55 45 65
rect 70 65 75 66
rect 77 81 87 85
rect 77 79 81 81
rect 83 79 87 81
rect 77 65 87 79
rect 89 65 97 85
<< alu1 >>
rect -2 95 102 100
rect -2 93 5 95
rect 7 93 102 95
rect -2 91 102 93
rect -2 89 17 91
rect 19 89 43 91
rect 45 89 69 91
rect 71 89 93 91
rect 95 89 102 91
rect -2 88 102 89
rect 19 81 93 82
rect 19 79 57 81
rect 59 79 81 81
rect 83 79 93 81
rect 19 78 93 79
rect 4 71 8 73
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 4 59 5 61
rect 7 59 8 61
rect 4 42 8 59
rect 19 52 23 78
rect 13 51 23 52
rect 13 49 15 51
rect 17 49 23 51
rect 13 48 23 49
rect 4 41 15 42
rect 4 39 11 41
rect 13 39 15 41
rect 4 38 15 39
rect 4 21 8 38
rect 19 32 23 48
rect 13 31 23 32
rect 13 29 15 31
rect 17 29 23 31
rect 13 28 23 29
rect 28 71 32 73
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 4 19 5 21
rect 7 19 8 21
rect 4 17 8 19
rect 28 21 32 59
rect 28 19 29 21
rect 31 19 32 21
rect 28 17 32 19
rect 48 31 52 73
rect 48 29 49 31
rect 51 29 52 31
rect 48 17 52 29
rect 58 41 62 73
rect 58 39 59 41
rect 61 39 62 41
rect 58 17 62 39
rect 68 51 72 73
rect 68 49 69 51
rect 71 49 72 51
rect 68 17 72 49
rect 78 41 82 73
rect 78 39 79 41
rect 81 39 82 41
rect 78 17 82 39
rect 89 22 93 78
rect 87 21 93 22
rect 87 19 89 21
rect 91 19 93 21
rect 87 18 93 19
rect -2 11 102 12
rect -2 9 17 11
rect 19 9 43 11
rect 45 9 102 11
rect -2 0 102 9
<< ntie >>
rect 3 95 9 97
rect 3 93 5 95
rect 7 93 9 95
rect 3 86 9 93
<< nmos >>
rect 11 14 13 24
rect 23 6 25 25
rect 35 6 37 25
rect 51 6 53 24
rect 59 6 61 24
rect 67 6 69 24
rect 75 6 77 24
<< pmos >>
rect 11 56 13 76
rect 23 55 25 94
rect 35 55 37 94
rect 51 65 53 85
rect 63 66 65 86
rect 75 65 77 85
rect 87 65 89 85
<< polyct1 >>
rect 15 49 17 51
rect 11 39 13 41
rect 15 29 17 31
rect 69 49 71 51
rect 59 39 61 41
rect 49 29 51 31
rect 79 39 81 41
<< ndifct1 >>
rect 5 19 7 21
rect 17 9 19 11
rect 29 19 31 21
rect 43 9 45 11
rect 89 19 91 21
<< ntiect1 >>
rect 5 93 7 95
<< pdifct1 >>
rect 17 89 19 91
rect 5 69 7 71
rect 5 59 7 61
rect 29 69 31 71
rect 29 59 31 61
rect 43 89 45 91
rect 69 89 71 91
rect 93 89 95 91
rect 57 79 59 81
rect 81 79 83 81
<< labels >>
rlabel alu1 30 45 30 45 6 nq
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 50 45 50 45 6 i0
rlabel alu1 70 45 70 45 6 i2
rlabel alu1 60 45 60 45 6 i1
rlabel alu1 50 94 50 94 6 vdd
rlabel alu1 80 45 80 45 6 i3
<< end >>
