magic
tech scmos
timestamp 1199543355
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 57 94 59 98
rect 11 85 13 89
rect 19 85 21 89
rect 27 85 29 89
rect 35 85 37 89
rect 11 43 13 56
rect 19 43 21 56
rect 27 43 29 56
rect 35 53 37 56
rect 35 51 43 53
rect 41 43 43 51
rect 57 43 59 55
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 47 41 59 43
rect 47 39 49 41
rect 51 39 59 41
rect 47 37 59 39
rect 11 25 13 37
rect 19 29 21 37
rect 31 29 33 37
rect 41 29 43 37
rect 19 27 25 29
rect 31 27 37 29
rect 41 27 49 29
rect 23 24 25 27
rect 35 24 37 27
rect 47 24 49 27
rect 57 25 59 37
rect 11 11 13 15
rect 23 10 25 14
rect 35 10 37 14
rect 47 11 49 15
rect 57 2 59 6
<< ndif >>
rect 3 15 11 25
rect 13 24 18 25
rect 52 24 57 25
rect 13 21 23 24
rect 13 19 17 21
rect 19 19 23 21
rect 13 15 23 19
rect 3 11 9 15
rect 15 14 23 15
rect 25 14 35 24
rect 37 21 47 24
rect 37 19 41 21
rect 43 19 47 21
rect 37 15 47 19
rect 49 15 57 24
rect 37 14 45 15
rect 3 9 5 11
rect 7 9 9 11
rect 27 11 33 14
rect 3 7 9 9
rect 27 9 29 11
rect 31 9 33 11
rect 51 9 57 15
rect 27 7 33 9
rect 49 7 57 9
rect 49 5 51 7
rect 53 6 57 7
rect 59 21 67 25
rect 59 19 63 21
rect 65 19 67 21
rect 59 6 67 19
rect 53 5 55 6
rect 49 3 55 5
<< pdif >>
rect 39 91 57 94
rect 39 89 43 91
rect 45 89 51 91
rect 53 89 57 91
rect 39 85 57 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 56 11 79
rect 13 56 19 85
rect 21 56 27 85
rect 29 56 35 85
rect 37 56 57 85
rect 47 55 57 56
rect 59 81 67 94
rect 59 79 63 81
rect 65 79 67 81
rect 59 71 67 79
rect 59 69 63 71
rect 65 69 67 71
rect 59 61 67 69
rect 59 59 63 61
rect 65 59 67 61
rect 59 55 67 59
<< alu1 >>
rect -2 95 72 100
rect -2 93 5 95
rect 7 93 17 95
rect 19 93 29 95
rect 31 93 72 95
rect -2 91 72 93
rect -2 89 43 91
rect 45 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 58 82 62 83
rect 3 81 53 82
rect 3 79 5 81
rect 7 79 53 81
rect 3 78 53 79
rect 8 41 12 73
rect 8 39 9 41
rect 11 39 12 41
rect 8 27 12 39
rect 18 41 22 73
rect 18 39 19 41
rect 21 39 22 41
rect 18 27 22 39
rect 28 41 32 73
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 41 42 73
rect 49 42 53 78
rect 38 39 39 41
rect 41 39 42 41
rect 38 27 42 39
rect 47 41 53 42
rect 47 39 49 41
rect 51 39 53 41
rect 47 38 53 39
rect 49 22 53 38
rect 15 21 53 22
rect 15 19 17 21
rect 19 19 41 21
rect 43 19 53 21
rect 15 18 53 19
rect 58 81 67 82
rect 58 79 63 81
rect 65 79 67 81
rect 58 78 67 79
rect 58 72 62 78
rect 58 71 67 72
rect 58 69 63 71
rect 65 69 67 71
rect 58 68 67 69
rect 58 62 62 68
rect 58 61 67 62
rect 58 59 63 61
rect 65 59 67 61
rect 58 58 67 59
rect 58 22 62 58
rect 58 21 67 22
rect 58 19 63 21
rect 65 19 67 21
rect 58 18 67 19
rect 58 17 62 18
rect -2 11 72 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 72 11
rect -2 7 72 9
rect -2 5 51 7
rect 53 5 72 7
rect -2 0 72 5
<< ntie >>
rect 3 95 33 97
rect 3 93 5 95
rect 7 93 17 95
rect 19 93 29 95
rect 31 93 33 95
rect 3 91 33 93
<< nmos >>
rect 11 15 13 25
rect 23 14 25 24
rect 35 14 37 24
rect 47 15 49 24
rect 57 6 59 25
<< pmos >>
rect 11 56 13 85
rect 19 56 21 85
rect 27 56 29 85
rect 35 56 37 85
rect 57 55 59 94
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 39 39 41 41
rect 49 39 51 41
<< ndifct1 >>
rect 17 19 19 21
rect 41 19 43 21
rect 5 9 7 11
rect 29 9 31 11
rect 51 5 53 7
rect 63 19 65 21
<< ntiect1 >>
rect 5 93 7 95
rect 17 93 19 95
rect 29 93 31 95
<< pdifct1 >>
rect 43 89 45 91
rect 51 89 53 91
rect 5 79 7 81
rect 63 79 65 81
rect 63 69 65 71
rect 63 59 65 61
<< labels >>
rlabel alu1 10 50 10 50 6 i3
rlabel alu1 30 50 30 50 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 50 40 50 6 i2
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 50 60 50 6 q
<< end >>
