magic
tech scmos
timestamp 1199541705
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 55 94 57 98
rect 67 94 69 98
rect 11 86 13 90
rect 31 85 33 89
rect 43 85 45 89
rect 11 63 13 66
rect 11 61 23 63
rect 17 59 19 61
rect 21 59 23 61
rect 17 57 23 59
rect 3 51 9 53
rect 31 51 33 65
rect 3 49 5 51
rect 7 49 33 51
rect 3 47 9 49
rect 31 29 33 49
rect 43 53 45 65
rect 43 51 51 53
rect 43 49 47 51
rect 49 49 51 51
rect 43 47 51 49
rect 37 41 43 43
rect 55 41 57 55
rect 67 41 69 55
rect 37 39 39 41
rect 41 39 69 41
rect 37 37 43 39
rect 43 31 51 33
rect 43 29 47 31
rect 49 29 51 31
rect 31 27 37 29
rect 17 25 23 27
rect 17 23 19 25
rect 21 23 23 25
rect 35 24 37 27
rect 43 27 51 29
rect 43 24 45 27
rect 55 25 57 39
rect 67 25 69 39
rect 11 21 23 23
rect 11 18 13 21
rect 11 4 13 8
rect 35 2 37 6
rect 43 2 45 6
rect 55 2 57 6
rect 67 2 69 6
<< ndif >>
rect 50 24 55 25
rect 3 21 9 23
rect 3 19 5 21
rect 7 19 9 21
rect 3 18 9 19
rect 27 21 35 24
rect 27 19 29 21
rect 31 19 35 21
rect 3 8 11 18
rect 13 11 21 18
rect 13 9 17 11
rect 19 9 21 11
rect 13 8 21 9
rect 15 7 21 8
rect 27 6 35 19
rect 37 6 43 24
rect 45 11 55 24
rect 45 9 49 11
rect 51 9 55 11
rect 45 6 55 9
rect 57 21 67 25
rect 57 19 61 21
rect 63 19 67 21
rect 57 6 67 19
rect 69 21 77 25
rect 69 19 73 21
rect 75 19 77 21
rect 69 11 77 19
rect 69 9 73 11
rect 75 9 77 11
rect 69 6 77 9
<< pdif >>
rect 15 91 29 93
rect 15 89 17 91
rect 19 89 25 91
rect 27 89 29 91
rect 47 91 55 94
rect 47 89 49 91
rect 51 89 55 91
rect 15 86 29 89
rect 3 81 11 86
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 66 11 69
rect 13 85 29 86
rect 47 85 55 89
rect 13 66 31 85
rect 15 65 31 66
rect 33 81 43 85
rect 33 79 37 81
rect 39 79 43 81
rect 33 71 43 79
rect 33 69 37 71
rect 39 69 43 71
rect 33 65 43 69
rect 45 65 55 85
rect 47 55 55 65
rect 57 81 67 94
rect 57 79 61 81
rect 63 79 67 81
rect 57 71 67 79
rect 57 69 61 71
rect 63 69 67 71
rect 57 61 67 69
rect 57 59 61 61
rect 63 59 67 61
rect 57 55 67 59
rect 69 91 77 94
rect 69 89 73 91
rect 75 89 77 91
rect 69 81 77 89
rect 69 79 73 81
rect 75 79 77 81
rect 69 71 77 79
rect 69 69 73 71
rect 75 69 77 71
rect 69 61 77 69
rect 69 59 73 61
rect 75 59 77 61
rect 69 55 77 59
<< alu1 >>
rect -2 91 82 100
rect -2 89 17 91
rect 19 89 25 91
rect 27 89 49 91
rect 51 89 73 91
rect 75 89 82 91
rect -2 88 82 89
rect 4 81 8 83
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 4 69 5 71
rect 7 69 8 71
rect 4 51 8 69
rect 4 49 5 51
rect 7 49 8 51
rect 4 21 8 49
rect 4 19 5 21
rect 7 19 8 21
rect 4 17 8 19
rect 18 61 22 83
rect 35 81 41 82
rect 35 79 37 81
rect 39 79 41 81
rect 35 78 41 79
rect 37 72 41 78
rect 35 71 41 72
rect 35 69 37 71
rect 39 69 41 71
rect 35 68 41 69
rect 18 59 19 61
rect 21 59 22 61
rect 18 25 22 59
rect 18 23 19 25
rect 21 23 22 25
rect 18 17 22 23
rect 37 42 41 68
rect 48 52 52 83
rect 45 51 52 52
rect 45 49 47 51
rect 49 49 52 51
rect 45 48 52 49
rect 37 41 43 42
rect 37 39 39 41
rect 41 39 43 41
rect 37 38 43 39
rect 37 22 41 38
rect 48 32 52 48
rect 45 31 52 32
rect 45 29 47 31
rect 49 29 52 31
rect 45 28 52 29
rect 27 21 41 22
rect 27 19 29 21
rect 31 19 41 21
rect 27 18 41 19
rect 48 17 52 28
rect 58 82 62 83
rect 58 81 65 82
rect 58 79 61 81
rect 63 79 65 81
rect 58 78 65 79
rect 72 81 76 88
rect 72 79 73 81
rect 75 79 76 81
rect 58 72 62 78
rect 58 71 65 72
rect 58 69 61 71
rect 63 69 65 71
rect 58 68 65 69
rect 72 71 76 79
rect 72 69 73 71
rect 75 69 76 71
rect 58 62 62 68
rect 58 61 65 62
rect 58 59 61 61
rect 63 59 65 61
rect 58 58 65 59
rect 72 61 76 69
rect 72 59 73 61
rect 75 59 76 61
rect 58 22 62 58
rect 72 57 76 59
rect 58 21 65 22
rect 58 19 61 21
rect 63 19 65 21
rect 58 18 65 19
rect 72 21 76 23
rect 72 19 73 21
rect 75 19 76 21
rect 58 17 62 18
rect 72 12 76 19
rect -2 11 82 12
rect -2 9 17 11
rect 19 9 49 11
rect 51 9 73 11
rect 75 9 82 11
rect -2 0 82 9
<< nmos >>
rect 11 8 13 18
rect 35 6 37 24
rect 43 6 45 24
rect 55 6 57 25
rect 67 6 69 25
<< pmos >>
rect 11 66 13 86
rect 31 65 33 85
rect 43 65 45 85
rect 55 55 57 94
rect 67 55 69 94
<< polyct1 >>
rect 19 59 21 61
rect 5 49 7 51
rect 47 49 49 51
rect 39 39 41 41
rect 47 29 49 31
rect 19 23 21 25
<< ndifct1 >>
rect 5 19 7 21
rect 29 19 31 21
rect 17 9 19 11
rect 49 9 51 11
rect 61 19 63 21
rect 73 19 75 21
rect 73 9 75 11
<< pdifct1 >>
rect 17 89 19 91
rect 25 89 27 91
rect 49 89 51 91
rect 5 79 7 81
rect 5 69 7 71
rect 37 79 39 81
rect 37 69 39 71
rect 61 79 63 81
rect 61 69 63 71
rect 61 59 63 61
rect 73 89 75 91
rect 73 79 75 81
rect 73 69 75 71
rect 73 59 75 61
<< labels >>
rlabel alu1 20 50 20 50 6 i0
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 50 50 50 50 6 i1
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 60 50 60 50 6 q
<< end >>
