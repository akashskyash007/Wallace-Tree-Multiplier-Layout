magic
tech scmos
timestamp 1199542521
<< ab >>
rect 0 0 110 100
<< nwell >>
rect -5 48 115 105
<< pwell >>
rect -5 -5 115 48
<< poly >>
rect 83 94 85 98
rect 95 94 97 98
rect 11 85 13 89
rect 23 85 25 89
rect 35 85 37 89
rect 47 85 49 89
rect 71 76 73 80
rect 11 43 13 65
rect 23 43 25 65
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 25 43
rect 17 39 19 41
rect 21 39 25 41
rect 17 37 25 39
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 65
rect 47 43 49 65
rect 71 53 73 56
rect 71 51 79 53
rect 71 49 75 51
rect 77 49 79 51
rect 71 47 79 49
rect 35 41 43 43
rect 35 39 39 41
rect 41 39 43 41
rect 35 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 35 25 37 37
rect 47 25 49 37
rect 71 25 73 47
rect 83 43 85 55
rect 95 43 97 55
rect 77 41 97 43
rect 77 39 79 41
rect 81 39 97 41
rect 77 37 97 39
rect 83 25 85 37
rect 95 25 97 37
rect 11 11 13 15
rect 23 11 25 15
rect 35 11 37 15
rect 47 11 49 15
rect 71 11 73 15
rect 83 2 85 6
rect 95 2 97 6
<< ndif >>
rect 15 31 21 33
rect 15 29 17 31
rect 19 29 21 31
rect 15 25 21 29
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 15 35 19
rect 37 15 47 25
rect 49 21 57 25
rect 49 19 53 21
rect 55 19 57 21
rect 49 15 57 19
rect 63 21 71 25
rect 63 19 65 21
rect 67 19 71 21
rect 63 15 71 19
rect 73 21 83 25
rect 73 19 77 21
rect 79 19 83 21
rect 73 15 83 19
rect 39 11 45 15
rect 75 11 83 15
rect 39 9 41 11
rect 43 9 45 11
rect 75 9 77 11
rect 79 9 83 11
rect 39 7 45 9
rect 75 6 83 9
rect 85 21 95 25
rect 85 19 89 21
rect 91 19 95 21
rect 85 6 95 19
rect 97 21 105 25
rect 97 19 101 21
rect 103 19 105 21
rect 97 11 105 19
rect 97 9 101 11
rect 103 9 105 11
rect 97 6 105 9
<< pdif >>
rect 3 91 9 93
rect 51 91 57 93
rect 3 89 5 91
rect 7 89 9 91
rect 51 89 53 91
rect 55 89 57 91
rect 3 85 9 89
rect 51 85 57 89
rect 75 91 83 94
rect 75 89 77 91
rect 79 89 83 91
rect 3 65 11 85
rect 13 65 23 85
rect 25 81 35 85
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 65 35 69
rect 37 65 47 85
rect 49 65 57 85
rect 75 81 83 89
rect 75 79 77 81
rect 79 79 83 81
rect 75 76 83 79
rect 63 61 71 76
rect 63 59 65 61
rect 67 59 71 61
rect 63 56 71 59
rect 73 56 83 76
rect 78 55 83 56
rect 85 81 95 94
rect 85 79 89 81
rect 91 79 95 81
rect 85 71 95 79
rect 85 69 89 71
rect 91 69 95 71
rect 85 61 95 69
rect 85 59 89 61
rect 91 59 95 61
rect 85 55 95 59
rect 97 91 105 94
rect 97 89 101 91
rect 103 89 105 91
rect 97 81 105 89
rect 97 79 101 81
rect 103 79 105 81
rect 97 71 105 79
rect 97 69 101 71
rect 103 69 105 71
rect 97 61 105 69
rect 97 59 101 61
rect 103 59 105 61
rect 97 55 105 59
<< alu1 >>
rect -2 95 112 100
rect -2 93 17 95
rect 19 93 29 95
rect 31 93 41 95
rect 43 93 65 95
rect 67 93 112 95
rect -2 91 112 93
rect -2 89 5 91
rect 7 89 53 91
rect 55 89 77 91
rect 79 89 101 91
rect 103 89 112 91
rect -2 88 112 89
rect 8 41 12 83
rect 8 39 9 41
rect 11 39 12 41
rect 8 37 12 39
rect 18 41 22 83
rect 18 39 19 41
rect 21 39 22 41
rect 18 37 22 39
rect 28 82 32 83
rect 28 81 68 82
rect 28 79 29 81
rect 31 79 68 81
rect 28 78 68 79
rect 28 71 32 78
rect 28 69 29 71
rect 31 69 32 71
rect 28 32 32 69
rect 15 31 32 32
rect 15 29 17 31
rect 19 29 32 31
rect 15 28 32 29
rect 38 41 42 73
rect 38 39 39 41
rect 41 39 42 41
rect 38 27 42 39
rect 48 41 52 73
rect 64 72 68 78
rect 76 81 80 88
rect 76 79 77 81
rect 79 79 80 81
rect 76 77 80 79
rect 88 81 92 83
rect 88 79 89 81
rect 91 79 92 81
rect 64 68 78 72
rect 48 39 49 41
rect 51 39 52 41
rect 48 27 52 39
rect 64 61 68 63
rect 64 59 65 61
rect 67 59 68 61
rect 64 42 68 59
rect 74 51 78 68
rect 74 49 75 51
rect 77 49 78 51
rect 74 47 78 49
rect 88 71 92 79
rect 88 69 89 71
rect 91 69 92 71
rect 88 61 92 69
rect 88 59 89 61
rect 91 59 92 61
rect 64 41 83 42
rect 64 39 79 41
rect 81 39 83 41
rect 64 38 83 39
rect 3 21 57 22
rect 3 19 5 21
rect 7 19 29 21
rect 31 19 53 21
rect 55 19 57 21
rect 3 18 57 19
rect 64 21 68 38
rect 64 19 65 21
rect 67 19 68 21
rect 64 17 68 19
rect 76 21 80 23
rect 76 19 77 21
rect 79 19 80 21
rect 76 12 80 19
rect 88 21 92 59
rect 100 81 104 88
rect 100 79 101 81
rect 103 79 104 81
rect 100 71 104 79
rect 100 69 101 71
rect 103 69 104 71
rect 100 61 104 69
rect 100 59 101 61
rect 103 59 104 61
rect 100 57 104 59
rect 88 19 89 21
rect 91 19 92 21
rect 88 17 92 19
rect 100 21 104 23
rect 100 19 101 21
rect 103 19 104 21
rect 100 12 104 19
rect -2 11 112 12
rect -2 9 41 11
rect 43 9 77 11
rect 79 9 101 11
rect 103 9 112 11
rect -2 7 112 9
rect -2 5 5 7
rect 7 5 17 7
rect 19 5 29 7
rect 31 5 53 7
rect 55 5 65 7
rect 67 5 112 7
rect -2 0 112 5
<< ptie >>
rect 3 7 33 9
rect 51 7 69 9
rect 3 5 5 7
rect 7 5 17 7
rect 19 5 29 7
rect 31 5 33 7
rect 3 3 33 5
rect 51 5 53 7
rect 55 5 65 7
rect 67 5 69 7
rect 51 3 69 5
<< ntie >>
rect 15 95 45 97
rect 15 93 17 95
rect 19 93 29 95
rect 31 93 41 95
rect 43 93 45 95
rect 63 95 69 97
rect 63 93 65 95
rect 67 93 69 95
rect 15 91 45 93
rect 63 86 69 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 15 49 25
rect 71 15 73 25
rect 83 6 85 25
rect 95 6 97 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 65 49 85
rect 71 56 73 76
rect 83 55 85 94
rect 95 55 97 94
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 75 49 77 51
rect 39 39 41 41
rect 49 39 51 41
rect 79 39 81 41
<< ndifct1 >>
rect 17 29 19 31
rect 5 19 7 21
rect 29 19 31 21
rect 53 19 55 21
rect 65 19 67 21
rect 77 19 79 21
rect 41 9 43 11
rect 77 9 79 11
rect 89 19 91 21
rect 101 19 103 21
rect 101 9 103 11
<< ntiect1 >>
rect 17 93 19 95
rect 29 93 31 95
rect 41 93 43 95
rect 65 93 67 95
<< ptiect1 >>
rect 5 5 7 7
rect 17 5 19 7
rect 29 5 31 7
rect 53 5 55 7
rect 65 5 67 7
<< pdifct1 >>
rect 5 89 7 91
rect 53 89 55 91
rect 77 89 79 91
rect 29 79 31 81
rect 29 69 31 71
rect 77 79 79 81
rect 65 59 67 61
rect 89 79 91 81
rect 89 69 91 71
rect 89 59 91 61
rect 101 89 103 91
rect 101 79 103 81
rect 101 69 103 71
rect 101 59 103 61
<< labels >>
rlabel alu1 10 60 10 60 6 i0
rlabel alu1 20 60 20 60 6 i1
rlabel alu1 40 50 40 50 6 i3
rlabel alu1 50 50 50 50 6 i2
rlabel alu1 55 6 55 6 6 vss
rlabel alu1 55 94 55 94 6 vdd
rlabel alu1 90 50 90 50 6 nq
<< end >>
