magic
tech scmos
timestamp 1199202712
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 9 35 11 38
rect 19 35 21 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 30 35
rect 19 31 26 33
rect 28 31 30 33
rect 19 29 30 31
rect 12 26 14 29
rect 19 26 21 29
rect 12 3 14 8
rect 19 3 21 8
<< ndif >>
rect 7 18 12 26
rect 5 16 12 18
rect 5 14 7 16
rect 9 14 12 16
rect 5 12 12 14
rect 7 8 12 12
rect 14 8 19 26
rect 21 19 30 26
rect 21 17 26 19
rect 28 17 30 19
rect 21 12 30 17
rect 21 10 26 12
rect 28 10 30 12
rect 21 8 30 10
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
<< alu1 >>
rect -2 64 34 72
rect 2 45 14 51
rect 2 17 6 45
rect 18 37 30 43
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 27 14 31
rect 26 33 30 37
rect 28 31 30 33
rect 26 29 30 31
rect 10 21 22 27
rect 2 16 11 17
rect 2 14 7 16
rect 9 14 11 16
rect 2 13 11 14
rect -2 0 34 8
<< nmos >>
rect 12 8 14 26
rect 19 8 21 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
<< polyct1 >>
rect 11 31 13 33
rect 26 31 28 33
<< ndifct0 >>
rect 26 17 28 19
rect 26 10 28 12
<< ndifct1 >>
rect 7 14 9 16
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 55 16 57
rect 14 48 16 50
rect 24 62 26 64
rect 24 55 26 57
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 51 17 55
rect 22 57 28 62
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 14 50 17 51
rect 16 48 17 50
rect 14 46 17 48
rect 24 30 26 37
rect 25 19 29 21
rect 25 17 26 19
rect 28 17 29 19
rect 25 12 29 17
rect 25 10 26 12
rect 28 10 29 12
rect 25 8 29 10
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 28 12 28 6 b
rlabel alu1 12 48 12 48 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 24 20 24 6 b
rlabel alu1 20 40 20 40 6 a
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 36 28 36 6 a
<< end >>
