magic
tech scmos
timestamp 1199203607
<< ab >>
rect 0 0 240 80
<< nwell >>
rect -5 36 245 88
<< pwell >>
rect -5 -8 245 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 69 41 74
rect 49 69 51 74
rect 59 69 61 74
rect 79 72 91 74
rect 79 69 81 72
rect 89 69 91 72
rect 119 69 121 74
rect 129 69 131 74
rect 139 69 141 74
rect 149 69 151 74
rect 159 69 161 74
rect 169 69 171 74
rect 179 69 181 74
rect 189 69 191 74
rect 199 69 201 74
rect 209 69 211 74
rect 219 69 221 74
rect 99 56 101 61
rect 109 56 111 61
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 37 61 39
rect 79 38 81 42
rect 89 39 91 42
rect 99 39 101 42
rect 109 39 111 42
rect 119 39 121 42
rect 129 39 131 42
rect 139 39 141 42
rect 149 39 151 42
rect 9 35 11 37
rect 13 35 61 37
rect 85 37 91 39
rect 85 35 87 37
rect 89 35 91 37
rect 9 33 61 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 59 30 61 33
rect 69 30 71 35
rect 79 30 81 34
rect 85 33 91 35
rect 95 37 115 39
rect 95 35 97 37
rect 99 35 111 37
rect 113 35 115 37
rect 95 33 115 35
rect 119 37 131 39
rect 119 35 124 37
rect 126 35 131 37
rect 119 33 131 35
rect 135 37 151 39
rect 135 35 137 37
rect 139 35 141 37
rect 135 33 141 35
rect 159 35 161 42
rect 169 39 171 42
rect 169 37 175 39
rect 169 35 171 37
rect 173 35 175 37
rect 159 33 175 35
rect 89 30 91 33
rect 96 30 98 33
rect 112 30 114 33
rect 119 30 121 33
rect 129 30 131 33
rect 136 30 138 33
rect 152 31 161 33
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 59 9 61 12
rect 69 9 71 12
rect 79 9 81 12
rect 152 29 154 31
rect 156 29 161 31
rect 172 30 174 33
rect 179 30 181 42
rect 189 39 191 42
rect 199 39 201 42
rect 209 39 211 42
rect 219 39 221 42
rect 189 37 231 39
rect 189 35 227 37
rect 229 35 231 37
rect 189 33 231 35
rect 189 30 191 33
rect 199 30 201 33
rect 209 30 211 33
rect 152 27 161 29
rect 172 12 174 16
rect 59 7 81 9
rect 89 6 91 10
rect 96 6 98 10
rect 112 6 114 10
rect 119 6 121 10
rect 129 7 131 12
rect 136 8 138 12
rect 179 8 181 16
rect 136 6 181 8
rect 189 7 191 12
rect 199 7 201 12
rect 209 7 211 12
<< ndif >>
rect 2 24 9 30
rect 2 22 4 24
rect 6 22 9 24
rect 2 16 9 22
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 12 19 19
rect 21 16 29 30
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 31 28 38 30
rect 31 26 34 28
rect 36 26 38 28
rect 31 21 38 26
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
rect 52 28 59 30
rect 52 26 54 28
rect 56 26 59 28
rect 52 21 59 26
rect 52 19 54 21
rect 56 19 59 21
rect 52 17 59 19
rect 31 12 36 17
rect 54 12 59 17
rect 61 21 69 30
rect 61 19 64 21
rect 66 19 69 21
rect 61 12 69 19
rect 71 28 79 30
rect 71 26 74 28
rect 76 26 79 28
rect 71 12 79 26
rect 81 21 89 30
rect 81 19 84 21
rect 86 19 89 21
rect 81 12 89 19
rect 84 10 89 12
rect 91 10 96 30
rect 98 14 112 30
rect 98 12 104 14
rect 106 12 112 14
rect 98 10 112 12
rect 114 10 119 30
rect 121 21 129 30
rect 121 19 124 21
rect 126 19 129 21
rect 121 12 129 19
rect 131 12 136 30
rect 138 14 147 30
rect 165 28 172 30
rect 165 26 167 28
rect 169 26 172 28
rect 165 24 172 26
rect 167 16 172 24
rect 174 16 179 30
rect 181 27 189 30
rect 181 25 184 27
rect 186 25 189 27
rect 181 20 189 25
rect 181 18 184 20
rect 186 18 189 20
rect 181 16 189 18
rect 138 12 142 14
rect 144 12 147 14
rect 121 10 126 12
rect 140 10 147 12
rect 184 12 189 16
rect 191 28 199 30
rect 191 26 194 28
rect 196 26 199 28
rect 191 21 199 26
rect 191 19 194 21
rect 196 19 199 21
rect 191 12 199 19
rect 201 24 209 30
rect 201 22 204 24
rect 206 22 209 24
rect 201 16 209 22
rect 201 14 204 16
rect 206 14 209 16
rect 201 12 209 14
rect 211 28 218 30
rect 211 26 214 28
rect 216 26 218 28
rect 211 21 218 26
rect 211 19 214 21
rect 216 19 218 21
rect 211 17 218 19
rect 211 12 216 17
<< pdif >>
rect 2 67 9 69
rect 2 65 4 67
rect 6 65 9 67
rect 2 60 9 65
rect 2 58 4 60
rect 6 58 9 60
rect 2 42 9 58
rect 11 53 19 69
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 53 39 69
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 67 49 69
rect 41 65 44 67
rect 46 65 49 67
rect 41 60 49 65
rect 41 58 44 60
rect 46 58 49 60
rect 41 42 49 58
rect 51 53 59 69
rect 51 51 54 53
rect 56 51 59 53
rect 51 46 59 51
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 67 68 69
rect 61 65 64 67
rect 66 65 68 67
rect 61 60 68 65
rect 74 62 79 69
rect 61 58 64 60
rect 66 58 68 60
rect 61 42 68 58
rect 72 60 79 62
rect 72 58 74 60
rect 76 58 79 60
rect 72 53 79 58
rect 72 51 74 53
rect 76 51 79 53
rect 72 49 79 51
rect 74 42 79 49
rect 81 53 89 69
rect 81 51 84 53
rect 86 51 89 53
rect 81 46 89 51
rect 81 44 84 46
rect 86 44 89 46
rect 81 42 89 44
rect 91 56 96 69
rect 114 56 119 69
rect 91 54 99 56
rect 91 52 94 54
rect 96 52 99 54
rect 91 42 99 52
rect 101 46 109 56
rect 101 44 104 46
rect 106 44 109 46
rect 101 42 109 44
rect 111 54 119 56
rect 111 52 114 54
rect 116 52 119 54
rect 111 42 119 52
rect 121 46 129 69
rect 121 44 124 46
rect 126 44 129 46
rect 121 42 129 44
rect 131 61 139 69
rect 131 59 134 61
rect 136 59 139 61
rect 131 42 139 59
rect 141 46 149 69
rect 141 44 144 46
rect 146 44 149 46
rect 141 42 149 44
rect 151 61 159 69
rect 151 59 154 61
rect 156 59 159 61
rect 151 42 159 59
rect 161 53 169 69
rect 161 51 164 53
rect 166 51 169 53
rect 161 42 169 51
rect 171 60 179 69
rect 171 58 174 60
rect 176 58 179 60
rect 171 53 179 58
rect 171 51 174 53
rect 176 51 179 53
rect 171 46 179 51
rect 171 44 174 46
rect 176 44 179 46
rect 171 42 179 44
rect 181 53 189 69
rect 181 51 184 53
rect 186 51 189 53
rect 181 46 189 51
rect 181 44 184 46
rect 186 44 189 46
rect 181 42 189 44
rect 191 67 199 69
rect 191 65 194 67
rect 196 65 199 67
rect 191 60 199 65
rect 191 58 194 60
rect 196 58 199 60
rect 191 42 199 58
rect 201 53 209 69
rect 201 51 204 53
rect 206 51 209 53
rect 201 46 209 51
rect 201 44 204 46
rect 206 44 209 46
rect 201 42 209 44
rect 211 67 219 69
rect 211 65 214 67
rect 216 65 219 67
rect 211 60 219 65
rect 211 58 214 60
rect 216 58 219 60
rect 211 42 219 58
rect 221 55 226 69
rect 221 53 228 55
rect 221 51 224 53
rect 226 51 228 53
rect 221 46 228 51
rect 221 44 224 46
rect 226 44 228 46
rect 221 42 228 44
<< alu1 >>
rect -2 81 242 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 203 81
rect 205 79 211 81
rect 213 79 219 81
rect 221 79 227 81
rect 229 79 235 81
rect 237 79 242 81
rect -2 68 242 79
rect 73 61 177 62
rect 73 60 134 61
rect 73 58 74 60
rect 76 59 134 60
rect 136 59 154 61
rect 156 60 177 61
rect 156 59 174 60
rect 76 58 174 59
rect 176 58 177 60
rect 2 38 6 47
rect 73 53 78 58
rect 73 51 74 53
rect 76 51 78 53
rect 73 49 78 51
rect 92 54 98 58
rect 92 52 94 54
rect 96 52 98 54
rect 92 51 98 52
rect 112 54 118 58
rect 112 52 114 54
rect 116 52 118 54
rect 112 51 118 52
rect 173 53 177 58
rect 173 51 174 53
rect 176 51 177 53
rect 2 37 15 38
rect 2 35 11 37
rect 13 35 15 37
rect 2 33 15 35
rect 173 46 177 51
rect 162 44 174 46
rect 176 44 177 46
rect 162 42 177 44
rect 162 22 166 42
rect 62 21 166 22
rect 62 19 64 21
rect 66 19 84 21
rect 86 19 124 21
rect 126 19 166 21
rect 62 18 166 19
rect 226 37 238 39
rect 226 35 227 37
rect 229 35 238 37
rect 226 33 238 35
rect 234 25 238 33
rect -2 1 242 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 203 1
rect 205 -1 211 1
rect 213 -1 219 1
rect 221 -1 227 1
rect 229 -1 235 1
rect 237 -1 242 1
rect -2 -2 242 -1
<< ptie >>
rect 0 1 240 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 203 1
rect 205 -1 211 1
rect 213 -1 219 1
rect 221 -1 227 1
rect 229 -1 235 1
rect 237 -1 240 1
rect 0 -3 240 -1
<< ntie >>
rect 0 81 240 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 203 81
rect 205 79 211 81
rect 213 79 219 81
rect 221 79 227 81
rect 229 79 235 81
rect 237 79 240 81
rect 0 77 240 79
<< nmos >>
rect 9 12 11 30
rect 19 12 21 30
rect 29 12 31 30
rect 59 12 61 30
rect 69 12 71 30
rect 79 12 81 30
rect 89 10 91 30
rect 96 10 98 30
rect 112 10 114 30
rect 119 10 121 30
rect 129 12 131 30
rect 136 12 138 30
rect 172 16 174 30
rect 179 16 181 30
rect 189 12 191 30
rect 199 12 201 30
rect 209 12 211 30
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 49 42 51 69
rect 59 42 61 69
rect 79 42 81 69
rect 89 42 91 69
rect 99 42 101 56
rect 109 42 111 56
rect 119 42 121 69
rect 129 42 131 69
rect 139 42 141 69
rect 149 42 151 69
rect 159 42 161 69
rect 169 42 171 69
rect 179 42 181 69
rect 189 42 191 69
rect 199 42 201 69
rect 209 42 211 69
rect 219 42 221 69
<< polyct0 >>
rect 87 35 89 37
rect 97 35 99 37
rect 111 35 113 37
rect 124 35 126 37
rect 137 35 139 37
rect 171 35 173 37
rect 154 29 156 31
<< polyct1 >>
rect 11 35 13 37
rect 227 35 229 37
<< ndifct0 >>
rect 4 22 6 24
rect 4 14 6 16
rect 14 26 16 28
rect 14 19 16 21
rect 24 14 26 16
rect 34 26 36 28
rect 34 19 36 21
rect 54 26 56 28
rect 54 19 56 21
rect 74 26 76 28
rect 104 12 106 14
rect 167 26 169 28
rect 184 25 186 27
rect 184 18 186 20
rect 142 12 144 14
rect 194 26 196 28
rect 194 19 196 21
rect 204 22 206 24
rect 204 14 206 16
rect 214 26 216 28
rect 214 19 216 21
<< ndifct1 >>
rect 64 19 66 21
rect 84 19 86 21
rect 124 19 126 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
rect 171 79 173 81
rect 179 79 181 81
rect 187 79 189 81
rect 195 79 197 81
rect 203 79 205 81
rect 211 79 213 81
rect 219 79 221 81
rect 227 79 229 81
rect 235 79 237 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
rect 171 -1 173 1
rect 179 -1 181 1
rect 187 -1 189 1
rect 195 -1 197 1
rect 203 -1 205 1
rect 211 -1 213 1
rect 219 -1 221 1
rect 227 -1 229 1
rect 235 -1 237 1
<< pdifct0 >>
rect 4 65 6 67
rect 4 58 6 60
rect 14 51 16 53
rect 14 44 16 46
rect 24 65 26 67
rect 24 58 26 60
rect 34 51 36 53
rect 34 44 36 46
rect 44 65 46 67
rect 44 58 46 60
rect 54 51 56 53
rect 54 44 56 46
rect 64 65 66 67
rect 64 58 66 60
rect 84 51 86 53
rect 84 44 86 46
rect 104 44 106 46
rect 124 44 126 46
rect 144 44 146 46
rect 164 51 166 53
rect 184 51 186 53
rect 184 44 186 46
rect 194 65 196 67
rect 194 58 196 60
rect 204 51 206 53
rect 204 44 206 46
rect 214 65 216 67
rect 214 58 216 60
rect 224 51 226 53
rect 224 44 226 46
<< pdifct1 >>
rect 74 58 76 60
rect 74 51 76 53
rect 94 52 96 54
rect 114 52 116 54
rect 134 59 136 61
rect 154 59 156 61
rect 174 58 176 60
rect 174 51 176 53
rect 174 44 176 46
<< alu0 >>
rect 3 67 7 68
rect 3 65 4 67
rect 6 65 7 67
rect 3 60 7 65
rect 3 58 4 60
rect 6 58 7 60
rect 3 56 7 58
rect 23 67 27 68
rect 23 65 24 67
rect 26 65 27 67
rect 23 60 27 65
rect 23 58 24 60
rect 26 58 27 60
rect 23 56 27 58
rect 43 67 47 68
rect 43 65 44 67
rect 46 65 47 67
rect 43 60 47 65
rect 43 58 44 60
rect 46 58 47 60
rect 43 56 47 58
rect 63 67 67 68
rect 63 65 64 67
rect 66 65 67 67
rect 63 60 67 65
rect 193 67 197 68
rect 193 65 194 67
rect 196 65 197 67
rect 63 58 64 60
rect 66 58 67 60
rect 63 56 67 58
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 13 46 17 51
rect 33 53 37 55
rect 33 51 34 53
rect 36 51 37 53
rect 33 46 37 51
rect 53 53 57 55
rect 53 51 54 53
rect 56 51 57 53
rect 53 46 57 51
rect 83 53 87 55
rect 83 51 84 53
rect 86 51 87 53
rect 134 53 168 54
rect 134 51 164 53
rect 166 51 168 53
rect 83 46 87 51
rect 134 50 168 51
rect 193 60 197 65
rect 193 58 194 60
rect 196 58 197 60
rect 193 56 197 58
rect 213 67 217 68
rect 213 65 214 67
rect 216 65 217 67
rect 213 60 217 65
rect 213 58 214 60
rect 216 58 217 60
rect 213 56 217 58
rect 103 46 107 48
rect 134 47 138 50
rect 13 44 14 46
rect 16 44 34 46
rect 36 44 54 46
rect 56 44 84 46
rect 86 44 100 46
rect 13 42 100 44
rect 33 29 37 42
rect 86 37 90 39
rect 86 35 87 37
rect 89 35 90 37
rect 86 30 90 35
rect 96 37 100 42
rect 96 35 97 37
rect 99 35 100 37
rect 96 33 100 35
rect 103 44 104 46
rect 106 44 107 46
rect 103 30 107 44
rect 110 46 138 47
rect 110 44 124 46
rect 126 44 138 46
rect 110 43 138 44
rect 142 46 149 47
rect 142 44 144 46
rect 146 44 149 46
rect 142 43 149 44
rect 110 37 114 43
rect 134 38 138 43
rect 110 35 111 37
rect 113 35 114 37
rect 110 33 114 35
rect 122 37 128 38
rect 122 35 124 37
rect 126 35 128 37
rect 122 30 128 35
rect 134 37 141 38
rect 134 35 137 37
rect 139 35 141 37
rect 134 34 141 35
rect 145 32 149 43
rect 183 53 187 55
rect 183 51 184 53
rect 186 51 187 53
rect 183 47 187 51
rect 203 53 207 55
rect 203 51 204 53
rect 206 51 207 53
rect 203 47 207 51
rect 223 53 228 55
rect 223 51 224 53
rect 226 51 228 53
rect 223 47 228 51
rect 183 46 228 47
rect 183 44 184 46
rect 186 44 204 46
rect 206 44 224 46
rect 226 44 228 46
rect 183 43 228 44
rect 145 31 158 32
rect 145 30 154 31
rect 12 28 37 29
rect 12 26 14 28
rect 16 26 34 28
rect 36 26 37 28
rect 3 24 7 26
rect 3 22 4 24
rect 6 22 7 24
rect 3 16 7 22
rect 12 25 37 26
rect 12 21 17 25
rect 12 19 14 21
rect 16 19 17 21
rect 12 17 17 19
rect 33 21 37 25
rect 33 19 34 21
rect 36 19 37 21
rect 3 14 4 16
rect 6 14 7 16
rect 3 12 7 14
rect 23 16 27 18
rect 33 17 37 19
rect 53 29 154 30
rect 156 29 158 31
rect 53 28 158 29
rect 53 26 54 28
rect 56 26 74 28
rect 76 26 149 28
rect 53 21 57 26
rect 72 25 78 26
rect 183 38 187 43
rect 169 37 187 38
rect 169 35 171 37
rect 173 35 187 37
rect 169 34 187 35
rect 166 28 171 29
rect 166 26 167 28
rect 169 26 171 28
rect 166 25 171 26
rect 183 27 187 29
rect 183 25 184 27
rect 186 25 187 27
rect 53 19 54 21
rect 56 19 57 21
rect 53 17 57 19
rect 183 20 187 25
rect 183 18 184 20
rect 186 18 187 20
rect 23 14 24 16
rect 26 14 27 16
rect 23 12 27 14
rect 102 14 108 15
rect 102 12 104 14
rect 106 12 108 14
rect 140 14 146 15
rect 140 12 142 14
rect 144 12 146 14
rect 155 12 161 15
rect 183 12 187 18
rect 193 28 197 43
rect 193 26 194 28
rect 196 26 197 28
rect 213 28 217 43
rect 213 26 214 28
rect 216 26 217 28
rect 193 21 197 26
rect 193 19 194 21
rect 196 19 197 21
rect 193 17 197 19
rect 203 24 207 26
rect 203 22 204 24
rect 206 22 207 24
rect 203 16 207 22
rect 213 21 217 26
rect 213 19 214 21
rect 216 19 217 21
rect 213 17 217 19
rect 203 14 204 16
rect 206 14 207 16
rect 203 12 207 14
<< labels >>
rlabel alu0 14 23 14 23 6 bn
rlabel alu0 15 48 15 48 6 bn
rlabel alu0 35 36 35 36 6 bn
rlabel alu0 55 23 55 23 6 an
rlabel alu0 88 32 88 32 6 an
rlabel alu0 85 48 85 48 6 bn
rlabel alu0 55 48 55 48 6 bn
rlabel alu0 125 32 125 32 6 an
rlabel alu0 112 40 112 40 6 bn
rlabel alu0 98 39 98 39 6 bn
rlabel alu0 124 45 124 45 6 bn
rlabel alu0 136 44 136 44 6 bn
rlabel alu0 105 37 105 37 6 an
rlabel alu0 101 28 101 28 6 an
rlabel alu0 151 30 151 30 6 an
rlabel pdifct0 145 45 145 45 6 an
rlabel alu0 178 36 178 36 6 an
rlabel alu0 151 52 151 52 6 bn
rlabel alu0 215 32 215 32 6 an
rlabel alu0 195 32 195 32 6 an
rlabel pdifct0 205 45 205 45 6 an
rlabel alu0 205 49 205 49 6 an
rlabel alu0 225 49 225 49 6 an
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 40 4 40 6 b
rlabel alu1 92 20 92 20 6 z
rlabel alu1 84 20 84 20 6 z
rlabel alu1 76 20 76 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 92 60 92 60 6 z
rlabel alu1 84 60 84 60 6 z
rlabel alu1 76 56 76 56 6 z
rlabel alu1 120 6 120 6 6 vss
rlabel alu1 100 20 100 20 6 z
rlabel alu1 108 20 108 20 6 z
rlabel alu1 116 20 116 20 6 z
rlabel alu1 124 20 124 20 6 z
rlabel alu1 132 20 132 20 6 z
rlabel alu1 140 20 140 20 6 z
rlabel alu1 140 60 140 60 6 z
rlabel alu1 132 60 132 60 6 z
rlabel alu1 124 60 124 60 6 z
rlabel alu1 116 60 116 60 6 z
rlabel alu1 108 60 108 60 6 z
rlabel alu1 100 60 100 60 6 z
rlabel alu1 120 74 120 74 6 vdd
rlabel alu1 148 20 148 20 6 z
rlabel alu1 156 20 156 20 6 z
rlabel alu1 164 32 164 32 6 z
rlabel alu1 172 44 172 44 6 z
rlabel alu1 148 60 148 60 6 z
rlabel alu1 172 60 172 60 6 z
rlabel alu1 164 60 164 60 6 z
rlabel alu1 156 60 156 60 6 z
rlabel alu1 236 32 236 32 6 a
rlabel polyct1 228 36 228 36 6 a
<< end >>
