magic
tech scmos
timestamp 1199203053
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 14 69 16 74
rect 21 69 23 74
rect 28 69 30 74
rect 35 69 37 74
rect 47 69 49 74
rect 54 69 56 74
rect 61 69 63 74
rect 68 69 70 74
rect 78 69 80 74
rect 85 69 87 74
rect 92 69 94 74
rect 99 69 101 74
rect 14 41 16 44
rect 9 39 16 41
rect 9 37 11 39
rect 13 37 16 39
rect 9 35 16 37
rect 10 22 12 35
rect 21 31 23 44
rect 17 29 23 31
rect 17 27 19 29
rect 21 27 23 29
rect 17 25 23 27
rect 28 31 30 44
rect 35 39 37 44
rect 47 39 49 42
rect 35 37 49 39
rect 38 35 40 37
rect 42 35 44 37
rect 38 33 44 35
rect 28 29 34 31
rect 28 27 30 29
rect 32 27 34 29
rect 28 25 34 27
rect 20 22 22 25
rect 32 22 34 25
rect 42 22 44 33
rect 54 31 56 42
rect 61 33 63 42
rect 68 39 70 42
rect 78 39 80 42
rect 68 37 81 39
rect 75 35 77 37
rect 79 35 81 37
rect 75 33 81 35
rect 61 31 71 33
rect 48 29 56 31
rect 48 27 50 29
rect 52 27 56 29
rect 65 29 67 31
rect 69 29 71 31
rect 85 29 87 42
rect 65 27 87 29
rect 48 25 56 27
rect 54 23 56 25
rect 92 23 94 42
rect 54 21 94 23
rect 99 23 101 42
rect 99 21 105 23
rect 99 19 101 21
rect 103 19 105 21
rect 99 17 105 19
rect 10 6 12 11
rect 20 6 22 11
rect 32 6 34 11
rect 42 6 44 11
<< ndif >>
rect 2 11 10 22
rect 12 20 20 22
rect 12 18 15 20
rect 17 18 20 20
rect 12 11 20 18
rect 22 11 32 22
rect 34 20 42 22
rect 34 18 37 20
rect 39 18 42 20
rect 34 11 42 18
rect 44 11 52 22
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
rect 24 9 26 11
rect 28 9 30 11
rect 24 7 30 9
rect 46 9 48 11
rect 50 9 52 11
rect 46 7 52 9
<< pdif >>
rect 39 71 45 73
rect 39 69 41 71
rect 43 69 45 71
rect 9 63 14 69
rect 7 61 14 63
rect 7 59 9 61
rect 11 59 14 61
rect 7 57 14 59
rect 9 44 14 57
rect 16 44 21 69
rect 23 44 28 69
rect 30 44 35 69
rect 37 44 47 69
rect 39 42 47 44
rect 49 42 54 69
rect 56 42 61 69
rect 63 42 68 69
rect 70 61 78 69
rect 70 59 73 61
rect 75 59 78 61
rect 70 42 78 59
rect 80 42 85 69
rect 87 42 92 69
rect 94 42 99 69
rect 101 67 108 69
rect 101 65 104 67
rect 106 65 108 67
rect 101 60 108 65
rect 101 58 104 60
rect 106 58 108 60
rect 101 42 108 58
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 71 114 79
rect -2 69 41 71
rect 43 69 114 71
rect -2 68 114 69
rect 2 61 79 62
rect 2 59 9 61
rect 11 59 73 61
rect 75 59 79 61
rect 2 58 79 59
rect 2 23 6 58
rect 10 50 80 54
rect 10 39 14 50
rect 10 37 11 39
rect 13 37 14 39
rect 10 33 14 37
rect 18 42 70 46
rect 18 29 22 42
rect 38 37 62 38
rect 38 35 40 37
rect 42 35 62 37
rect 38 34 62 35
rect 18 27 19 29
rect 21 27 22 29
rect 18 25 22 27
rect 28 29 54 30
rect 28 27 30 29
rect 32 27 50 29
rect 52 27 54 29
rect 28 26 54 27
rect 2 21 14 23
rect 33 21 41 22
rect 2 20 41 21
rect 2 18 15 20
rect 17 18 37 20
rect 39 18 41 20
rect 2 17 41 18
rect 50 17 54 26
rect 58 22 62 34
rect 66 31 70 42
rect 74 37 80 50
rect 74 35 77 37
rect 79 35 80 37
rect 74 33 80 35
rect 66 29 67 31
rect 69 29 70 31
rect 66 27 70 29
rect 58 21 105 22
rect 58 19 101 21
rect 103 19 105 21
rect 58 18 105 19
rect -2 11 114 12
rect -2 9 4 11
rect 6 9 26 11
rect 28 9 48 11
rect 50 9 114 11
rect -2 1 114 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 10 11 12 22
rect 20 11 22 22
rect 32 11 34 22
rect 42 11 44 22
<< pmos >>
rect 14 44 16 69
rect 21 44 23 69
rect 28 44 30 69
rect 35 44 37 69
rect 47 42 49 69
rect 54 42 56 69
rect 61 42 63 69
rect 68 42 70 69
rect 78 42 80 69
rect 85 42 87 69
rect 92 42 94 69
rect 99 42 101 69
<< polyct1 >>
rect 11 37 13 39
rect 19 27 21 29
rect 40 35 42 37
rect 30 27 32 29
rect 77 35 79 37
rect 50 27 52 29
rect 67 29 69 31
rect 101 19 103 21
<< ndifct1 >>
rect 15 18 17 20
rect 37 18 39 20
rect 4 9 6 11
rect 26 9 28 11
rect 48 9 50 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 104 65 106 67
rect 104 58 106 60
<< pdifct1 >>
rect 41 69 43 71
rect 9 59 11 61
rect 73 59 75 61
<< alu0 >>
rect 102 67 108 68
rect 102 65 104 67
rect 106 65 108 67
rect 102 60 108 65
rect 102 58 104 60
rect 106 58 108 60
rect 102 57 108 58
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 40 12 40 6 d
rlabel alu1 12 60 12 60 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 b
rlabel alu1 20 32 20 32 6 c
rlabel alu1 28 44 28 44 6 c
rlabel alu1 36 44 36 44 6 c
rlabel alu1 28 52 28 52 6 d
rlabel alu1 36 52 36 52 6 d
rlabel alu1 20 52 20 52 6 d
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 56 6 56 6 6 vss
rlabel alu1 44 28 44 28 6 b
rlabel alu1 52 20 52 20 6 b
rlabel alu1 60 28 60 28 6 a
rlabel alu1 44 36 44 36 6 a
rlabel alu1 44 44 44 44 6 c
rlabel alu1 52 36 52 36 6 a
rlabel alu1 52 44 52 44 6 c
rlabel alu1 60 44 60 44 6 c
rlabel alu1 52 52 52 52 6 d
rlabel alu1 60 52 60 52 6 d
rlabel alu1 44 52 44 52 6 d
rlabel alu1 44 60 44 60 6 z
rlabel alu1 52 60 52 60 6 z
rlabel alu1 60 60 60 60 6 z
rlabel alu1 56 74 56 74 6 vdd
rlabel alu1 68 20 68 20 6 a
rlabel alu1 76 20 76 20 6 a
rlabel alu1 84 20 84 20 6 a
rlabel alu1 68 36 68 36 6 c
rlabel alu1 76 44 76 44 6 d
rlabel alu1 68 52 68 52 6 d
rlabel alu1 68 60 68 60 6 z
rlabel alu1 76 60 76 60 6 z
rlabel alu1 92 20 92 20 6 a
rlabel alu1 100 20 100 20 6 a
<< end >>
