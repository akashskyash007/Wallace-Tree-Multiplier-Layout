magic
tech scmos
timestamp 1199202957
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 12 69 14 74
rect 19 69 21 74
rect 29 69 31 74
rect 36 69 38 74
rect 12 39 14 42
rect 19 39 21 42
rect 29 39 31 42
rect 36 39 38 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 32 39
rect 19 35 28 37
rect 30 35 32 37
rect 19 33 32 35
rect 36 37 49 39
rect 36 35 45 37
rect 47 35 49 37
rect 36 33 49 35
rect 9 23 11 33
rect 19 23 21 33
rect 29 23 31 33
rect 39 30 41 33
rect 39 12 41 17
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
<< ndif >>
rect 34 23 39 30
rect 2 14 9 23
rect 2 12 4 14
rect 6 12 9 14
rect 2 10 9 12
rect 11 21 19 23
rect 11 19 14 21
rect 16 19 19 21
rect 11 10 19 19
rect 21 14 29 23
rect 21 12 24 14
rect 26 12 29 14
rect 21 10 29 12
rect 31 21 39 23
rect 31 19 34 21
rect 36 19 39 21
rect 31 17 39 19
rect 41 21 49 30
rect 41 19 44 21
rect 46 19 49 21
rect 41 17 49 19
rect 31 10 36 17
<< pdif >>
rect 4 67 12 69
rect 4 65 7 67
rect 9 65 12 67
rect 4 59 12 65
rect 4 57 7 59
rect 9 57 12 59
rect 4 42 12 57
rect 14 42 19 69
rect 21 53 29 69
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 42 36 69
rect 38 63 43 69
rect 38 61 46 63
rect 38 59 41 61
rect 43 59 46 61
rect 38 54 46 59
rect 38 52 41 54
rect 43 52 46 54
rect 38 42 46 52
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 22 53 31 54
rect 22 51 24 53
rect 26 51 31 53
rect 22 50 31 51
rect 22 47 28 50
rect 2 46 28 47
rect 2 44 24 46
rect 26 44 28 46
rect 2 43 28 44
rect 2 22 6 43
rect 33 42 47 46
rect 10 37 22 39
rect 33 38 39 42
rect 10 35 11 37
rect 13 35 22 37
rect 10 33 22 35
rect 26 37 39 38
rect 26 35 28 37
rect 30 35 39 37
rect 26 34 39 35
rect 43 37 49 38
rect 43 35 45 37
rect 47 35 49 37
rect 17 30 22 33
rect 43 30 49 35
rect 17 26 49 30
rect 2 21 39 22
rect 2 19 14 21
rect 16 19 34 21
rect 36 19 39 21
rect 2 18 39 19
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 10 11 23
rect 19 10 21 23
rect 29 10 31 23
rect 39 17 41 30
<< pmos >>
rect 12 42 14 69
rect 19 42 21 69
rect 29 42 31 69
rect 36 42 38 69
<< polyct1 >>
rect 11 35 13 37
rect 28 35 30 37
rect 45 35 47 37
<< ndifct0 >>
rect 4 12 6 14
rect 24 12 26 14
rect 44 19 46 21
<< ndifct1 >>
rect 14 19 16 21
rect 34 19 36 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 7 65 9 67
rect 7 57 9 59
rect 41 59 43 61
rect 41 52 43 54
<< pdifct1 >>
rect 24 51 26 53
rect 24 44 26 46
<< alu0 >>
rect 6 67 10 68
rect 6 65 7 67
rect 9 65 10 67
rect 6 59 10 65
rect 6 57 7 59
rect 9 57 10 59
rect 6 55 10 57
rect 40 61 44 68
rect 40 59 41 61
rect 43 59 44 61
rect 40 54 44 59
rect 40 52 41 54
rect 43 52 44 54
rect 40 50 44 52
rect 43 21 47 23
rect 43 19 44 21
rect 46 19 47 21
rect 2 14 8 15
rect 2 12 4 14
rect 6 12 8 14
rect 22 14 28 15
rect 22 12 24 14
rect 26 12 28 14
rect 43 12 47 19
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 32 20 32 6 a
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 40 36 40 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 44 44 44 6 b
<< end >>
