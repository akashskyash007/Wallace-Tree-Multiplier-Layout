magic
tech scmos
timestamp 1199203200
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 39 69 41 74
rect 46 69 48 74
rect 29 62 31 67
rect 9 54 11 59
rect 29 47 31 54
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 9 39 11 42
rect 29 41 35 43
rect 9 37 18 39
rect 9 35 14 37
rect 16 35 18 37
rect 9 33 18 35
rect 9 30 11 33
rect 29 30 31 41
rect 39 39 41 54
rect 46 47 48 54
rect 46 45 57 47
rect 51 43 53 45
rect 55 43 57 45
rect 51 41 57 43
rect 39 37 47 39
rect 39 35 43 37
rect 45 35 47 37
rect 39 33 47 35
rect 39 30 41 33
rect 9 19 11 24
rect 51 23 53 41
rect 29 18 31 23
rect 39 18 41 23
rect 51 11 53 16
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 11 28 18 30
rect 11 26 14 28
rect 16 26 18 28
rect 11 24 18 26
rect 22 28 29 30
rect 22 26 24 28
rect 26 26 29 28
rect 22 23 29 26
rect 31 27 39 30
rect 31 25 34 27
rect 36 25 39 27
rect 31 23 39 25
rect 41 23 49 30
rect 43 16 51 23
rect 53 20 60 23
rect 53 18 56 20
rect 58 18 60 20
rect 53 16 60 18
rect 43 11 49 16
rect 43 9 45 11
rect 47 9 49 11
rect 43 7 49 9
<< pdif >>
rect 13 62 27 64
rect 34 62 39 69
rect 13 60 15 62
rect 17 60 29 62
rect 13 54 29 60
rect 31 60 39 62
rect 31 58 34 60
rect 36 58 39 60
rect 31 54 39 58
rect 41 54 46 69
rect 48 67 56 69
rect 48 65 51 67
rect 53 65 56 67
rect 48 60 56 65
rect 48 58 51 60
rect 53 58 56 60
rect 48 54 56 58
rect 4 48 9 54
rect 2 46 9 48
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 52 15 54
rect 17 52 27 54
rect 11 42 27 52
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 46 15 47
rect 2 44 4 46
rect 6 44 15 46
rect 2 42 15 44
rect 2 30 6 42
rect 42 50 46 55
rect 34 47 46 50
rect 30 46 46 47
rect 30 45 38 46
rect 30 43 31 45
rect 33 43 38 45
rect 30 41 38 43
rect 50 45 62 47
rect 50 43 53 45
rect 55 43 62 45
rect 50 41 62 43
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 24 7 26
rect 2 17 6 24
rect 42 37 46 39
rect 42 35 43 37
rect 45 35 46 37
rect 42 31 46 35
rect 58 33 62 41
rect 42 25 54 31
rect -2 11 66 12
rect -2 9 45 11
rect 47 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 24 11 30
rect 29 23 31 30
rect 39 23 41 30
rect 51 16 53 23
<< pmos >>
rect 29 54 31 62
rect 39 54 41 69
rect 46 54 48 69
rect 9 42 11 54
<< polyct0 >>
rect 14 35 16 37
<< polyct1 >>
rect 31 43 33 45
rect 53 43 55 45
rect 43 35 45 37
<< ndifct0 >>
rect 14 26 16 28
rect 24 26 26 28
rect 34 25 36 27
rect 56 18 58 20
<< ndifct1 >>
rect 4 26 6 28
rect 45 9 47 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 15 60 17 62
rect 34 58 36 60
rect 51 65 53 67
rect 51 58 53 60
rect 15 52 17 54
<< pdifct1 >>
rect 4 44 6 46
<< alu0 >>
rect 13 62 19 68
rect 13 60 15 62
rect 17 60 19 62
rect 50 67 54 68
rect 50 65 51 67
rect 53 65 54 67
rect 13 54 19 60
rect 13 52 15 54
rect 17 52 19 54
rect 13 51 19 52
rect 23 60 38 61
rect 23 58 34 60
rect 36 58 38 60
rect 23 57 38 58
rect 50 60 54 65
rect 50 58 51 60
rect 53 58 54 60
rect 23 38 27 57
rect 50 56 54 58
rect 12 37 27 38
rect 12 35 14 37
rect 16 35 27 37
rect 12 34 27 35
rect 13 28 17 30
rect 13 26 14 28
rect 16 26 17 28
rect 13 12 17 26
rect 23 28 27 34
rect 23 26 24 28
rect 26 26 27 28
rect 23 24 27 26
rect 33 27 37 29
rect 33 25 34 27
rect 36 25 37 27
rect 33 21 37 25
rect 33 20 60 21
rect 33 18 56 20
rect 58 18 60 20
rect 33 17 60 18
<< labels >>
rlabel alu0 19 36 19 36 6 zn
rlabel alu0 25 42 25 42 6 zn
rlabel alu0 35 23 35 23 6 n1
rlabel alu0 30 59 30 59 6 zn
rlabel alu0 46 19 46 19 6 n1
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 32 44 32 6 a2
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 52 44 52 6 b
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 a2
rlabel alu1 60 40 60 40 6 a1
rlabel alu1 52 44 52 44 6 a1
<< end >>
