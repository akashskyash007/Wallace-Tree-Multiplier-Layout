magic
tech scmos
timestamp 1199203097
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 12 66 14 71
rect 22 66 24 71
rect 29 66 31 71
rect 12 55 14 58
rect 9 53 15 55
rect 9 51 11 53
rect 13 51 15 53
rect 9 49 15 51
rect 40 60 42 65
rect 9 30 11 49
rect 22 39 24 50
rect 29 47 31 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 40 46 42 50
rect 40 44 57 46
rect 29 41 35 43
rect 51 42 53 44
rect 55 42 57 44
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 19 30 21 33
rect 9 18 11 23
rect 19 18 21 23
rect 31 22 33 41
rect 51 40 57 42
rect 51 30 53 40
rect 51 19 53 24
rect 31 10 33 15
<< ndif >>
rect 2 27 9 30
rect 2 25 4 27
rect 6 25 9 27
rect 2 23 9 25
rect 11 27 19 30
rect 11 25 14 27
rect 16 25 19 27
rect 11 23 19 25
rect 21 23 29 30
rect 23 22 29 23
rect 44 28 51 30
rect 44 26 46 28
rect 48 26 51 28
rect 44 24 51 26
rect 53 28 60 30
rect 53 26 56 28
rect 58 26 60 28
rect 53 24 60 26
rect 23 15 31 22
rect 33 20 40 22
rect 33 18 36 20
rect 38 18 40 20
rect 33 15 40 18
rect 23 11 29 15
rect 23 9 25 11
rect 27 9 29 11
rect 23 7 29 9
<< pdif >>
rect 3 71 10 73
rect 3 69 6 71
rect 8 69 10 71
rect 3 66 10 69
rect 3 58 12 66
rect 14 62 22 66
rect 14 60 17 62
rect 19 60 22 62
rect 14 58 22 60
rect 17 50 22 58
rect 24 50 29 66
rect 31 61 38 66
rect 31 59 34 61
rect 36 60 38 61
rect 36 59 40 60
rect 31 50 40 59
rect 42 56 47 60
rect 42 54 49 56
rect 42 52 45 54
rect 47 52 49 54
rect 42 50 49 52
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 6 71
rect 8 69 66 71
rect -2 68 66 69
rect 2 62 23 63
rect 2 60 17 62
rect 19 60 23 62
rect 2 58 23 60
rect 2 27 6 58
rect 10 45 35 46
rect 10 43 31 45
rect 33 43 35 45
rect 10 42 35 43
rect 10 33 14 42
rect 19 37 38 38
rect 19 35 21 37
rect 23 35 38 37
rect 19 34 38 35
rect 2 25 4 27
rect 2 17 6 25
rect 34 25 38 34
rect 58 47 62 55
rect 50 44 62 47
rect 50 42 53 44
rect 55 42 62 44
rect 50 41 62 42
rect -2 11 66 12
rect -2 9 25 11
rect 27 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 23 11 30
rect 19 23 21 30
rect 51 24 53 30
rect 31 15 33 22
<< pmos >>
rect 12 58 14 66
rect 22 50 24 66
rect 29 50 31 66
rect 40 50 42 60
<< polyct0 >>
rect 11 51 13 53
<< polyct1 >>
rect 31 43 33 45
rect 53 42 55 44
rect 21 35 23 37
<< ndifct0 >>
rect 14 25 16 27
rect 46 26 48 28
rect 56 26 58 28
rect 36 18 38 20
<< ndifct1 >>
rect 4 25 6 27
rect 25 9 27 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 34 59 36 61
rect 45 52 47 54
<< pdifct1 >>
rect 6 69 8 71
rect 17 60 19 62
<< alu0 >>
rect 32 61 38 68
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 42 54 49 55
rect 9 53 45 54
rect 9 51 11 53
rect 13 52 45 53
rect 47 52 49 54
rect 13 51 49 52
rect 9 50 46 51
rect 6 23 7 29
rect 13 27 17 29
rect 13 25 14 27
rect 16 25 17 27
rect 42 29 46 50
rect 42 28 50 29
rect 42 26 46 28
rect 48 26 50 28
rect 42 25 50 26
rect 55 28 59 30
rect 55 26 56 28
rect 58 26 59 28
rect 13 21 17 25
rect 13 20 40 21
rect 13 18 36 20
rect 38 18 40 20
rect 13 17 40 18
rect 55 12 59 26
<< labels >>
rlabel alu0 15 23 15 23 6 n1
rlabel alu0 26 19 26 19 6 n1
rlabel alu0 27 52 27 52 6 bn
rlabel alu0 46 27 46 27 6 bn
rlabel alu0 45 53 45 53 6 bn
rlabel alu1 12 36 12 36 6 a1
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 36 28 36 6 a2
rlabel alu1 28 44 28 44 6 a1
rlabel alu1 20 44 20 44 6 a1
rlabel alu1 20 60 20 60 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 44 52 44 6 b
rlabel alu1 60 48 60 48 6 b
<< end >>
