magic
tech scmos
timestamp 1199202332
<< ab >>
rect 0 0 24 72
<< nwell >>
rect -5 32 29 77
<< pwell >>
rect -5 -5 29 32
<< poly >>
rect 9 62 11 67
rect 9 35 11 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 9 25 11 29
rect 9 14 11 19
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 19 19 25
rect 13 17 19 19
rect 13 15 15 17
rect 17 15 19 17
rect 13 13 19 15
<< pdif >>
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 38 9 58
rect 11 51 16 62
rect 11 49 18 51
rect 11 47 14 49
rect 16 47 18 49
rect 11 42 18 47
rect 11 40 14 42
rect 16 40 18 42
rect 11 38 18 40
<< alu1 >>
rect -2 64 26 72
rect 2 49 22 51
rect 2 47 14 49
rect 16 47 22 49
rect 2 45 22 47
rect 2 25 6 45
rect 10 33 22 35
rect 10 31 11 33
rect 13 31 22 33
rect 10 29 22 31
rect 2 23 7 25
rect 2 21 4 23
rect 6 21 7 23
rect 18 21 22 29
rect 2 19 7 21
rect -2 7 26 8
rect -2 5 5 7
rect 7 5 14 7
rect 16 5 26 7
rect -2 0 26 5
<< ptie >>
rect 3 7 18 9
rect 3 5 5 7
rect 7 5 14 7
rect 16 5 18 7
rect 3 3 18 5
<< nmos >>
rect 9 19 11 25
<< pmos >>
rect 9 38 11 62
<< polyct1 >>
rect 11 31 13 33
<< ndifct0 >>
rect 15 15 17 17
<< ndifct1 >>
rect 4 21 6 23
<< ptiect1 >>
rect 5 5 7 7
rect 14 5 16 7
<< pdifct0 >>
rect 4 58 6 60
rect 14 40 16 42
<< pdifct1 >>
rect 14 47 16 49
<< alu0 >>
rect 3 60 7 64
rect 3 58 4 60
rect 6 58 7 60
rect 3 56 7 58
rect 13 42 17 45
rect 13 40 14 42
rect 16 40 17 42
rect 13 38 17 40
rect 13 17 19 18
rect 13 15 15 17
rect 17 15 19 17
rect 13 8 19 15
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 4 12 4 6 vss
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 12 48 12 48 6 z
rlabel alu1 12 68 12 68 6 vdd
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 48 20 48 6 z
<< end >>
