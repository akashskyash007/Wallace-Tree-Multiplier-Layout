magic
tech scmos
timestamp 1199201773
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 57 11 61
rect 20 60 22 65
rect 30 60 32 65
rect 42 60 44 65
rect 52 60 54 65
rect 9 35 11 39
rect 20 35 22 54
rect 30 43 32 54
rect 42 43 44 54
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 29 37 35 39
rect 42 41 48 43
rect 42 39 44 41
rect 46 39 48 41
rect 42 37 48 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 9 21 11 29
rect 22 21 24 29
rect 29 21 31 37
rect 42 32 44 37
rect 36 30 44 32
rect 52 35 54 54
rect 52 33 58 35
rect 52 31 54 33
rect 56 31 58 33
rect 36 21 38 30
rect 52 29 58 31
rect 52 26 54 29
rect 43 24 54 26
rect 43 21 45 24
rect 9 7 11 12
rect 22 8 24 13
rect 29 8 31 13
rect 36 8 38 13
rect 43 8 45 13
<< ndif >>
rect 4 18 9 21
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 13 22 21
rect 24 13 29 21
rect 31 13 36 21
rect 38 13 43 21
rect 45 19 50 21
rect 45 17 52 19
rect 45 15 48 17
rect 50 15 52 17
rect 45 13 52 15
rect 11 12 20 13
rect 13 7 20 12
rect 13 5 15 7
rect 17 5 20 7
rect 13 3 20 5
<< pdif >>
rect 34 67 40 69
rect 34 65 36 67
rect 38 65 40 67
rect 34 60 40 65
rect 13 58 20 60
rect 13 57 15 58
rect 4 52 9 57
rect 2 50 9 52
rect 2 48 4 50
rect 6 48 9 50
rect 2 43 9 48
rect 2 41 4 43
rect 6 41 9 43
rect 2 39 9 41
rect 11 56 15 57
rect 17 56 20 58
rect 11 54 20 56
rect 22 58 30 60
rect 22 56 25 58
rect 27 56 30 58
rect 22 54 30 56
rect 32 54 42 60
rect 44 58 52 60
rect 44 56 47 58
rect 49 56 52 58
rect 44 54 52 56
rect 54 58 61 60
rect 54 56 57 58
rect 59 56 61 58
rect 54 54 61 56
rect 11 39 18 54
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 36 67
rect 38 65 66 67
rect -2 64 66 65
rect 2 50 7 59
rect 2 48 4 50
rect 6 48 7 50
rect 2 43 7 48
rect 2 41 4 43
rect 6 41 7 43
rect 2 39 7 41
rect 33 46 47 50
rect 2 18 6 39
rect 33 42 37 46
rect 58 42 62 51
rect 25 41 37 42
rect 25 39 31 41
rect 33 39 37 41
rect 25 38 37 39
rect 41 41 62 42
rect 41 39 44 41
rect 46 39 62 41
rect 41 38 62 39
rect 19 33 31 34
rect 19 31 21 33
rect 23 31 31 33
rect 19 30 31 31
rect 41 33 62 34
rect 41 31 54 33
rect 56 31 62 33
rect 41 30 62 31
rect 27 26 31 30
rect 27 22 47 26
rect 2 16 15 18
rect 2 14 4 16
rect 6 14 15 16
rect 2 13 15 14
rect 58 13 62 30
rect -2 7 66 8
rect -2 5 15 7
rect 17 5 58 7
rect 60 5 66 7
rect -2 0 66 5
<< ptie >>
rect 56 7 62 24
rect 56 5 58 7
rect 60 5 62 7
rect 56 3 62 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 12 11 21
rect 22 13 24 21
rect 29 13 31 21
rect 36 13 38 21
rect 43 13 45 21
<< pmos >>
rect 9 39 11 57
rect 20 54 22 60
rect 30 54 32 60
rect 42 54 44 60
rect 52 54 54 60
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 31 39 33 41
rect 44 39 46 41
rect 21 31 23 33
rect 54 31 56 33
<< ndifct0 >>
rect 48 15 50 17
<< ndifct1 >>
rect 4 14 6 16
rect 15 5 17 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 58 5 60 7
<< pdifct0 >>
rect 15 56 17 58
rect 25 56 27 58
rect 47 56 49 58
rect 57 56 59 58
<< pdifct1 >>
rect 36 65 38 67
rect 4 48 6 50
rect 4 41 6 43
<< alu0 >>
rect 14 58 18 64
rect 14 56 15 58
rect 17 56 18 58
rect 14 54 18 56
rect 23 58 51 59
rect 23 56 25 58
rect 27 56 47 58
rect 49 56 51 58
rect 23 55 51 56
rect 55 58 61 64
rect 55 56 57 58
rect 59 56 61 58
rect 55 55 61 56
rect 23 50 27 55
rect 11 46 27 50
rect 11 35 15 46
rect 10 33 15 35
rect 10 31 11 33
rect 13 31 15 33
rect 10 29 15 31
rect 11 26 15 29
rect 11 22 23 26
rect 19 18 23 22
rect 19 17 52 18
rect 19 15 48 17
rect 50 15 52 17
rect 19 14 52 15
<< labels >>
rlabel alu0 13 36 13 36 6 zn
rlabel alu0 35 16 35 16 6 zn
rlabel alu0 37 57 37 57 6 zn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 32 44 32 6 d
rlabel alu1 44 24 44 24 6 a
rlabel alu1 44 40 44 40 6 c
rlabel alu1 36 48 36 48 6 b
rlabel alu1 44 48 44 48 6 b
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 60 20 60 20 6 d
rlabel alu1 52 32 52 32 6 d
rlabel alu1 52 40 52 40 6 c
rlabel alu1 60 48 60 48 6 c
<< end >>
