magic
tech scmos
timestamp 1199203536
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 31 70 33 74
rect 38 70 40 74
rect 48 70 50 74
rect 58 70 60 74
rect 68 70 70 74
rect 75 70 77 74
rect 85 70 87 74
rect 12 39 14 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 30 11 33
rect 19 30 21 42
rect 31 39 33 50
rect 38 47 40 50
rect 48 47 50 50
rect 58 47 60 50
rect 68 47 70 50
rect 38 45 43 47
rect 48 45 61 47
rect 41 41 43 45
rect 55 43 57 45
rect 59 43 61 45
rect 55 41 61 43
rect 65 45 70 47
rect 41 39 51 41
rect 31 37 37 39
rect 31 35 33 37
rect 35 35 37 37
rect 49 35 51 39
rect 65 35 67 45
rect 75 39 77 50
rect 85 39 87 42
rect 31 33 44 35
rect 49 33 67 35
rect 71 37 77 39
rect 71 35 73 37
rect 75 35 77 37
rect 71 33 77 35
rect 81 37 87 39
rect 81 35 83 37
rect 85 35 87 37
rect 81 33 87 35
rect 42 30 44 33
rect 52 30 54 33
rect 28 20 34 22
rect 28 18 30 20
rect 32 18 34 20
rect 28 16 34 18
rect 61 29 67 33
rect 61 27 63 29
rect 65 27 67 29
rect 84 28 86 33
rect 61 25 67 27
rect 9 11 11 16
rect 19 13 21 16
rect 28 13 30 16
rect 19 11 30 13
rect 42 13 44 18
rect 52 13 54 18
rect 84 10 86 15
<< ndif >>
rect 4 22 9 30
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 16 19 26
rect 21 28 28 30
rect 21 26 24 28
rect 26 26 28 28
rect 21 24 28 26
rect 21 16 26 24
rect 36 18 42 30
rect 44 28 52 30
rect 44 26 47 28
rect 49 26 52 28
rect 44 18 52 26
rect 54 22 59 30
rect 77 26 84 28
rect 77 24 79 26
rect 81 24 84 26
rect 77 22 84 24
rect 54 18 62 22
rect 36 14 40 18
rect 34 11 40 14
rect 34 9 36 11
rect 38 9 40 11
rect 34 7 40 9
rect 56 11 62 18
rect 79 15 84 22
rect 86 19 94 28
rect 86 17 89 19
rect 91 17 94 19
rect 86 15 94 17
rect 56 9 58 11
rect 60 9 62 11
rect 56 7 62 9
<< pdif >>
rect 7 62 12 70
rect 5 60 12 62
rect 5 58 7 60
rect 9 58 12 60
rect 5 53 12 58
rect 5 51 7 53
rect 9 51 12 53
rect 5 49 12 51
rect 7 42 12 49
rect 14 42 19 70
rect 21 68 31 70
rect 21 66 25 68
rect 27 66 31 68
rect 21 50 31 66
rect 33 50 38 70
rect 40 54 48 70
rect 40 52 43 54
rect 45 52 48 54
rect 40 50 48 52
rect 50 61 58 70
rect 50 59 53 61
rect 55 59 58 61
rect 50 50 58 59
rect 60 61 68 70
rect 60 59 63 61
rect 65 59 68 61
rect 60 54 68 59
rect 60 52 63 54
rect 65 52 68 54
rect 60 50 68 52
rect 70 50 75 70
rect 77 68 85 70
rect 77 66 80 68
rect 82 66 85 68
rect 77 61 85 66
rect 77 59 80 61
rect 82 59 85 61
rect 77 50 85 59
rect 21 42 26 50
rect 80 42 85 50
rect 87 63 92 70
rect 87 61 94 63
rect 87 59 90 61
rect 92 59 94 61
rect 87 54 94 59
rect 87 52 90 54
rect 92 52 94 54
rect 87 50 94 52
rect 87 42 92 50
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 2 54 10 55
rect 25 61 57 62
rect 25 59 53 61
rect 55 59 57 61
rect 25 58 57 59
rect 25 54 30 58
rect 2 53 30 54
rect 2 51 7 53
rect 9 51 30 53
rect 2 50 30 51
rect 2 29 6 50
rect 42 38 46 47
rect 73 46 79 54
rect 55 45 86 46
rect 55 43 57 45
rect 59 43 86 45
rect 55 42 86 43
rect 31 37 77 38
rect 31 35 33 37
rect 35 35 73 37
rect 75 35 77 37
rect 31 34 77 35
rect 82 37 86 42
rect 82 35 83 37
rect 85 35 86 37
rect 82 33 86 35
rect 57 29 71 30
rect 2 28 18 29
rect 2 26 14 28
rect 16 26 18 28
rect 2 25 18 26
rect 57 27 63 29
rect 65 27 71 29
rect 57 26 71 27
rect -2 11 98 12
rect -2 9 36 11
rect 38 9 58 11
rect 60 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 42 18 44 30
rect 52 18 54 30
rect 84 15 86 28
<< pmos >>
rect 12 42 14 70
rect 19 42 21 70
rect 31 50 33 70
rect 38 50 40 70
rect 48 50 50 70
rect 58 50 60 70
rect 68 50 70 70
rect 75 50 77 70
rect 85 42 87 70
<< polyct0 >>
rect 11 35 13 37
rect 30 18 32 20
<< polyct1 >>
rect 57 43 59 45
rect 33 35 35 37
rect 73 35 75 37
rect 83 35 85 37
rect 63 27 65 29
<< ndifct0 >>
rect 4 18 6 20
rect 24 26 26 28
rect 47 26 49 28
rect 79 24 81 26
rect 89 17 91 19
<< ndifct1 >>
rect 14 26 16 28
rect 36 9 38 11
rect 58 9 60 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 7 58 9 60
rect 25 66 27 68
rect 43 52 45 54
rect 63 59 65 61
rect 63 52 65 54
rect 80 66 82 68
rect 80 59 82 61
rect 90 59 92 61
rect 90 52 92 54
<< pdifct1 >>
rect 7 51 9 53
rect 53 59 55 61
<< alu0 >>
rect 23 66 25 68
rect 27 66 29 68
rect 23 65 29 66
rect 78 66 80 68
rect 82 66 84 68
rect 6 60 10 62
rect 6 58 7 60
rect 9 58 10 60
rect 6 55 10 58
rect 62 61 67 63
rect 62 59 63 61
rect 65 59 67 61
rect 30 50 31 58
rect 62 55 67 59
rect 78 61 84 66
rect 78 59 80 61
rect 82 59 84 61
rect 78 58 84 59
rect 89 61 94 63
rect 89 59 90 61
rect 92 59 94 61
rect 34 54 67 55
rect 89 54 94 59
rect 34 52 43 54
rect 45 52 63 54
rect 65 52 67 54
rect 34 51 67 52
rect 34 46 38 51
rect 22 42 38 46
rect 22 38 26 42
rect 89 52 90 54
rect 92 52 94 54
rect 89 50 94 52
rect 9 37 26 38
rect 9 35 11 37
rect 13 35 26 37
rect 9 34 26 35
rect 22 29 26 34
rect 90 29 94 50
rect 22 28 51 29
rect 22 26 24 28
rect 26 26 47 28
rect 49 26 51 28
rect 78 26 94 29
rect 22 25 51 26
rect 78 24 79 26
rect 81 25 94 26
rect 81 24 82 25
rect 78 21 82 24
rect 2 20 82 21
rect 2 18 4 20
rect 6 18 30 20
rect 32 18 82 20
rect 2 17 82 18
rect 88 19 92 21
rect 88 17 89 19
rect 91 17 92 19
rect 88 12 92 17
<< labels >>
rlabel alu0 17 36 17 36 6 an
rlabel alu0 36 27 36 27 6 an
rlabel alu0 50 53 50 53 6 an
rlabel alu0 64 57 64 57 6 an
rlabel alu0 80 23 80 23 6 bn
rlabel alu0 42 19 42 19 6 bn
rlabel alu0 92 44 92 44 6 bn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 36 36 36 36 6 a1
rlabel alu1 44 40 44 40 6 a1
rlabel alu1 28 56 28 56 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 52 36 52 36 6 a1
rlabel alu1 68 36 68 36 6 a1
rlabel alu1 60 36 60 36 6 a1
rlabel alu1 68 28 68 28 6 a2
rlabel alu1 60 28 60 28 6 a2
rlabel alu1 60 44 60 44 6 b
rlabel alu1 68 44 68 44 6 b
rlabel alu1 52 60 52 60 6 z
rlabel alu1 48 74 48 74 6 vdd
rlabel polyct1 84 36 84 36 6 b
rlabel alu1 76 48 76 48 6 b
<< end >>
