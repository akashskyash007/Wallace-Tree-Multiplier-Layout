magic
tech scmos
timestamp 1199203217
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 22 70 24 74
rect 29 70 31 74
rect 9 39 11 42
rect 22 39 24 42
rect 29 39 31 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 29 37 38 39
rect 29 35 34 37
rect 36 35 38 37
rect 29 33 38 35
rect 9 30 11 33
rect 19 25 21 33
rect 29 27 31 33
rect 9 11 11 16
rect 19 12 21 17
rect 29 15 31 19
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 16 9 19
rect 11 25 16 30
rect 24 25 29 27
rect 11 21 19 25
rect 11 19 14 21
rect 16 19 19 21
rect 11 17 19 19
rect 21 23 29 25
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 31 23 38 27
rect 31 21 34 23
rect 36 21 38 23
rect 31 19 38 21
rect 21 17 26 19
rect 11 16 16 17
<< pdif >>
rect 13 71 20 73
rect 13 70 15 71
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 55 9 60
rect 2 53 4 55
rect 6 53 9 55
rect 2 51 9 53
rect 4 42 9 51
rect 11 69 15 70
rect 17 70 20 71
rect 17 69 22 70
rect 11 42 22 69
rect 24 42 29 70
rect 31 64 36 70
rect 31 62 38 64
rect 31 60 34 62
rect 36 60 38 62
rect 31 58 38 60
rect 31 42 36 58
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 71 42 79
rect -2 69 15 71
rect 17 69 42 71
rect -2 68 42 69
rect 2 62 14 63
rect 2 60 4 62
rect 6 60 14 62
rect 2 57 14 60
rect 2 55 6 57
rect 2 53 4 55
rect 2 30 6 53
rect 26 49 38 55
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 18 39 22 47
rect 18 37 30 39
rect 18 35 21 37
rect 23 35 30 37
rect 18 33 30 35
rect 34 37 38 49
rect 36 35 38 37
rect 34 33 38 35
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 16 11 30
rect 19 17 21 25
rect 29 19 31 27
<< pmos >>
rect 9 42 11 70
rect 22 42 24 70
rect 29 42 31 70
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 21 35 23 37
rect 34 35 36 37
<< ndifct0 >>
rect 14 19 16 21
rect 24 21 26 23
rect 34 21 36 23
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 34 60 36 62
<< pdifct1 >>
rect 4 60 6 62
rect 4 53 6 55
rect 15 69 17 71
<< alu0 >>
rect 18 62 38 63
rect 18 60 34 62
rect 36 60 38 62
rect 18 59 38 60
rect 6 51 7 57
rect 18 54 22 59
rect 10 50 22 54
rect 10 37 14 50
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 33 33 34 49
rect 10 25 27 29
rect 23 23 27 25
rect 12 21 18 22
rect 12 19 14 21
rect 16 19 18 21
rect 23 21 24 23
rect 26 21 27 23
rect 23 19 27 21
rect 32 23 38 24
rect 32 21 34 23
rect 36 21 38 23
rect 12 12 18 19
rect 32 12 38 21
<< labels >>
rlabel alu0 12 39 12 39 6 zn
rlabel alu0 25 24 25 24 6 zn
rlabel alu0 28 61 28 61 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 36 28 36 6 a
rlabel alu1 20 40 20 40 6 a
rlabel alu1 28 52 28 52 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 44 36 44 6 b
<< end >>
