magic
tech scmos
timestamp 1199470007
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -2 48 52 104
<< pwell >>
rect -2 -4 52 48
<< poly >>
rect 15 78 17 82
rect 23 78 25 82
rect 37 73 39 78
rect 15 43 17 56
rect 23 52 25 56
rect 37 52 39 56
rect 23 49 27 52
rect 13 41 21 43
rect 13 39 17 41
rect 19 39 21 41
rect 13 37 21 39
rect 25 42 27 49
rect 32 50 39 52
rect 32 48 34 50
rect 36 48 39 50
rect 32 46 39 48
rect 25 40 32 42
rect 25 38 28 40
rect 30 38 32 40
rect 13 23 15 37
rect 25 36 32 38
rect 25 23 27 36
rect 37 26 39 46
rect 13 12 15 17
rect 25 12 27 17
rect 37 12 39 17
<< ndif >>
rect 30 23 37 26
rect 4 17 13 23
rect 15 21 25 23
rect 15 19 19 21
rect 21 19 25 21
rect 15 17 25 19
rect 27 21 37 23
rect 27 19 31 21
rect 33 19 37 21
rect 27 17 37 19
rect 39 24 47 26
rect 39 22 43 24
rect 45 22 47 24
rect 39 20 47 22
rect 39 17 44 20
rect 4 11 11 17
rect 4 9 7 11
rect 9 9 11 11
rect 4 7 11 9
<< pdif >>
rect 10 70 15 78
rect 7 68 15 70
rect 7 66 9 68
rect 11 66 15 68
rect 7 60 15 66
rect 7 58 9 60
rect 11 58 15 60
rect 7 56 15 58
rect 17 56 23 78
rect 25 73 35 78
rect 25 71 37 73
rect 25 69 29 71
rect 31 69 37 71
rect 25 56 37 69
rect 39 70 44 73
rect 39 68 47 70
rect 39 66 43 68
rect 45 66 47 68
rect 39 60 47 66
rect 39 58 43 60
rect 45 58 47 60
rect 39 56 47 58
<< alu1 >>
rect -2 95 52 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 52 95
rect -2 88 52 93
rect 8 68 12 73
rect 8 66 9 68
rect 11 66 12 68
rect 8 60 12 66
rect 8 58 9 60
rect 11 58 12 60
rect 8 23 12 58
rect 18 63 22 73
rect 28 71 32 88
rect 28 69 29 71
rect 31 69 32 71
rect 28 67 32 69
rect 42 68 46 70
rect 42 66 43 68
rect 45 66 46 68
rect 18 57 32 63
rect 18 44 22 53
rect 28 51 32 57
rect 42 60 46 66
rect 42 58 43 60
rect 45 58 46 60
rect 28 50 38 51
rect 28 48 34 50
rect 36 48 38 50
rect 28 47 38 48
rect 16 41 22 44
rect 42 41 46 58
rect 16 39 17 41
rect 19 39 22 41
rect 16 38 22 39
rect 18 32 22 38
rect 26 40 46 41
rect 26 38 28 40
rect 30 38 46 40
rect 26 37 46 38
rect 18 27 33 32
rect 42 24 46 37
rect 8 21 22 23
rect 8 19 19 21
rect 21 19 22 21
rect 8 17 22 19
rect 30 21 34 23
rect 30 19 31 21
rect 33 19 34 21
rect 42 22 43 24
rect 45 22 46 24
rect 42 20 46 22
rect 30 12 34 19
rect -2 11 52 12
rect -2 9 7 11
rect 9 9 52 11
rect -2 7 52 9
rect -2 5 19 7
rect 21 5 29 7
rect 31 5 52 7
rect -2 0 52 5
<< ptie >>
rect 17 7 33 9
rect 17 5 19 7
rect 21 5 29 7
rect 31 5 33 7
rect 17 3 33 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 13 17 15 23
rect 25 17 27 23
rect 37 17 39 26
<< pmos >>
rect 15 56 17 78
rect 23 56 25 78
rect 37 56 39 73
<< polyct1 >>
rect 17 39 19 41
rect 34 48 36 50
rect 28 38 30 40
<< ndifct1 >>
rect 19 19 21 21
rect 31 19 33 21
rect 43 22 45 24
rect 7 9 9 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 19 5 21 7
rect 29 5 31 7
<< pdifct1 >>
rect 9 66 11 68
rect 9 58 11 60
rect 29 69 31 71
rect 43 66 45 68
rect 43 58 45 60
<< labels >>
rlabel ndifct1 20 20 20 20 6 z
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 65 20 65 6 a
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 30 30 30 6 b
rlabel alu1 30 55 30 55 6 a
rlabel alu1 25 94 25 94 6 vdd
rlabel alu1 36 39 36 39 6 an
rlabel alu1 44 45 44 45 6 an
<< end >>
