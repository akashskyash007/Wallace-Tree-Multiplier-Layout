magic
tech scmos
timestamp 1199202651
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 65 41 70
rect 9 45 11 48
rect 9 43 15 45
rect 9 41 11 43
rect 13 41 15 43
rect 9 39 15 41
rect 19 39 21 48
rect 29 39 31 48
rect 10 30 12 39
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 39 39 41 48
rect 39 37 48 39
rect 39 35 43 37
rect 45 35 48 37
rect 17 33 31 35
rect 17 30 19 33
rect 29 30 31 33
rect 36 33 48 35
rect 36 30 38 33
rect 46 30 48 33
rect 53 37 59 39
rect 53 35 55 37
rect 57 35 59 37
rect 53 33 59 35
rect 53 30 55 33
rect 10 8 12 13
rect 17 8 19 13
rect 29 6 31 10
rect 36 6 38 10
rect 46 6 48 10
rect 53 6 55 10
<< ndif >>
rect 3 28 10 30
rect 3 26 5 28
rect 7 26 10 28
rect 3 21 10 26
rect 3 19 5 21
rect 7 19 10 21
rect 3 17 10 19
rect 5 13 10 17
rect 12 13 17 30
rect 19 14 29 30
rect 19 13 23 14
rect 21 12 23 13
rect 25 12 29 14
rect 21 10 29 12
rect 31 10 36 30
rect 38 21 46 30
rect 38 19 41 21
rect 43 19 46 21
rect 38 10 46 19
rect 48 10 53 30
rect 55 21 62 30
rect 55 19 58 21
rect 60 19 62 21
rect 55 14 62 19
rect 55 12 58 14
rect 60 12 62 14
rect 55 10 62 12
<< pdif >>
rect 2 63 9 65
rect 2 61 4 63
rect 6 61 9 63
rect 2 48 9 61
rect 11 61 19 65
rect 11 59 14 61
rect 16 59 19 61
rect 11 53 19 59
rect 11 51 14 53
rect 16 51 19 53
rect 11 48 19 51
rect 21 63 29 65
rect 21 61 24 63
rect 26 61 29 63
rect 21 48 29 61
rect 31 61 39 65
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 48 39 51
rect 41 63 49 65
rect 41 61 44 63
rect 46 61 49 63
rect 41 55 49 61
rect 41 53 44 55
rect 46 53 49 55
rect 41 48 49 53
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 2 53 38 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 51 38 53
rect 2 50 38 51
rect 2 28 6 50
rect 10 43 21 45
rect 10 41 11 43
rect 13 41 21 43
rect 10 39 21 41
rect 17 30 21 39
rect 25 42 55 46
rect 25 37 31 42
rect 51 38 55 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 30 47 35
rect 51 37 59 38
rect 51 35 55 37
rect 57 35 59 37
rect 51 34 59 35
rect 2 26 5 28
rect 17 26 47 30
rect 2 22 6 26
rect 2 21 47 22
rect 2 19 5 21
rect 7 19 41 21
rect 43 19 47 21
rect 2 18 47 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 10 13 12 30
rect 17 13 19 30
rect 29 10 31 30
rect 36 10 38 30
rect 46 10 48 30
rect 53 10 55 30
<< pmos >>
rect 9 48 11 65
rect 19 48 21 65
rect 29 48 31 65
rect 39 48 41 65
<< polyct1 >>
rect 11 41 13 43
rect 27 35 29 37
rect 43 35 45 37
rect 55 35 57 37
<< ndifct0 >>
rect 6 26 7 28
rect 23 12 25 14
rect 58 19 60 21
rect 58 12 60 14
<< ndifct1 >>
rect 5 26 6 28
rect 5 19 7 21
rect 41 19 43 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 61 6 63
rect 14 59 16 61
rect 24 61 26 63
rect 44 61 46 63
rect 44 53 46 55
<< pdifct1 >>
rect 14 51 16 53
rect 34 59 36 61
rect 34 51 36 53
<< alu0 >>
rect 3 63 7 68
rect 23 63 27 68
rect 43 63 47 68
rect 3 61 4 63
rect 6 61 7 63
rect 3 59 7 61
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 23 61 24 63
rect 26 61 27 63
rect 23 59 27 61
rect 13 54 17 59
rect 43 61 44 63
rect 46 61 47 63
rect 43 55 47 61
rect 43 53 44 55
rect 46 53 47 55
rect 43 51 47 53
rect 6 28 8 30
rect 7 26 8 28
rect 6 22 8 26
rect 56 21 62 22
rect 56 19 58 21
rect 60 19 62 21
rect 21 14 27 15
rect 21 12 23 14
rect 25 12 27 14
rect 56 14 62 19
rect 56 12 58 14
rect 60 12 62 14
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 b
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 40 28 40 6 a
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 b
rlabel alu1 44 32 44 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 36 60 36 60 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 44 52 44 6 a
<< end >>
