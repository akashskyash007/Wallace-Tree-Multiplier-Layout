magic
tech scmos
timestamp 1199543205
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 11 41 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 67 75 69 79
rect 23 51 43 53
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 17 41 23 43
rect 47 41 49 55
rect 67 43 69 55
rect 11 39 19 41
rect 21 39 49 41
rect 11 25 13 39
rect 17 37 23 39
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 23 27 43 29
rect 23 24 25 27
rect 35 24 37 27
rect 47 25 49 39
rect 57 41 69 43
rect 57 39 59 41
rect 61 39 69 41
rect 57 37 69 39
rect 67 25 69 37
rect 67 11 69 15
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 11 11 19
rect 3 9 5 11
rect 7 9 11 11
rect 3 6 11 9
rect 13 24 18 25
rect 42 24 47 25
rect 13 6 23 24
rect 25 21 35 24
rect 25 19 29 21
rect 31 19 35 21
rect 25 6 35 19
rect 37 6 47 24
rect 49 15 67 25
rect 69 21 77 25
rect 69 19 73 21
rect 75 19 77 21
rect 69 15 77 19
rect 49 11 65 15
rect 49 9 53 11
rect 55 9 61 11
rect 63 9 65 11
rect 49 6 65 9
<< pdif >>
rect 3 91 11 94
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 56 23 94
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 56 35 59
rect 37 56 47 94
rect 13 55 18 56
rect 42 55 47 56
rect 49 91 65 94
rect 49 89 53 91
rect 55 89 61 91
rect 63 89 65 91
rect 49 75 65 89
rect 49 55 67 75
rect 69 71 77 75
rect 69 69 73 71
rect 75 69 77 71
rect 69 61 77 69
rect 69 59 73 61
rect 75 59 77 61
rect 69 55 77 59
<< alu1 >>
rect -2 95 82 100
rect -2 93 73 95
rect 75 93 82 95
rect -2 91 82 93
rect -2 89 5 91
rect 7 89 53 91
rect 55 89 61 91
rect 63 89 82 91
rect -2 88 82 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 4 59 5 61
rect 7 59 8 61
rect 4 57 8 59
rect 18 41 22 83
rect 18 39 19 41
rect 21 39 22 41
rect 4 21 8 23
rect 4 19 5 21
rect 7 19 8 21
rect 4 12 8 19
rect 18 17 22 39
rect 28 81 32 83
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 28 21 32 59
rect 38 78 76 82
rect 38 51 42 78
rect 38 49 39 51
rect 41 49 42 51
rect 38 47 42 49
rect 58 41 62 73
rect 58 39 59 41
rect 61 39 62 41
rect 58 32 62 39
rect 37 31 62 32
rect 37 29 39 31
rect 41 29 62 31
rect 37 28 62 29
rect 28 19 29 21
rect 31 19 32 21
rect 28 17 32 19
rect 58 17 62 28
rect 72 71 76 78
rect 72 69 73 71
rect 75 69 76 71
rect 72 61 76 69
rect 72 59 73 61
rect 75 59 76 61
rect 72 21 76 59
rect 72 19 73 21
rect 75 19 76 21
rect 72 17 76 19
rect -2 11 82 12
rect -2 9 5 11
rect 7 9 53 11
rect 55 9 61 11
rect 63 9 82 11
rect -2 0 82 9
<< ntie >>
rect 71 95 77 97
rect 71 93 73 95
rect 75 93 77 95
rect 71 86 77 93
<< nmos >>
rect 11 6 13 25
rect 23 6 25 24
rect 35 6 37 24
rect 47 6 49 25
rect 67 15 69 25
<< pmos >>
rect 11 55 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 47 55 49 94
rect 67 55 69 75
<< polyct1 >>
rect 39 49 41 51
rect 19 39 21 41
rect 39 29 41 31
rect 59 39 61 41
<< ndifct1 >>
rect 5 19 7 21
rect 5 9 7 11
rect 29 19 31 21
rect 73 19 75 21
rect 53 9 55 11
rect 61 9 63 11
<< ntiect1 >>
rect 73 93 75 95
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 5 69 7 71
rect 5 59 7 61
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
rect 53 89 55 91
rect 61 89 63 91
rect 73 69 75 71
rect 73 59 75 61
<< labels >>
rlabel alu1 30 50 30 50 6 nq
rlabel alu1 20 50 20 50 6 i
rlabel alu1 40 6 40 6 6 vss
rlabel polyct1 40 30 40 30 6 cmd
rlabel alu1 50 30 50 30 6 cmd
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 60 45 60 45 6 cmd
<< end >>
