magic
tech scmos
timestamp 1199203043
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 13 64 15 69
rect 20 64 22 69
rect 27 64 29 69
rect 34 64 36 69
rect 44 57 46 61
rect 51 57 53 61
rect 58 57 60 61
rect 65 57 67 61
rect 13 36 15 39
rect 2 34 15 36
rect 2 32 4 34
rect 6 32 11 34
rect 2 30 11 32
rect 9 18 11 30
rect 20 29 22 39
rect 27 36 29 39
rect 34 36 36 39
rect 44 36 46 39
rect 27 33 30 36
rect 34 34 46 36
rect 17 27 23 29
rect 17 25 19 27
rect 21 25 23 27
rect 17 23 23 25
rect 28 27 30 33
rect 28 25 34 27
rect 28 23 30 25
rect 32 23 34 25
rect 19 18 21 23
rect 28 21 34 23
rect 31 18 33 21
rect 41 18 43 34
rect 51 27 53 39
rect 58 30 60 39
rect 65 36 67 39
rect 65 34 73 36
rect 67 32 69 34
rect 71 32 73 34
rect 67 30 73 32
rect 47 25 53 27
rect 47 23 49 25
rect 51 23 53 25
rect 57 28 63 30
rect 57 26 59 28
rect 61 26 63 28
rect 57 24 63 26
rect 47 21 53 23
rect 57 17 63 19
rect 57 15 59 17
rect 61 15 63 17
rect 57 13 63 15
rect 9 7 11 12
rect 19 7 21 12
rect 31 7 33 12
rect 41 9 43 12
rect 57 9 59 13
rect 41 7 59 9
<< ndif >>
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 16 19 18
rect 11 14 14 16
rect 16 14 19 16
rect 11 12 19 14
rect 21 12 31 18
rect 33 16 41 18
rect 33 14 36 16
rect 38 14 41 16
rect 33 12 41 14
rect 43 16 50 18
rect 43 14 46 16
rect 48 14 50 16
rect 43 12 50 14
rect 23 7 29 12
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< pdif >>
rect 4 67 11 69
rect 4 65 7 67
rect 9 65 11 67
rect 4 64 11 65
rect 4 39 13 64
rect 15 39 20 64
rect 22 39 27 64
rect 29 39 34 64
rect 36 57 41 64
rect 36 49 44 57
rect 36 47 39 49
rect 41 47 44 49
rect 36 39 44 47
rect 46 39 51 57
rect 53 39 58 57
rect 60 39 65 57
rect 67 55 74 57
rect 67 53 70 55
rect 72 53 74 55
rect 67 48 74 53
rect 67 46 70 48
rect 72 46 74 48
rect 67 39 74 46
<< alu1 >>
rect -2 67 82 72
rect -2 65 7 67
rect 9 65 47 67
rect 49 65 69 67
rect 71 65 82 67
rect -2 64 82 65
rect 2 54 62 58
rect 2 34 6 54
rect 10 49 43 50
rect 10 47 39 49
rect 41 47 43 49
rect 10 46 43 47
rect 2 32 4 34
rect 2 30 6 32
rect 10 18 14 46
rect 58 42 62 54
rect 18 38 53 42
rect 58 38 73 42
rect 18 27 22 38
rect 49 34 53 38
rect 67 34 73 38
rect 18 25 19 27
rect 21 25 22 27
rect 33 26 39 34
rect 49 30 62 34
rect 67 32 69 34
rect 71 32 73 34
rect 67 31 73 32
rect 58 28 62 30
rect 58 26 59 28
rect 61 26 62 28
rect 18 23 22 25
rect 28 25 53 26
rect 28 23 30 25
rect 32 23 49 25
rect 51 23 53 25
rect 58 24 62 26
rect 28 22 53 23
rect 66 19 70 27
rect 10 16 40 18
rect 10 14 14 16
rect 16 14 36 16
rect 38 14 40 16
rect 10 13 40 14
rect 58 17 70 19
rect 58 15 59 17
rect 61 15 70 17
rect 58 13 70 15
rect -2 7 82 8
rect -2 5 25 7
rect 27 5 69 7
rect 71 5 82 7
rect -2 0 82 5
<< ptie >>
rect 67 7 73 24
rect 67 5 69 7
rect 71 5 73 7
rect 67 3 73 5
<< ntie >>
rect 45 67 73 69
rect 45 65 47 67
rect 49 65 69 67
rect 71 65 73 67
rect 45 63 73 65
<< nmos >>
rect 9 12 11 18
rect 19 12 21 18
rect 31 12 33 18
rect 41 12 43 18
<< pmos >>
rect 13 39 15 64
rect 20 39 22 64
rect 27 39 29 64
rect 34 39 36 64
rect 44 39 46 57
rect 51 39 53 57
rect 58 39 60 57
rect 65 39 67 57
<< polyct1 >>
rect 4 32 6 34
rect 19 25 21 27
rect 30 23 32 25
rect 69 32 71 34
rect 49 23 51 25
rect 59 26 61 28
rect 59 15 61 17
<< ndifct0 >>
rect 4 14 6 16
rect 46 14 48 16
<< ndifct1 >>
rect 14 14 16 16
rect 36 14 38 16
rect 25 5 27 7
<< ntiect1 >>
rect 47 65 49 67
rect 69 65 71 67
<< ptiect1 >>
rect 69 5 71 7
<< pdifct0 >>
rect 70 53 72 55
rect 70 46 72 48
<< pdifct1 >>
rect 7 65 9 67
rect 39 47 41 49
<< alu0 >>
rect 6 30 7 36
rect 68 55 74 64
rect 68 53 70 55
rect 72 53 74 55
rect 68 48 74 53
rect 68 46 70 48
rect 72 46 74 48
rect 68 45 74 46
rect 3 16 7 18
rect 3 14 4 16
rect 6 14 7 16
rect 3 8 7 14
rect 45 16 49 18
rect 45 14 46 16
rect 48 14 49 16
rect 45 8 49 14
<< labels >>
rlabel alu1 4 44 4 44 6 a
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 32 20 32 6 b
rlabel alu1 12 28 12 28 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 56 28 56 6 a
rlabel alu1 20 56 20 56 6 a
rlabel alu1 12 56 12 56 6 a
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 36 16 36 16 6 z
rlabel alu1 44 24 44 24 6 c
rlabel alu1 36 28 36 28 6 c
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 56 44 56 6 a
rlabel alu1 36 56 36 56 6 a
rlabel alu1 40 68 40 68 6 vdd
rlabel polyct1 60 16 60 16 6 d
rlabel alu1 52 32 52 32 6 b
rlabel alu1 60 48 60 48 6 a
rlabel alu1 52 56 52 56 6 a
rlabel alu1 68 20 68 20 6 d
rlabel alu1 68 40 68 40 6 a
<< end >>
