magic
tech scmos
timestamp 1199202253
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 10 69 12 73
rect 20 61 22 65
rect 10 40 12 45
rect 20 40 22 45
rect 10 38 30 40
rect 10 30 12 38
rect 20 36 26 38
rect 28 36 30 38
rect 20 34 30 36
rect 20 30 22 34
rect 10 15 12 20
rect 20 15 22 20
<< ndif >>
rect 2 21 10 30
rect 2 19 4 21
rect 6 20 10 21
rect 12 28 20 30
rect 12 26 15 28
rect 17 26 20 28
rect 12 20 20 26
rect 22 24 30 30
rect 22 22 26 24
rect 28 22 30 24
rect 22 20 30 22
rect 6 19 8 20
rect 2 17 8 19
<< pdif >>
rect 2 67 10 69
rect 2 65 5 67
rect 7 65 10 67
rect 2 60 10 65
rect 2 58 5 60
rect 7 58 10 60
rect 2 45 10 58
rect 12 61 17 69
rect 12 53 20 61
rect 12 51 15 53
rect 17 51 20 53
rect 12 45 20 51
rect 22 59 30 61
rect 22 57 25 59
rect 27 57 30 59
rect 22 52 30 57
rect 22 50 25 52
rect 27 50 30 52
rect 22 45 30 50
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 53 19 54
rect 2 51 15 53
rect 17 51 19 53
rect 2 50 19 51
rect 2 31 6 50
rect 17 42 30 46
rect 26 38 30 42
rect 28 36 30 38
rect 26 33 30 36
rect 2 28 22 31
rect 2 26 15 28
rect 17 26 22 28
rect 2 25 22 26
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 10 20 12 30
rect 20 20 22 30
<< pmos >>
rect 10 45 12 69
rect 20 45 22 61
<< polyct1 >>
rect 26 36 28 38
<< ndifct0 >>
rect 4 19 6 21
rect 26 22 28 24
<< ndifct1 >>
rect 15 26 17 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 5 65 7 67
rect 5 58 7 60
rect 25 57 27 59
rect 25 50 27 52
<< pdifct1 >>
rect 15 51 17 53
<< alu0 >>
rect 3 67 9 68
rect 3 65 5 67
rect 7 65 9 67
rect 3 60 9 65
rect 3 58 5 60
rect 7 58 9 60
rect 3 57 9 58
rect 23 59 29 68
rect 23 57 25 59
rect 27 57 29 59
rect 23 52 29 57
rect 23 50 25 52
rect 27 50 29 52
rect 23 49 29 50
rect 24 35 26 42
rect 25 24 29 26
rect 25 22 26 24
rect 28 22 29 24
rect 2 21 8 22
rect 2 19 4 21
rect 6 19 8 21
rect 2 12 8 19
rect 25 12 29 22
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 28 20 28 6 z
rlabel alu1 20 44 20 44 6 a
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 36 28 36 6 a
<< end >>
