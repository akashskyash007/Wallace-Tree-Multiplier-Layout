magic
tech scmos
timestamp 1199542711
<< ab >>
rect 0 0 40 100
<< nwell >>
rect -5 48 45 105
<< pwell >>
rect -5 -5 45 48
<< poly >>
rect 19 94 21 98
rect 27 94 29 98
rect 19 53 21 56
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 13 47 23 49
rect 13 25 15 47
rect 27 43 29 56
rect 27 41 33 43
rect 25 39 29 41
rect 31 39 33 41
rect 25 37 33 39
rect 25 25 27 37
rect 13 11 15 15
rect 25 11 27 15
<< ndif >>
rect 5 15 13 25
rect 15 21 25 25
rect 15 19 19 21
rect 21 19 25 21
rect 15 15 25 19
rect 27 15 35 25
rect 5 11 11 15
rect 29 11 35 15
rect 5 9 7 11
rect 9 9 11 11
rect 5 7 11 9
rect 29 9 31 11
rect 33 9 35 11
rect 29 7 35 9
<< pdif >>
rect 14 85 19 94
rect 7 81 19 85
rect 7 79 9 81
rect 11 79 19 81
rect 7 71 19 79
rect 7 69 9 71
rect 11 69 19 71
rect 7 61 19 69
rect 7 59 9 61
rect 11 59 19 61
rect 7 56 19 59
rect 21 56 27 94
rect 29 91 37 94
rect 29 89 33 91
rect 35 89 37 91
rect 29 56 37 89
rect 7 55 13 56
<< alu1 >>
rect -2 91 42 100
rect -2 89 33 91
rect 35 89 42 91
rect -2 88 42 89
rect 8 81 12 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 71 12 79
rect 8 69 9 71
rect 11 69 12 71
rect 8 61 12 69
rect 8 59 9 61
rect 11 59 12 61
rect 8 22 12 59
rect 18 51 22 83
rect 18 49 19 51
rect 21 49 22 51
rect 18 27 22 49
rect 28 41 32 83
rect 28 39 29 41
rect 31 39 32 41
rect 8 21 23 22
rect 8 19 19 21
rect 21 19 23 21
rect 8 18 23 19
rect 8 17 12 18
rect 28 17 32 39
rect -2 11 42 12
rect -2 9 7 11
rect 9 9 31 11
rect 33 9 42 11
rect -2 0 42 9
<< nmos >>
rect 13 15 15 25
rect 25 15 27 25
<< pmos >>
rect 19 56 21 94
rect 27 56 29 94
<< polyct1 >>
rect 19 49 21 51
rect 29 39 31 41
<< ndifct1 >>
rect 19 19 21 21
rect 7 9 9 11
rect 31 9 33 11
<< pdifct1 >>
rect 9 79 11 81
rect 9 69 11 71
rect 9 59 11 61
rect 33 89 35 91
<< labels >>
rlabel alu1 20 6 20 6 6 vss
rlabel ndifct1 20 20 20 20 6 nq
rlabel alu1 10 50 10 50 6 nq
rlabel alu1 20 55 20 55 6 i1
rlabel alu1 20 94 20 94 6 vdd
rlabel alu1 30 50 30 50 6 i0
<< end >>
