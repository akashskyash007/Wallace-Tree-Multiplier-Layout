magic
tech scmos
timestamp 1199202721
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 15 62 17 67
rect 25 62 27 67
rect 35 62 37 67
rect 45 62 47 67
rect 15 39 17 42
rect 25 39 27 42
rect 9 37 27 39
rect 9 35 11 37
rect 13 35 27 37
rect 9 33 27 35
rect 15 30 17 33
rect 25 30 27 33
rect 35 39 37 42
rect 45 39 47 42
rect 35 37 47 39
rect 35 35 43 37
rect 45 35 47 37
rect 35 33 47 35
rect 35 30 37 33
rect 45 30 47 33
rect 15 12 17 17
rect 25 12 27 17
rect 35 12 37 17
rect 45 13 47 17
<< ndif >>
rect 10 23 15 30
rect 8 21 15 23
rect 8 19 10 21
rect 12 19 15 21
rect 8 17 15 19
rect 17 28 25 30
rect 17 26 20 28
rect 22 26 25 28
rect 17 17 25 26
rect 27 28 35 30
rect 27 26 30 28
rect 32 26 35 28
rect 27 21 35 26
rect 27 19 30 21
rect 32 19 35 21
rect 27 17 35 19
rect 37 21 45 30
rect 37 19 40 21
rect 42 19 45 21
rect 37 17 45 19
rect 47 28 54 30
rect 47 26 50 28
rect 52 26 54 28
rect 47 24 54 26
rect 47 17 52 24
<< pdif >>
rect 6 60 15 62
rect 6 58 9 60
rect 11 58 15 60
rect 6 53 15 58
rect 6 51 9 53
rect 11 51 15 53
rect 6 42 15 51
rect 17 53 25 62
rect 17 51 20 53
rect 22 51 25 53
rect 17 46 25 51
rect 17 44 20 46
rect 22 44 25 46
rect 17 42 25 44
rect 27 60 35 62
rect 27 58 30 60
rect 32 58 35 60
rect 27 53 35 58
rect 27 51 30 53
rect 32 51 35 53
rect 27 42 35 51
rect 37 53 45 62
rect 37 51 40 53
rect 42 51 45 53
rect 37 46 45 51
rect 37 44 40 46
rect 42 44 45 46
rect 37 42 45 44
rect 47 60 54 62
rect 47 58 50 60
rect 52 58 54 60
rect 47 42 54 58
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 18 53 23 55
rect 18 51 20 53
rect 22 51 23 53
rect 18 46 23 51
rect 39 53 43 55
rect 39 51 40 53
rect 42 51 43 53
rect 39 46 43 51
rect 18 44 20 46
rect 22 44 40 46
rect 42 44 43 46
rect 18 42 43 44
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 2 25 6 33
rect 18 28 23 42
rect 50 38 54 47
rect 41 37 54 38
rect 41 35 43 37
rect 45 35 54 37
rect 41 33 54 35
rect 18 26 20 28
rect 22 26 23 28
rect 18 24 23 26
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 15 17 17 30
rect 25 17 27 30
rect 35 17 37 30
rect 45 17 47 30
<< pmos >>
rect 15 42 17 62
rect 25 42 27 62
rect 35 42 37 62
rect 45 42 47 62
<< polyct1 >>
rect 11 35 13 37
rect 43 35 45 37
<< ndifct0 >>
rect 10 19 12 21
rect 30 26 32 28
rect 30 19 32 21
rect 40 19 42 21
rect 50 26 52 28
<< ndifct1 >>
rect 20 26 22 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 9 58 11 60
rect 9 51 11 53
rect 30 58 32 60
rect 30 51 32 53
rect 50 58 52 60
<< pdifct1 >>
rect 20 51 22 53
rect 20 44 22 46
rect 40 51 42 53
rect 40 44 42 46
<< alu0 >>
rect 8 60 12 68
rect 8 58 9 60
rect 11 58 12 60
rect 8 53 12 58
rect 29 60 33 68
rect 29 58 30 60
rect 32 58 33 60
rect 8 51 9 53
rect 11 51 12 53
rect 8 49 12 51
rect 29 53 33 58
rect 49 60 53 68
rect 49 58 50 60
rect 52 58 53 60
rect 49 56 53 58
rect 29 51 30 53
rect 32 51 33 53
rect 29 49 33 51
rect 28 28 54 29
rect 28 26 30 28
rect 32 26 50 28
rect 52 26 54 28
rect 28 25 54 26
rect 8 21 14 22
rect 28 21 33 25
rect 8 19 10 21
rect 12 19 30 21
rect 32 19 33 21
rect 8 17 33 19
rect 38 21 44 22
rect 38 19 40 21
rect 42 19 44 21
rect 38 12 44 19
<< labels >>
rlabel alu0 30 23 30 23 6 n1
rlabel alu0 20 19 20 19 6 n1
rlabel alu0 41 27 41 27 6 n1
rlabel alu1 4 32 4 32 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 40 20 40 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 44 36 44 6 z
rlabel alu1 28 44 28 44 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 36 44 36 6 a
rlabel alu1 52 40 52 40 6 a
<< end >>
