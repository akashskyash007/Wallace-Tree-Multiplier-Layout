magic
tech scmos
timestamp 1199203623
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 6 72 30 74
rect 6 63 8 72
rect 18 64 20 68
rect 28 64 30 72
rect 38 72 60 74
rect 38 64 40 72
rect 48 64 50 68
rect 58 64 60 72
rect 2 61 8 63
rect 2 59 4 61
rect 6 59 8 61
rect 2 57 8 59
rect 18 39 20 42
rect 8 37 20 39
rect 28 37 30 42
rect 38 38 40 42
rect 48 38 50 42
rect 58 39 60 42
rect 8 35 10 37
rect 12 35 14 37
rect 28 35 34 37
rect 8 33 14 35
rect 12 30 14 33
rect 22 29 24 33
rect 32 29 34 35
rect 48 36 54 38
rect 48 34 50 36
rect 52 34 54 36
rect 42 32 54 34
rect 58 37 64 39
rect 58 35 60 37
rect 62 35 64 37
rect 58 33 64 35
rect 42 29 44 32
rect 61 29 63 33
rect 12 14 14 19
rect 22 10 24 18
rect 32 14 34 18
rect 42 14 44 18
rect 61 10 63 18
rect 22 8 63 10
<< ndif >>
rect 2 23 12 30
rect 2 21 4 23
rect 6 21 12 23
rect 2 19 12 21
rect 14 29 19 30
rect 14 26 22 29
rect 14 24 17 26
rect 19 24 22 26
rect 14 19 22 24
rect 17 18 22 19
rect 24 27 32 29
rect 24 25 27 27
rect 29 25 32 27
rect 24 18 32 25
rect 34 27 42 29
rect 34 25 37 27
rect 39 25 42 27
rect 34 18 42 25
rect 44 22 61 29
rect 44 20 56 22
rect 58 20 61 22
rect 44 18 61 20
rect 63 27 70 29
rect 63 25 66 27
rect 68 25 70 27
rect 63 23 70 25
rect 63 18 68 23
<< pdif >>
rect 11 62 18 64
rect 11 60 13 62
rect 15 60 18 62
rect 11 42 18 60
rect 20 46 28 64
rect 20 44 23 46
rect 25 44 28 46
rect 20 42 28 44
rect 30 46 38 64
rect 30 44 33 46
rect 35 44 38 46
rect 30 42 38 44
rect 40 46 48 64
rect 40 44 43 46
rect 45 44 48 46
rect 40 42 48 44
rect 50 62 58 64
rect 50 60 53 62
rect 55 60 58 62
rect 50 42 58 60
rect 60 56 65 64
rect 60 54 67 56
rect 60 52 63 54
rect 65 52 67 54
rect 60 50 67 52
rect 60 42 65 50
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 39 6 47
rect 30 46 38 47
rect 30 44 33 46
rect 35 44 38 46
rect 2 37 14 39
rect 2 35 10 37
rect 12 35 14 37
rect 2 33 14 35
rect 30 41 38 44
rect 30 38 34 41
rect 50 41 62 47
rect 58 39 62 41
rect 25 34 34 38
rect 25 27 31 34
rect 58 37 63 39
rect 58 35 60 37
rect 62 35 63 37
rect 58 33 63 35
rect 25 25 27 27
rect 29 25 31 27
rect 25 24 31 25
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 12 19 14 30
rect 22 18 24 29
rect 32 18 34 29
rect 42 18 44 29
rect 61 18 63 29
<< pmos >>
rect 18 42 20 64
rect 28 42 30 64
rect 38 42 40 64
rect 48 42 50 64
rect 58 42 60 64
<< polyct0 >>
rect 4 59 6 61
rect 50 34 52 36
<< polyct1 >>
rect 10 35 12 37
rect 60 35 62 37
<< ndifct0 >>
rect 4 21 6 23
rect 17 24 19 26
rect 37 25 39 27
rect 56 20 58 22
rect 66 25 68 27
<< ndifct1 >>
rect 27 25 29 27
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 13 60 15 62
rect 23 44 25 46
rect 43 44 45 46
rect 53 60 55 62
rect 63 52 65 54
<< pdifct1 >>
rect 33 44 35 46
<< alu0 >>
rect 3 61 7 63
rect 3 59 4 61
rect 6 59 7 61
rect 11 62 17 68
rect 11 60 13 62
rect 15 60 17 62
rect 11 59 17 60
rect 51 62 57 68
rect 51 60 53 62
rect 55 60 57 62
rect 51 59 57 60
rect 3 55 7 59
rect 3 54 70 55
rect 3 52 63 54
rect 65 52 70 54
rect 3 51 70 52
rect 17 46 27 47
rect 17 44 23 46
rect 25 44 27 46
rect 17 43 27 44
rect 17 28 21 43
rect 42 46 46 48
rect 42 44 43 46
rect 45 44 46 46
rect 42 38 46 44
rect 16 26 21 28
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 16 24 17 26
rect 19 24 21 26
rect 38 34 46 38
rect 49 36 53 38
rect 49 34 50 36
rect 52 34 53 36
rect 38 28 42 34
rect 49 31 53 34
rect 35 27 42 28
rect 35 25 37 27
rect 39 25 42 27
rect 35 24 42 25
rect 47 27 53 31
rect 66 29 70 51
rect 65 27 70 29
rect 16 22 21 24
rect 3 12 7 21
rect 17 21 21 22
rect 47 21 51 27
rect 65 25 66 27
rect 68 25 70 27
rect 17 17 51 21
rect 55 22 59 24
rect 65 23 70 25
rect 55 20 56 22
rect 58 20 59 22
rect 55 12 59 20
<< labels >>
rlabel alu0 5 57 5 57 6 bn
rlabel alu0 19 32 19 32 6 an
rlabel alu0 22 45 22 45 6 an
rlabel alu0 40 31 40 31 6 ai
rlabel alu0 51 32 51 32 6 an
rlabel alu0 44 41 44 41 6 ai
rlabel alu0 68 39 68 39 6 bn
rlabel alu0 36 53 36 53 6 bn
rlabel alu1 12 36 12 36 6 a
rlabel alu1 4 40 4 40 6 a
rlabel alu1 28 32 28 32 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 52 44 52 44 6 b
rlabel alu1 36 44 36 44 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 40 60 40 6 b
<< end >>
