magic
tech scmos
timestamp 1199542067
<< ab >>
rect 0 0 180 100
<< nwell >>
rect -5 48 185 105
<< pwell >>
rect -5 -5 185 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 155 94 157 98
rect 167 94 169 98
rect 35 83 37 87
rect 47 84 49 88
rect 83 78 85 82
rect 95 78 97 82
rect 71 72 73 76
rect 11 43 13 55
rect 23 43 25 55
rect 35 53 37 65
rect 47 63 49 66
rect 47 61 53 63
rect 47 59 49 61
rect 51 59 53 61
rect 47 57 53 59
rect 107 77 109 81
rect 119 77 121 81
rect 131 78 133 82
rect 29 51 37 53
rect 71 53 73 56
rect 83 53 85 56
rect 71 51 85 53
rect 95 53 97 56
rect 95 51 103 53
rect 29 49 31 51
rect 33 49 37 51
rect 29 47 37 49
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 97 49 99 51
rect 101 49 103 51
rect 97 47 103 49
rect 11 41 25 43
rect 37 41 43 43
rect 11 39 39 41
rect 41 39 43 41
rect 11 37 25 39
rect 37 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 63 41 69 43
rect 107 41 109 55
rect 119 43 121 55
rect 131 53 133 56
rect 127 51 133 53
rect 127 49 129 51
rect 131 49 133 51
rect 127 47 133 49
rect 155 43 157 55
rect 167 43 169 55
rect 63 39 65 41
rect 67 39 109 41
rect 63 37 69 39
rect 11 25 13 37
rect 23 25 25 37
rect 29 31 37 33
rect 29 29 31 31
rect 33 29 37 31
rect 47 29 49 37
rect 97 33 103 35
rect 77 31 83 33
rect 97 31 99 33
rect 101 31 103 33
rect 77 29 79 31
rect 81 29 83 31
rect 95 29 103 31
rect 29 27 37 29
rect 35 24 37 27
rect 71 27 85 29
rect 71 24 73 27
rect 83 24 85 27
rect 95 26 97 29
rect 107 27 109 39
rect 117 41 123 43
rect 137 41 143 43
rect 117 39 119 41
rect 121 39 139 41
rect 141 39 143 41
rect 117 37 123 39
rect 137 37 143 39
rect 147 41 169 43
rect 147 39 149 41
rect 151 39 169 41
rect 147 37 169 39
rect 127 31 133 33
rect 127 29 129 31
rect 131 29 133 31
rect 119 27 133 29
rect 35 11 37 15
rect 47 11 49 15
rect 71 12 73 16
rect 119 24 121 27
rect 131 24 133 27
rect 155 25 157 37
rect 167 25 169 37
rect 83 11 85 15
rect 95 11 97 15
rect 107 11 109 15
rect 119 11 121 15
rect 131 12 133 16
rect 11 2 13 6
rect 23 2 25 6
rect 155 2 157 6
rect 167 2 169 6
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 11 11 19
rect 3 9 5 11
rect 7 9 11 11
rect 3 6 11 9
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 6 23 19
rect 25 24 30 25
rect 39 24 47 29
rect 25 15 35 24
rect 37 15 47 24
rect 49 21 57 29
rect 102 26 107 27
rect 87 24 95 26
rect 49 19 53 21
rect 55 19 57 21
rect 49 15 57 19
rect 63 21 71 24
rect 63 19 65 21
rect 67 19 71 21
rect 63 17 71 19
rect 66 16 71 17
rect 73 16 83 24
rect 25 11 33 15
rect 75 15 83 16
rect 85 15 95 24
rect 97 23 107 26
rect 97 21 101 23
rect 103 21 107 23
rect 97 15 107 21
rect 109 24 117 27
rect 135 31 143 33
rect 135 29 139 31
rect 141 29 143 31
rect 135 27 143 29
rect 135 24 141 27
rect 109 15 119 24
rect 121 16 131 24
rect 133 16 141 24
rect 150 21 155 25
rect 121 15 129 16
rect 75 11 81 15
rect 123 11 129 15
rect 25 9 29 11
rect 31 9 33 11
rect 75 9 77 11
rect 79 9 81 11
rect 123 9 125 11
rect 127 9 129 11
rect 25 6 33 9
rect 75 7 81 9
rect 123 7 129 9
rect 147 11 155 21
rect 147 9 149 11
rect 151 9 155 11
rect 147 6 155 9
rect 157 21 167 25
rect 157 19 161 21
rect 163 19 167 21
rect 157 6 167 19
rect 169 21 177 25
rect 169 19 173 21
rect 175 19 177 21
rect 169 11 177 19
rect 169 9 173 11
rect 175 9 177 11
rect 169 6 177 9
<< pdif >>
rect 3 91 11 94
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 81 23 94
rect 13 79 17 81
rect 19 79 23 81
rect 13 71 23 79
rect 13 69 17 71
rect 19 69 23 71
rect 13 61 23 69
rect 13 59 17 61
rect 19 59 23 61
rect 13 55 23 59
rect 25 91 33 94
rect 25 89 29 91
rect 31 89 33 91
rect 25 83 33 89
rect 51 91 57 93
rect 51 89 53 91
rect 55 89 57 91
rect 51 84 57 89
rect 75 91 81 93
rect 123 91 129 93
rect 75 89 77 91
rect 79 89 81 91
rect 39 83 47 84
rect 25 65 35 83
rect 37 71 47 83
rect 37 69 41 71
rect 43 69 47 71
rect 37 66 47 69
rect 49 66 57 84
rect 75 78 81 89
rect 123 89 125 91
rect 127 89 129 91
rect 75 72 83 78
rect 37 65 42 66
rect 25 55 33 65
rect 63 61 71 72
rect 63 59 65 61
rect 67 59 71 61
rect 63 56 71 59
rect 73 56 83 72
rect 85 71 95 78
rect 85 69 89 71
rect 91 69 95 71
rect 85 56 95 69
rect 97 77 105 78
rect 123 78 129 89
rect 147 91 155 94
rect 147 89 149 91
rect 151 89 155 91
rect 147 81 155 89
rect 147 79 149 81
rect 151 79 155 81
rect 123 77 131 78
rect 97 61 107 77
rect 97 59 101 61
rect 103 59 107 61
rect 97 56 107 59
rect 102 55 107 56
rect 109 71 119 77
rect 109 69 113 71
rect 115 69 119 71
rect 109 61 119 69
rect 109 59 113 61
rect 115 59 119 61
rect 109 55 119 59
rect 121 56 131 77
rect 133 61 141 78
rect 147 71 155 79
rect 147 69 149 71
rect 151 69 155 71
rect 147 67 155 69
rect 133 59 143 61
rect 133 57 139 59
rect 141 57 143 59
rect 133 56 143 57
rect 121 55 126 56
rect 137 55 143 56
rect 150 55 155 67
rect 157 81 167 94
rect 157 79 161 81
rect 163 79 167 81
rect 157 71 167 79
rect 157 69 161 71
rect 163 69 167 71
rect 157 61 167 69
rect 157 59 161 61
rect 163 59 167 61
rect 157 55 167 59
rect 169 91 177 94
rect 169 89 173 91
rect 175 89 177 91
rect 169 81 177 89
rect 169 79 173 81
rect 175 79 177 81
rect 169 71 177 79
rect 169 69 173 71
rect 175 69 177 71
rect 169 61 177 69
rect 169 59 173 61
rect 175 59 177 61
rect 169 55 177 59
<< alu1 >>
rect -2 95 182 100
rect -2 93 65 95
rect 67 93 89 95
rect 91 93 101 95
rect 103 93 113 95
rect 115 93 137 95
rect 139 93 182 95
rect -2 91 182 93
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 53 91
rect 55 89 77 91
rect 79 89 125 91
rect 127 89 149 91
rect 151 89 173 91
rect 175 89 182 91
rect -2 88 182 89
rect 4 81 8 88
rect 18 82 22 83
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 15 81 22 82
rect 15 79 17 81
rect 19 79 22 81
rect 15 78 22 79
rect 18 72 22 78
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 15 71 22 72
rect 15 69 17 71
rect 19 69 22 71
rect 15 68 22 69
rect 18 62 22 68
rect 4 59 5 61
rect 7 59 8 61
rect 4 57 8 59
rect 15 61 22 62
rect 15 59 17 61
rect 19 59 22 61
rect 15 58 22 59
rect 4 21 8 23
rect 18 22 22 58
rect 4 19 5 21
rect 7 19 8 21
rect 4 12 8 19
rect 15 21 22 22
rect 15 19 17 21
rect 19 19 22 21
rect 15 18 22 19
rect 18 17 22 18
rect 28 82 32 83
rect 28 78 132 82
rect 28 52 32 78
rect 78 72 82 73
rect 112 72 116 73
rect 39 71 45 72
rect 39 69 41 71
rect 43 69 45 71
rect 39 68 45 69
rect 50 68 82 72
rect 87 71 116 72
rect 87 69 89 71
rect 91 69 113 71
rect 115 69 116 71
rect 87 68 116 69
rect 28 51 35 52
rect 28 49 31 51
rect 33 49 35 51
rect 28 48 35 49
rect 28 32 32 48
rect 39 42 43 68
rect 50 63 54 68
rect 37 41 43 42
rect 37 39 39 41
rect 41 39 43 41
rect 37 38 43 39
rect 28 31 35 32
rect 28 29 31 31
rect 33 29 35 31
rect 28 28 35 29
rect 28 17 32 28
rect 39 22 43 38
rect 48 61 54 63
rect 48 59 49 61
rect 51 59 54 61
rect 48 58 54 59
rect 64 61 68 63
rect 64 59 65 61
rect 67 59 68 61
rect 48 41 52 58
rect 48 39 49 41
rect 51 39 52 41
rect 48 37 52 39
rect 64 41 68 59
rect 64 39 65 41
rect 67 39 68 41
rect 39 21 57 22
rect 39 19 53 21
rect 55 19 57 21
rect 39 18 57 19
rect 64 21 68 39
rect 64 19 65 21
rect 67 19 68 21
rect 64 17 68 19
rect 78 51 82 68
rect 78 49 79 51
rect 81 49 82 51
rect 78 31 82 49
rect 78 29 79 31
rect 81 29 82 31
rect 78 17 82 29
rect 88 61 105 62
rect 88 59 101 61
rect 103 59 105 61
rect 88 58 105 59
rect 112 61 116 68
rect 112 59 113 61
rect 115 59 116 61
rect 88 22 92 58
rect 112 57 116 59
rect 128 52 132 78
rect 148 81 152 88
rect 148 79 149 81
rect 151 79 152 81
rect 148 71 152 79
rect 148 69 149 71
rect 151 69 152 71
rect 148 67 152 69
rect 158 82 162 83
rect 158 81 165 82
rect 158 79 161 81
rect 163 79 165 81
rect 158 78 165 79
rect 172 81 176 88
rect 172 79 173 81
rect 175 79 176 81
rect 158 72 162 78
rect 158 71 165 72
rect 158 69 161 71
rect 163 69 165 71
rect 158 68 165 69
rect 172 71 176 79
rect 172 69 173 71
rect 175 69 176 71
rect 158 62 162 68
rect 158 61 165 62
rect 97 51 132 52
rect 97 49 99 51
rect 101 49 129 51
rect 131 49 132 51
rect 97 48 132 49
rect 108 41 123 42
rect 108 39 119 41
rect 121 39 123 41
rect 108 38 123 39
rect 108 34 112 38
rect 97 33 112 34
rect 97 31 99 33
rect 101 31 112 33
rect 97 30 112 31
rect 128 31 132 48
rect 128 29 129 31
rect 131 29 132 31
rect 128 27 132 29
rect 138 59 142 61
rect 138 57 139 59
rect 141 57 142 59
rect 138 41 142 57
rect 158 59 161 61
rect 163 59 165 61
rect 158 58 165 59
rect 172 61 176 69
rect 172 59 173 61
rect 175 59 176 61
rect 138 39 139 41
rect 141 39 142 41
rect 138 31 142 39
rect 138 29 139 31
rect 141 29 142 31
rect 138 27 142 29
rect 148 41 152 43
rect 148 39 149 41
rect 151 39 152 41
rect 99 23 105 24
rect 99 22 101 23
rect 88 21 101 22
rect 103 22 105 23
rect 148 22 152 39
rect 103 21 152 22
rect 88 18 152 21
rect 158 22 162 58
rect 172 57 176 59
rect 158 21 165 22
rect 158 19 161 21
rect 163 19 165 21
rect 158 18 165 19
rect 172 21 176 23
rect 172 19 173 21
rect 175 19 176 21
rect 158 17 162 18
rect 172 12 176 19
rect -2 11 182 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 77 11
rect 79 9 125 11
rect 127 9 149 11
rect 151 9 173 11
rect 175 9 182 11
rect -2 7 182 9
rect -2 5 41 7
rect 43 5 53 7
rect 55 5 65 7
rect 67 5 89 7
rect 91 5 101 7
rect 103 5 113 7
rect 115 5 182 7
rect -2 0 182 5
<< ptie >>
rect 39 7 69 9
rect 87 7 117 9
rect 39 5 41 7
rect 43 5 53 7
rect 55 5 65 7
rect 67 5 69 7
rect 39 3 69 5
rect 87 5 89 7
rect 91 5 101 7
rect 103 5 113 7
rect 115 5 117 7
rect 87 3 117 5
<< ntie >>
rect 63 95 69 97
rect 63 93 65 95
rect 67 93 69 95
rect 87 95 117 97
rect 87 93 89 95
rect 91 93 101 95
rect 103 93 113 95
rect 115 93 117 95
rect 135 95 141 97
rect 135 93 137 95
rect 139 93 141 95
rect 63 86 69 93
rect 87 91 117 93
rect 135 86 141 93
<< nmos >>
rect 11 6 13 25
rect 23 6 25 25
rect 35 15 37 24
rect 47 15 49 29
rect 71 16 73 24
rect 83 15 85 24
rect 95 15 97 26
rect 107 15 109 27
rect 119 15 121 24
rect 131 16 133 24
rect 155 6 157 25
rect 167 6 169 25
<< pmos >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 65 37 83
rect 47 66 49 84
rect 71 56 73 72
rect 83 56 85 78
rect 95 56 97 78
rect 107 55 109 77
rect 119 55 121 77
rect 131 56 133 78
rect 155 55 157 94
rect 167 55 169 94
<< polyct1 >>
rect 49 59 51 61
rect 31 49 33 51
rect 79 49 81 51
rect 99 49 101 51
rect 39 39 41 41
rect 49 39 51 41
rect 129 49 131 51
rect 65 39 67 41
rect 31 29 33 31
rect 99 31 101 33
rect 79 29 81 31
rect 119 39 121 41
rect 139 39 141 41
rect 149 39 151 41
rect 129 29 131 31
<< ndifct1 >>
rect 5 19 7 21
rect 5 9 7 11
rect 17 19 19 21
rect 53 19 55 21
rect 65 19 67 21
rect 101 21 103 23
rect 139 29 141 31
rect 29 9 31 11
rect 77 9 79 11
rect 125 9 127 11
rect 149 9 151 11
rect 161 19 163 21
rect 173 19 175 21
rect 173 9 175 11
<< ntiect1 >>
rect 65 93 67 95
rect 89 93 91 95
rect 101 93 103 95
rect 113 93 115 95
rect 137 93 139 95
<< ptiect1 >>
rect 41 5 43 7
rect 53 5 55 7
rect 65 5 67 7
rect 89 5 91 7
rect 101 5 103 7
rect 113 5 115 7
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 5 69 7 71
rect 5 59 7 61
rect 17 79 19 81
rect 17 69 19 71
rect 17 59 19 61
rect 29 89 31 91
rect 53 89 55 91
rect 77 89 79 91
rect 41 69 43 71
rect 125 89 127 91
rect 65 59 67 61
rect 89 69 91 71
rect 149 89 151 91
rect 149 79 151 81
rect 101 59 103 61
rect 113 69 115 71
rect 113 59 115 61
rect 149 69 151 71
rect 139 57 141 59
rect 161 79 163 81
rect 161 69 163 71
rect 161 59 163 61
rect 173 89 175 91
rect 173 79 175 81
rect 173 69 175 71
rect 173 59 175 61
<< labels >>
rlabel alu1 30 50 30 50 6 a
rlabel alu1 20 50 20 50 6 cout
rlabel polyct1 50 40 50 40 6 b
rlabel alu1 50 50 50 50 6 b
rlabel polyct1 50 60 50 60 6 b
rlabel alu1 60 70 60 70 6 b
rlabel ptiect1 90 6 90 6 6 vss
rlabel alu1 80 45 80 45 6 b
rlabel alu1 70 70 70 70 6 b
rlabel ntiect1 90 94 90 94 6 vdd
rlabel alu1 160 50 160 50 6 sout
<< end >>
