magic
tech scmos
timestamp 1199203565
<< ab >>
rect 0 0 200 72
<< nwell >>
rect -5 32 205 77
<< pwell >>
rect -5 -5 205 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 99 66 101 70
rect 109 66 111 70
rect 119 66 121 70
rect 126 66 128 70
rect 136 66 138 70
rect 143 66 145 70
rect 153 66 155 70
rect 160 66 162 70
rect 170 66 172 70
rect 177 66 179 70
rect 79 43 81 46
rect 89 43 91 46
rect 99 43 101 46
rect 79 41 101 43
rect 79 39 81 41
rect 83 39 85 41
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 33 31 35
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 69 35 71 38
rect 79 37 85 39
rect 99 39 101 41
rect 109 39 111 42
rect 99 37 111 39
rect 79 35 81 37
rect 39 33 64 35
rect 9 26 11 33
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 58 31 60 33
rect 62 31 64 33
rect 58 29 64 31
rect 19 26 21 29
rect 42 25 44 29
rect 52 25 54 29
rect 62 25 64 29
rect 69 33 81 35
rect 69 25 71 33
rect 79 25 81 33
rect 89 34 95 36
rect 89 32 91 34
rect 93 32 95 34
rect 119 33 121 38
rect 126 35 128 38
rect 136 35 138 38
rect 126 33 138 35
rect 143 35 145 38
rect 153 35 155 38
rect 143 33 155 35
rect 86 30 95 32
rect 114 31 121 33
rect 86 25 88 30
rect 114 29 116 31
rect 118 29 121 31
rect 129 31 131 33
rect 133 31 135 33
rect 129 29 135 31
rect 114 27 121 29
rect 9 6 11 9
rect 19 6 21 9
rect 42 6 44 9
rect 52 6 54 9
rect 9 4 54 6
rect 62 4 64 9
rect 69 4 71 9
rect 79 4 81 9
rect 86 4 88 9
rect 133 23 135 29
rect 143 31 147 33
rect 149 31 155 33
rect 143 29 155 31
rect 160 35 162 38
rect 170 35 172 38
rect 160 33 172 35
rect 160 31 163 33
rect 165 31 167 33
rect 160 29 167 31
rect 143 23 145 29
rect 153 23 155 29
rect 163 23 165 29
rect 177 27 179 38
rect 177 25 183 27
rect 177 23 179 25
rect 181 23 183 25
rect 177 21 183 23
rect 133 2 135 6
rect 143 2 145 6
rect 153 2 155 6
rect 163 2 165 6
<< ndif >>
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 13 9 19
rect 2 11 4 13
rect 6 11 9 13
rect 2 9 9 11
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 11 15 14 17
rect 16 15 19 17
rect 11 9 19 15
rect 21 13 29 26
rect 21 11 24 13
rect 26 11 29 13
rect 35 23 42 25
rect 35 21 37 23
rect 39 21 42 23
rect 35 16 42 21
rect 35 14 37 16
rect 39 14 42 16
rect 35 12 42 14
rect 21 9 29 11
rect 37 9 42 12
rect 44 23 52 25
rect 44 21 47 23
rect 49 21 52 23
rect 44 9 52 21
rect 54 23 62 25
rect 54 21 57 23
rect 59 21 62 23
rect 54 16 62 21
rect 54 14 57 16
rect 59 14 62 16
rect 54 9 62 14
rect 64 9 69 25
rect 71 13 79 25
rect 71 11 74 13
rect 76 11 79 13
rect 71 9 79 11
rect 81 9 86 25
rect 88 23 95 25
rect 88 21 91 23
rect 93 21 95 23
rect 88 16 95 21
rect 88 14 91 16
rect 93 14 95 16
rect 88 12 95 14
rect 88 9 93 12
rect 124 17 133 23
rect 124 15 127 17
rect 129 15 133 17
rect 124 10 133 15
rect 124 8 127 10
rect 129 8 133 10
rect 124 6 133 8
rect 135 17 143 23
rect 135 15 138 17
rect 140 15 143 17
rect 135 6 143 15
rect 145 10 153 23
rect 145 8 148 10
rect 150 8 153 10
rect 145 6 153 8
rect 155 17 163 23
rect 155 15 158 17
rect 160 15 163 17
rect 155 6 163 15
rect 165 10 173 23
rect 165 8 168 10
rect 170 8 173 10
rect 165 6 173 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 50 19 66
rect 11 48 14 50
rect 16 48 19 50
rect 11 43 19 48
rect 11 41 14 43
rect 16 41 19 43
rect 11 38 19 41
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 50 39 55
rect 31 48 34 50
rect 36 48 39 50
rect 31 38 39 48
rect 41 58 49 66
rect 41 56 44 58
rect 46 56 49 58
rect 41 42 49 56
rect 41 40 44 42
rect 46 40 49 42
rect 41 38 49 40
rect 51 49 59 66
rect 51 47 54 49
rect 56 47 59 49
rect 51 42 59 47
rect 51 40 54 42
rect 56 40 59 42
rect 51 38 59 40
rect 61 58 69 66
rect 61 56 64 58
rect 66 56 69 58
rect 61 51 69 56
rect 61 49 64 51
rect 66 49 69 51
rect 61 38 69 49
rect 71 50 79 66
rect 71 48 74 50
rect 76 48 79 50
rect 71 46 79 48
rect 81 58 89 66
rect 81 56 84 58
rect 86 56 89 58
rect 81 46 89 56
rect 91 50 99 66
rect 91 48 94 50
rect 96 48 99 50
rect 91 46 99 48
rect 101 58 109 66
rect 101 56 104 58
rect 106 56 109 58
rect 101 46 109 56
rect 71 38 76 46
rect 104 42 109 46
rect 111 57 119 66
rect 111 55 114 57
rect 116 55 119 57
rect 111 50 119 55
rect 111 48 114 50
rect 116 48 119 50
rect 111 42 119 48
rect 114 38 119 42
rect 121 38 126 66
rect 128 64 136 66
rect 128 62 131 64
rect 133 62 136 64
rect 128 57 136 62
rect 128 55 131 57
rect 133 55 136 57
rect 128 38 136 55
rect 138 38 143 66
rect 145 57 153 66
rect 145 55 148 57
rect 150 55 153 57
rect 145 50 153 55
rect 145 48 148 50
rect 150 48 153 50
rect 145 38 153 48
rect 155 38 160 66
rect 162 64 170 66
rect 162 62 165 64
rect 167 62 170 64
rect 162 57 170 62
rect 162 55 165 57
rect 167 55 170 57
rect 162 38 170 55
rect 172 38 177 66
rect 179 51 184 66
rect 179 49 186 51
rect 179 47 182 49
rect 184 47 186 49
rect 179 42 186 47
rect 179 40 182 42
rect 184 40 186 42
rect 179 38 186 40
<< alu1 >>
rect -2 67 202 72
rect -2 65 190 67
rect 192 65 202 67
rect -2 64 202 65
rect 26 35 30 43
rect 18 33 30 35
rect 18 31 21 33
rect 23 31 30 33
rect 18 29 30 31
rect 26 21 30 29
rect 34 42 48 43
rect 34 40 44 42
rect 46 40 48 42
rect 34 38 48 40
rect 34 23 38 38
rect 129 38 167 42
rect 113 31 119 34
rect 34 21 37 23
rect 34 17 38 21
rect 113 29 116 31
rect 118 29 119 31
rect 129 33 135 38
rect 129 31 131 33
rect 133 31 135 33
rect 129 30 135 31
rect 113 26 119 29
rect 146 33 150 34
rect 146 31 147 33
rect 149 31 150 33
rect 146 26 150 31
rect 161 33 167 38
rect 161 31 163 33
rect 165 31 167 33
rect 161 30 167 31
rect 56 23 95 26
rect 56 21 57 23
rect 59 22 91 23
rect 59 21 61 22
rect 56 17 61 21
rect 34 16 61 17
rect 34 14 37 16
rect 39 14 57 16
rect 59 14 61 16
rect 89 21 91 22
rect 93 21 95 23
rect 89 16 95 21
rect 34 13 61 14
rect 89 14 91 16
rect 93 14 95 16
rect 113 25 183 26
rect 113 23 179 25
rect 181 23 183 25
rect 113 22 183 23
rect 113 14 119 22
rect 89 13 95 14
rect -2 7 202 8
rect -2 5 103 7
rect 105 5 189 7
rect 191 5 202 7
rect -2 0 202 5
<< ptie >>
rect 101 7 107 24
rect 101 5 103 7
rect 105 5 107 7
rect 187 7 193 24
rect 101 3 107 5
rect 187 5 189 7
rect 191 5 193 7
rect 187 3 193 5
<< ntie >>
rect 188 67 194 69
rect 188 65 190 67
rect 192 65 194 67
rect 188 59 194 65
rect 188 57 190 59
rect 192 57 194 59
rect 188 55 194 57
<< nmos >>
rect 9 9 11 26
rect 19 9 21 26
rect 42 9 44 25
rect 52 9 54 25
rect 62 9 64 25
rect 69 9 71 25
rect 79 9 81 25
rect 86 9 88 25
rect 133 6 135 23
rect 143 6 145 23
rect 153 6 155 23
rect 163 6 165 23
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 79 46 81 66
rect 89 46 91 66
rect 99 46 101 66
rect 109 42 111 66
rect 119 38 121 66
rect 126 38 128 66
rect 136 38 138 66
rect 143 38 145 66
rect 153 38 155 66
rect 160 38 162 66
rect 170 38 172 66
rect 177 38 179 66
<< polyct0 >>
rect 81 39 83 41
rect 60 31 62 33
rect 91 32 93 34
<< polyct1 >>
rect 21 31 23 33
rect 116 29 118 31
rect 131 31 133 33
rect 147 31 149 33
rect 163 31 165 33
rect 179 23 181 25
<< ndifct0 >>
rect 4 19 6 21
rect 4 11 6 13
rect 14 22 16 24
rect 14 15 16 17
rect 24 11 26 13
rect 38 21 39 23
rect 47 21 49 23
rect 74 11 76 13
rect 127 15 129 17
rect 127 8 129 10
rect 138 15 140 17
rect 148 8 150 10
rect 158 15 160 17
rect 168 8 170 10
<< ndifct1 >>
rect 37 21 38 23
rect 37 14 39 16
rect 57 21 59 23
rect 57 14 59 16
rect 91 21 93 23
rect 91 14 93 16
<< ntiect0 >>
rect 190 57 192 59
<< ntiect1 >>
rect 190 65 192 67
<< ptiect1 >>
rect 103 5 105 7
rect 189 5 191 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 48 16 50
rect 14 41 16 43
rect 24 62 26 64
rect 24 55 26 57
rect 34 55 36 57
rect 34 48 36 50
rect 44 56 46 58
rect 54 47 56 49
rect 54 40 56 42
rect 64 56 66 58
rect 64 49 66 51
rect 74 48 76 50
rect 84 56 86 58
rect 94 48 96 50
rect 104 56 106 58
rect 114 55 116 57
rect 114 48 116 50
rect 131 62 133 64
rect 131 55 133 57
rect 148 55 150 57
rect 148 48 150 50
rect 165 62 167 64
rect 165 55 167 57
rect 182 47 184 49
rect 182 40 184 42
<< pdifct1 >>
rect 44 40 46 42
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 22 62 24 64
rect 26 62 28 64
rect 22 57 28 62
rect 129 62 131 64
rect 133 62 135 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 33 57 37 59
rect 33 55 34 57
rect 36 55 37 57
rect 42 58 108 59
rect 42 56 44 58
rect 46 56 64 58
rect 66 56 84 58
rect 86 56 104 58
rect 106 56 108 58
rect 42 55 108 56
rect 113 57 117 59
rect 113 55 114 57
rect 116 55 117 57
rect 33 51 37 55
rect 63 51 67 55
rect 113 51 117 55
rect 129 57 135 62
rect 163 62 165 64
rect 167 62 169 64
rect 129 55 131 57
rect 133 55 135 57
rect 129 54 135 55
rect 147 57 151 59
rect 147 55 148 57
rect 150 55 151 57
rect 147 51 151 55
rect 163 57 169 62
rect 163 55 165 57
rect 167 55 169 57
rect 189 59 193 64
rect 189 57 190 59
rect 192 57 193 59
rect 189 55 193 57
rect 163 54 169 55
rect 12 50 57 51
rect 12 48 14 50
rect 16 48 34 50
rect 36 49 57 50
rect 36 48 54 49
rect 12 47 54 48
rect 56 47 57 49
rect 63 49 64 51
rect 66 49 67 51
rect 63 47 67 49
rect 72 50 185 51
rect 72 48 74 50
rect 76 48 94 50
rect 96 48 114 50
rect 116 48 148 50
rect 150 49 185 50
rect 150 48 182 49
rect 72 47 182 48
rect 184 47 185 49
rect 12 43 17 47
rect 10 41 14 43
rect 16 41 17 43
rect 10 39 17 41
rect 10 25 14 39
rect 10 24 18 25
rect 3 21 7 23
rect 10 22 14 24
rect 16 22 18 24
rect 10 21 18 22
rect 53 42 57 47
rect 53 40 54 42
rect 56 41 85 42
rect 56 40 81 41
rect 53 39 81 40
rect 83 39 85 41
rect 53 38 85 39
rect 90 34 94 47
rect 181 42 185 47
rect 181 40 182 42
rect 184 40 190 42
rect 181 38 190 40
rect 45 33 91 34
rect 45 31 60 33
rect 62 32 91 33
rect 93 32 94 34
rect 62 31 94 32
rect 45 30 94 31
rect 38 23 40 25
rect 39 21 40 23
rect 3 19 4 21
rect 6 19 7 21
rect 3 13 7 19
rect 12 17 18 21
rect 12 15 14 17
rect 16 15 18 17
rect 38 17 40 21
rect 45 23 51 30
rect 145 26 146 34
rect 150 26 151 34
rect 45 21 47 23
rect 49 21 51 23
rect 45 20 51 21
rect 12 14 18 15
rect 3 11 4 13
rect 6 11 7 13
rect 3 8 7 11
rect 23 13 27 15
rect 73 13 77 15
rect 126 17 130 19
rect 186 18 190 38
rect 126 15 127 17
rect 129 15 130 17
rect 23 11 24 13
rect 26 11 27 13
rect 23 8 27 11
rect 73 11 74 13
rect 76 11 77 13
rect 73 8 77 11
rect 126 10 130 15
rect 136 17 190 18
rect 136 15 138 17
rect 140 15 158 17
rect 160 15 190 17
rect 136 14 190 15
rect 126 8 127 10
rect 129 8 130 10
rect 146 10 152 11
rect 146 8 148 10
rect 150 8 152 10
rect 166 10 172 11
rect 166 8 168 10
rect 170 8 172 10
<< labels >>
rlabel alu0 15 19 15 19 6 bn
rlabel alu0 14 45 14 45 6 bn
rlabel alu0 35 53 35 53 6 bn
rlabel alu0 48 27 48 27 6 an
rlabel alu0 69 40 69 40 6 bn
rlabel alu0 55 44 55 44 6 bn
rlabel alu0 34 49 34 49 6 bn
rlabel alu0 115 53 115 53 6 an
rlabel alu0 163 16 163 16 6 an
rlabel alu0 183 44 183 44 6 an
rlabel alu0 128 49 128 49 6 an
rlabel alu0 149 53 149 53 6 an
rlabel alu1 20 32 20 32 6 b
rlabel alu1 28 32 28 32 6 b
rlabel alu1 60 24 60 24 6 z
rlabel alu1 68 24 68 24 6 z
rlabel alu1 76 24 76 24 6 z
rlabel alu1 36 28 36 28 6 z
rlabel alu1 44 40 44 40 6 z
rlabel alu1 100 4 100 4 6 vss
rlabel alu1 116 24 116 24 6 a2
rlabel alu1 84 24 84 24 6 z
rlabel alu1 92 20 92 20 6 z
rlabel alu1 100 68 100 68 6 vdd
rlabel alu1 124 24 124 24 6 a2
rlabel alu1 132 24 132 24 6 a2
rlabel alu1 140 24 140 24 6 a2
rlabel alu1 156 24 156 24 6 a2
rlabel alu1 148 28 148 28 6 a2
rlabel alu1 140 40 140 40 6 a1
rlabel alu1 148 40 148 40 6 a1
rlabel alu1 156 40 156 40 6 a1
rlabel alu1 132 36 132 36 6 a1
rlabel alu1 164 24 164 24 6 a2
rlabel alu1 172 24 172 24 6 a2
rlabel polyct1 180 24 180 24 6 a2
rlabel alu1 164 36 164 36 6 a1
rlabel alu1 164 40 164 40 6 a1
<< end >>
