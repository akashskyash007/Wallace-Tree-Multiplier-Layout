magic
tech scmos
timestamp 1199202788
<< ab >>
rect 0 0 88 72
<< nwell >>
rect -5 32 93 77
<< pwell >>
rect -5 -5 93 32
<< poly >>
rect 25 66 27 70
rect 35 66 37 70
rect 47 66 49 70
rect 57 66 59 70
rect 67 66 69 70
rect 77 66 79 70
rect 15 58 17 63
rect 15 43 17 46
rect 11 41 17 43
rect 11 39 13 41
rect 15 39 17 41
rect 11 37 21 39
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 9 27 15 29
rect 12 24 14 27
rect 19 24 21 37
rect 25 35 27 43
rect 47 44 49 47
rect 44 42 50 44
rect 44 40 46 42
rect 48 40 50 42
rect 77 44 79 47
rect 77 42 86 44
rect 35 35 37 39
rect 44 38 50 40
rect 57 38 59 41
rect 67 38 69 41
rect 25 33 37 35
rect 25 31 33 33
rect 35 31 37 33
rect 25 29 41 31
rect 26 24 28 29
rect 39 24 41 29
rect 46 24 48 38
rect 57 36 69 38
rect 77 40 82 42
rect 84 40 86 42
rect 77 38 86 40
rect 77 36 79 38
rect 60 31 66 36
rect 73 34 79 36
rect 73 32 75 34
rect 60 29 62 31
rect 64 29 66 31
rect 53 27 66 29
rect 70 30 75 32
rect 53 24 55 27
rect 63 20 65 27
rect 70 20 72 30
rect 79 27 85 29
rect 79 26 81 27
rect 77 25 81 26
rect 83 25 85 27
rect 77 23 85 25
rect 77 20 79 23
rect 12 2 14 6
rect 19 2 21 6
rect 26 2 28 6
rect 39 2 41 6
rect 46 2 48 6
rect 53 2 55 6
rect 63 2 65 6
rect 70 2 72 6
rect 77 2 79 6
<< ndif >>
rect 7 19 12 24
rect 5 17 12 19
rect 5 15 7 17
rect 9 15 12 17
rect 5 13 12 15
rect 7 6 12 13
rect 14 6 19 24
rect 21 6 26 24
rect 28 10 39 24
rect 28 8 32 10
rect 34 8 39 10
rect 28 6 39 8
rect 41 6 46 24
rect 48 6 53 24
rect 55 20 60 24
rect 55 17 63 20
rect 55 15 58 17
rect 60 15 63 17
rect 55 6 63 15
rect 65 6 70 20
rect 72 6 77 20
rect 79 17 86 20
rect 79 15 82 17
rect 84 15 86 17
rect 79 10 86 15
rect 79 8 82 10
rect 84 8 86 10
rect 79 6 86 8
<< pdif >>
rect 19 58 25 66
rect 10 52 15 58
rect 8 50 15 52
rect 8 48 10 50
rect 12 48 15 50
rect 8 46 15 48
rect 17 56 25 58
rect 17 54 20 56
rect 22 54 25 56
rect 17 46 25 54
rect 19 43 25 46
rect 27 56 35 66
rect 27 54 30 56
rect 32 54 35 56
rect 27 49 35 54
rect 27 47 30 49
rect 32 47 35 49
rect 27 43 35 47
rect 30 39 35 43
rect 37 64 47 66
rect 37 62 41 64
rect 43 62 47 64
rect 37 47 47 62
rect 49 57 57 66
rect 49 55 52 57
rect 54 55 57 57
rect 49 47 57 55
rect 37 39 42 47
rect 52 41 57 47
rect 59 64 67 66
rect 59 62 62 64
rect 64 62 67 64
rect 59 41 67 62
rect 69 57 77 66
rect 69 55 72 57
rect 74 55 77 57
rect 69 47 77 55
rect 79 64 86 66
rect 79 62 82 64
rect 84 62 86 64
rect 79 47 86 62
rect 69 41 74 47
<< alu1 >>
rect -2 67 90 72
rect -2 65 5 67
rect 7 65 90 67
rect -2 64 90 65
rect 29 57 79 58
rect 29 56 52 57
rect 29 54 30 56
rect 32 55 52 56
rect 54 55 72 57
rect 74 55 79 57
rect 32 54 79 55
rect 2 50 14 51
rect 29 50 34 54
rect 2 48 10 50
rect 12 49 34 50
rect 12 48 30 49
rect 2 47 30 48
rect 32 47 34 49
rect 2 46 34 47
rect 45 46 86 50
rect 2 18 6 46
rect 45 42 49 46
rect 11 41 46 42
rect 11 39 13 41
rect 15 40 46 41
rect 48 40 49 42
rect 15 39 49 40
rect 11 38 49 39
rect 53 38 78 42
rect 82 42 86 46
rect 84 40 86 42
rect 53 34 57 38
rect 17 26 23 34
rect 31 33 57 34
rect 31 31 33 33
rect 35 31 57 33
rect 31 30 57 31
rect 61 31 65 33
rect 61 29 62 31
rect 64 29 65 31
rect 61 26 65 29
rect 17 22 65 26
rect 74 21 78 38
rect 82 37 86 40
rect 2 17 63 18
rect 2 15 7 17
rect 9 15 58 17
rect 60 15 63 17
rect 2 14 63 15
rect -2 0 90 8
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 12 6 14 24
rect 19 6 21 24
rect 26 6 28 24
rect 39 6 41 24
rect 46 6 48 24
rect 53 6 55 24
rect 63 6 65 20
rect 70 6 72 20
rect 77 6 79 20
<< pmos >>
rect 15 46 17 58
rect 25 43 27 66
rect 35 39 37 66
rect 47 47 49 66
rect 57 41 59 66
rect 67 41 69 66
rect 77 47 79 66
<< polyct0 >>
rect 11 29 13 31
rect 81 25 83 27
<< polyct1 >>
rect 13 39 15 41
rect 46 40 48 42
rect 33 31 35 33
rect 82 40 84 42
rect 62 29 64 31
<< ndifct0 >>
rect 32 8 34 10
rect 82 15 84 17
rect 82 8 84 10
<< ndifct1 >>
rect 7 15 9 17
rect 58 15 60 17
<< ntiect1 >>
rect 5 65 7 67
<< pdifct0 >>
rect 20 54 22 56
rect 41 62 43 64
rect 62 62 64 64
rect 82 62 84 64
<< pdifct1 >>
rect 10 48 12 50
rect 30 54 32 56
rect 30 47 32 49
rect 52 55 54 57
rect 72 55 74 57
<< alu0 >>
rect 18 56 24 64
rect 39 62 41 64
rect 43 62 45 64
rect 39 61 45 62
rect 60 62 62 64
rect 64 62 66 64
rect 60 61 66 62
rect 80 62 82 64
rect 84 62 86 64
rect 80 61 86 62
rect 18 54 20 56
rect 22 54 24 56
rect 18 53 24 54
rect 81 38 82 46
rect 10 31 17 33
rect 10 29 11 31
rect 13 29 17 31
rect 10 27 17 29
rect 78 27 85 28
rect 78 25 81 27
rect 83 25 85 27
rect 78 24 85 25
rect 80 17 86 18
rect 80 15 82 17
rect 84 15 86 17
rect 30 10 36 11
rect 30 8 32 10
rect 34 8 36 10
rect 80 10 86 15
rect 80 8 82 10
rect 84 8 86 10
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 28 24 28 24 6 c
rlabel alu1 20 28 20 28 6 c
rlabel alu1 20 40 20 40 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 44 4 44 4 6 vss
rlabel alu1 44 16 44 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 36 24 36 24 6 c
rlabel alu1 44 24 44 24 6 c
rlabel alu1 44 32 44 32 6 a
rlabel alu1 36 32 36 32 6 a
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 44 56 44 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 44 68 44 68 6 vdd
rlabel alu1 60 16 60 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 52 24 52 24 6 c
rlabel alu1 60 24 60 24 6 c
rlabel alu1 52 32 52 32 6 a
rlabel alu1 60 40 60 40 6 a
rlabel alu1 68 40 68 40 6 a
rlabel alu1 52 48 52 48 6 b
rlabel alu1 60 48 60 48 6 b
rlabel alu1 68 48 68 48 6 b
rlabel alu1 60 56 60 56 6 z
rlabel alu1 68 56 68 56 6 z
rlabel alu1 52 56 52 56 6 z
rlabel alu1 76 28 76 28 6 a
rlabel alu1 84 40 84 40 6 b
rlabel alu1 76 48 76 48 6 b
rlabel alu1 76 56 76 56 6 z
<< end >>
