magic
tech scmos
timestamp 1199203260
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 24 70 26 74
rect 31 70 33 74
rect 38 70 40 74
rect 13 61 15 66
rect 13 39 15 42
rect 24 39 26 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 26 39
rect 19 35 21 37
rect 23 36 26 37
rect 23 35 25 36
rect 19 33 25 35
rect 9 25 11 33
rect 19 22 21 33
rect 31 31 33 42
rect 38 39 40 42
rect 38 37 46 39
rect 40 35 42 37
rect 44 35 46 37
rect 40 33 46 35
rect 29 29 36 31
rect 29 27 32 29
rect 34 27 36 29
rect 29 25 36 27
rect 29 22 31 25
rect 41 22 43 33
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 41 11 43 16
<< ndif >>
rect 4 22 9 25
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 22 17 25
rect 11 20 19 22
rect 11 18 14 20
rect 16 18 19 20
rect 11 16 19 18
rect 21 20 29 22
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 31 16 41 22
rect 43 20 50 22
rect 43 18 46 20
rect 48 18 50 20
rect 43 16 50 18
rect 33 11 39 16
rect 33 9 35 11
rect 37 9 39 11
rect 33 7 39 9
<< pdif >>
rect 17 64 24 70
rect 17 62 19 64
rect 21 62 24 64
rect 17 61 24 62
rect 6 59 13 61
rect 6 57 8 59
rect 10 57 13 59
rect 6 55 13 57
rect 8 42 13 55
rect 15 42 24 61
rect 26 42 31 70
rect 33 42 38 70
rect 40 64 45 70
rect 40 62 47 64
rect 40 60 43 62
rect 45 60 47 62
rect 40 58 47 60
rect 40 42 45 58
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 59 15 62
rect 2 57 8 59
rect 10 57 15 59
rect 2 56 15 57
rect 2 21 6 56
rect 34 49 46 55
rect 26 39 30 47
rect 42 41 46 49
rect 17 37 30 39
rect 17 35 21 37
rect 23 35 30 37
rect 17 34 30 35
rect 34 30 38 39
rect 30 29 47 30
rect 30 27 32 29
rect 34 27 47 29
rect 30 26 47 27
rect 2 20 8 21
rect 2 18 4 20
rect 6 18 8 20
rect 2 17 8 18
rect -2 11 58 12
rect -2 9 35 11
rect 37 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 16 11 25
rect 19 16 21 22
rect 29 16 31 22
rect 41 16 43 22
<< pmos >>
rect 13 42 15 61
rect 24 42 26 70
rect 31 42 33 70
rect 38 42 40 70
<< polyct0 >>
rect 11 35 13 37
rect 42 35 44 37
<< polyct1 >>
rect 21 35 23 37
rect 32 27 34 29
<< ndifct0 >>
rect 14 18 16 20
rect 24 18 26 20
rect 46 18 48 20
<< ndifct1 >>
rect 4 18 6 20
rect 35 9 37 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 19 62 21 64
rect 43 60 45 62
<< pdifct1 >>
rect 8 57 10 59
<< alu0 >>
rect 18 64 22 68
rect 18 62 19 64
rect 21 62 22 64
rect 18 60 22 62
rect 26 62 47 63
rect 26 60 43 62
rect 45 60 47 62
rect 26 59 47 60
rect 26 55 30 59
rect 18 51 30 55
rect 18 48 22 51
rect 10 44 22 48
rect 10 37 14 44
rect 41 41 42 49
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 41 37 45 41
rect 41 35 42 37
rect 44 35 45 37
rect 41 33 45 35
rect 10 25 26 29
rect 22 21 26 25
rect 12 20 18 21
rect 12 18 14 20
rect 16 18 18 20
rect 12 12 18 18
rect 22 20 50 21
rect 22 18 24 20
rect 26 18 46 20
rect 48 18 50 20
rect 22 17 50 18
<< labels >>
rlabel polyct0 12 36 12 36 6 zn
rlabel alu0 36 19 36 19 6 zn
rlabel alu0 36 61 36 61 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 36 20 36 6 a
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 32 36 32 6 b
rlabel alu1 28 44 28 44 6 a
rlabel alu1 36 52 36 52 6 c
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 b
rlabel alu1 44 48 44 48 6 c
<< end >>
