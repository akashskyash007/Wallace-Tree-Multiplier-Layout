magic
tech scmos
timestamp 1199203416
<< ab >>
rect 0 0 152 80
<< nwell >>
rect -5 36 157 88
<< pwell >>
rect -5 -8 157 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 51 70 53 74
rect 58 70 60 74
rect 68 70 70 74
rect 78 70 80 74
rect 88 70 90 74
rect 95 70 97 74
rect 111 70 113 74
rect 121 70 123 74
rect 131 70 133 74
rect 141 70 143 74
rect 35 45 41 47
rect 35 43 37 45
rect 39 43 41 45
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 21 39
rect 9 35 17 37
rect 19 35 21 37
rect 35 39 41 43
rect 51 39 53 42
rect 35 37 53 39
rect 35 35 41 37
rect 9 33 21 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 33 41 35
rect 29 30 31 33
rect 39 30 41 33
rect 58 30 60 42
rect 68 39 70 42
rect 78 39 80 42
rect 64 37 80 39
rect 88 39 90 42
rect 95 39 97 42
rect 111 39 113 42
rect 121 39 123 42
rect 131 39 133 42
rect 64 35 66 37
rect 68 35 70 37
rect 88 36 91 39
rect 95 37 107 39
rect 64 33 70 35
rect 54 28 60 30
rect 79 28 81 33
rect 89 30 91 36
rect 101 35 103 37
rect 105 35 107 37
rect 101 33 107 35
rect 111 37 117 39
rect 111 35 113 37
rect 115 35 117 37
rect 111 33 117 35
rect 121 37 133 39
rect 121 35 123 37
rect 125 35 133 37
rect 141 39 143 42
rect 141 37 150 39
rect 141 35 146 37
rect 148 35 150 37
rect 121 33 133 35
rect 114 30 116 33
rect 121 30 123 33
rect 131 30 133 33
rect 138 33 150 35
rect 138 30 140 33
rect 54 26 56 28
rect 58 26 60 28
rect 54 24 70 26
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 39 11 41 16
rect 68 8 70 24
rect 79 8 81 11
rect 89 8 91 11
rect 68 6 91 8
rect 114 7 116 12
rect 121 7 123 12
rect 131 7 133 12
rect 138 7 140 12
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 16 9 19
rect 11 20 19 30
rect 11 18 14 20
rect 16 18 19 20
rect 11 16 19 18
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 21 29 26
rect 21 19 24 21
rect 26 19 29 21
rect 21 16 29 19
rect 31 21 39 30
rect 31 19 34 21
rect 36 19 39 21
rect 31 16 39 19
rect 41 28 48 30
rect 41 26 44 28
rect 46 26 48 28
rect 41 24 48 26
rect 84 28 89 30
rect 41 16 46 24
rect 74 23 79 28
rect 72 21 79 23
rect 72 19 74 21
rect 76 19 79 21
rect 72 17 79 19
rect 74 11 79 17
rect 81 20 89 28
rect 81 18 84 20
rect 86 18 89 20
rect 81 11 89 18
rect 91 28 98 30
rect 91 26 94 28
rect 96 26 98 28
rect 91 24 98 26
rect 91 11 96 24
rect 105 12 114 30
rect 116 12 121 30
rect 123 20 131 30
rect 123 18 126 20
rect 128 18 131 20
rect 123 12 131 18
rect 133 12 138 30
rect 140 25 148 30
rect 140 23 143 25
rect 145 23 148 25
rect 140 17 148 23
rect 140 15 143 17
rect 145 15 148 17
rect 140 12 148 15
rect 105 11 112 12
rect 105 9 108 11
rect 110 9 112 11
rect 105 7 112 9
<< pdif >>
rect 99 70 109 72
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 60 9 66
rect 2 58 4 60
rect 6 58 9 60
rect 2 42 9 58
rect 11 54 19 70
rect 11 52 14 54
rect 16 52 19 54
rect 11 47 19 52
rect 11 45 14 47
rect 16 45 19 47
rect 11 42 19 45
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 43 68 51 70
rect 43 66 46 68
rect 48 66 51 68
rect 43 61 51 66
rect 43 59 46 61
rect 48 59 51 61
rect 43 42 51 59
rect 53 42 58 70
rect 60 46 68 70
rect 60 44 63 46
rect 65 44 68 46
rect 60 42 68 44
rect 70 61 78 70
rect 70 59 73 61
rect 75 59 78 61
rect 70 54 78 59
rect 70 52 73 54
rect 75 52 78 54
rect 70 42 78 52
rect 80 46 88 70
rect 80 44 83 46
rect 85 44 88 46
rect 80 42 88 44
rect 90 42 95 70
rect 97 69 111 70
rect 97 67 103 69
rect 105 67 111 69
rect 97 62 111 67
rect 97 60 103 62
rect 105 60 111 62
rect 97 42 111 60
rect 113 61 121 70
rect 113 59 116 61
rect 118 59 121 61
rect 113 54 121 59
rect 113 52 116 54
rect 118 52 121 54
rect 113 42 121 52
rect 123 68 131 70
rect 123 66 126 68
rect 128 66 131 68
rect 123 61 131 66
rect 123 59 126 61
rect 128 59 131 61
rect 123 42 131 59
rect 133 61 141 70
rect 133 59 136 61
rect 138 59 141 61
rect 133 54 141 59
rect 133 52 136 54
rect 138 52 141 54
rect 133 42 141 52
rect 143 68 150 70
rect 143 66 146 68
rect 148 66 150 68
rect 143 61 150 66
rect 143 59 146 61
rect 148 59 150 61
rect 143 42 150 59
<< alu1 >>
rect -2 81 154 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 154 81
rect -2 69 154 79
rect -2 68 103 69
rect 105 68 154 69
rect 26 38 30 55
rect 57 46 87 47
rect 57 44 63 46
rect 65 44 83 46
rect 85 44 87 46
rect 57 42 87 44
rect 15 37 71 38
rect 15 35 17 37
rect 19 35 66 37
rect 68 35 71 37
rect 15 34 71 35
rect 82 30 87 42
rect 146 46 150 55
rect 73 28 98 30
rect 73 26 94 28
rect 96 26 98 28
rect 73 25 98 26
rect 73 22 78 25
rect 32 21 78 22
rect 111 42 150 46
rect 111 37 117 42
rect 111 35 113 37
rect 115 35 117 37
rect 111 34 117 35
rect 121 37 127 38
rect 121 35 123 37
rect 125 35 127 37
rect 121 30 127 35
rect 145 37 150 42
rect 145 35 146 37
rect 148 35 150 37
rect 145 33 150 35
rect 121 26 135 30
rect 32 19 34 21
rect 36 19 74 21
rect 76 19 78 21
rect 32 18 78 19
rect -2 11 154 12
rect -2 9 108 11
rect 110 9 154 11
rect -2 1 154 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 154 1
rect -2 -2 154 -1
<< ptie >>
rect 0 1 152 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 152 1
rect 0 -3 152 -1
<< ntie >>
rect 0 81 152 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 152 81
rect 0 77 152 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 30
rect 39 16 41 30
rect 79 11 81 28
rect 89 11 91 30
rect 114 12 116 30
rect 121 12 123 30
rect 131 12 133 30
rect 138 12 140 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 51 42 53 70
rect 58 42 60 70
rect 68 42 70 70
rect 78 42 80 70
rect 88 42 90 70
rect 95 42 97 70
rect 111 42 113 70
rect 121 42 123 70
rect 131 42 133 70
rect 141 42 143 70
<< polyct0 >>
rect 37 43 39 45
rect 103 35 105 37
rect 56 26 58 28
<< polyct1 >>
rect 17 35 19 37
rect 66 35 68 37
rect 113 35 115 37
rect 123 35 125 37
rect 146 35 148 37
<< ndifct0 >>
rect 4 26 6 28
rect 4 19 6 21
rect 14 18 16 20
rect 24 26 26 28
rect 24 19 26 21
rect 44 26 46 28
rect 84 18 86 20
rect 126 18 128 20
rect 143 23 145 25
rect 143 15 145 17
<< ndifct1 >>
rect 34 19 36 21
rect 74 19 76 21
rect 94 26 96 28
rect 108 9 110 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 58 6 60
rect 14 52 16 54
rect 14 45 16 47
rect 24 66 26 68
rect 24 59 26 61
rect 46 66 48 68
rect 46 59 48 61
rect 73 59 75 61
rect 73 52 75 54
rect 103 67 105 68
rect 103 60 105 62
rect 116 59 118 61
rect 116 52 118 54
rect 126 66 128 68
rect 126 59 128 61
rect 136 59 138 61
rect 136 52 138 54
rect 146 66 148 68
rect 146 59 148 61
<< pdifct1 >>
rect 63 44 65 46
rect 83 44 85 46
rect 103 68 105 69
<< alu0 >>
rect 3 66 4 68
rect 6 66 7 68
rect 3 60 7 66
rect 3 58 4 60
rect 6 58 7 60
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 44 66 46 68
rect 48 66 50 68
rect 44 61 50 66
rect 101 67 103 68
rect 105 67 107 68
rect 44 59 46 61
rect 48 59 50 61
rect 44 58 50 59
rect 72 61 76 63
rect 72 59 73 61
rect 75 59 76 61
rect 101 62 107 67
rect 124 66 126 68
rect 128 66 130 68
rect 101 60 103 62
rect 105 60 107 62
rect 101 59 107 60
rect 115 61 119 63
rect 115 59 116 61
rect 118 59 119 61
rect 3 56 7 58
rect 13 54 17 56
rect 72 55 76 59
rect 115 55 119 59
rect 124 61 130 66
rect 144 66 146 68
rect 148 66 150 68
rect 124 59 126 61
rect 128 59 130 61
rect 124 58 130 59
rect 135 61 140 63
rect 135 59 136 61
rect 138 59 140 61
rect 135 55 140 59
rect 144 61 150 66
rect 144 59 146 61
rect 148 59 150 61
rect 144 58 150 59
rect 13 52 14 54
rect 16 52 17 54
rect 13 47 17 52
rect 2 45 14 47
rect 16 45 17 47
rect 2 43 17 45
rect 2 29 6 43
rect 46 54 140 55
rect 46 52 73 54
rect 75 52 116 54
rect 118 52 136 54
rect 138 52 140 54
rect 46 51 140 52
rect 46 46 50 51
rect 35 45 50 46
rect 35 43 37 45
rect 39 43 50 45
rect 35 42 50 43
rect 102 37 106 51
rect 102 35 103 37
rect 105 35 106 37
rect 2 28 60 29
rect 2 26 4 28
rect 6 26 24 28
rect 26 26 44 28
rect 46 26 56 28
rect 58 26 60 28
rect 2 25 60 26
rect 3 21 7 25
rect 23 21 27 25
rect 3 19 4 21
rect 6 19 7 21
rect 3 17 7 19
rect 12 20 18 21
rect 12 18 14 20
rect 16 18 18 20
rect 12 12 18 18
rect 23 19 24 21
rect 26 19 27 21
rect 23 17 27 19
rect 102 21 106 35
rect 142 25 146 27
rect 142 23 143 25
rect 145 23 146 25
rect 82 20 130 21
rect 82 18 84 20
rect 86 18 126 20
rect 128 18 130 20
rect 82 17 130 18
rect 142 17 146 23
rect 142 15 143 17
rect 145 15 146 17
rect 142 12 146 15
<< labels >>
rlabel alu0 25 23 25 23 6 bn
rlabel alu0 5 23 5 23 6 bn
rlabel alu0 15 49 15 49 6 bn
rlabel alu0 31 27 31 27 6 bn
rlabel alu0 42 44 42 44 6 an
rlabel alu0 74 57 74 57 6 an
rlabel polyct0 104 36 104 36 6 an
rlabel alu0 117 57 117 57 6 an
rlabel alu0 106 19 106 19 6 an
rlabel alu0 93 53 93 53 6 an
rlabel alu0 137 57 137 57 6 an
rlabel alu1 20 36 20 36 6 b
rlabel alu1 36 20 36 20 6 z
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 28 44 28 44 6 b
rlabel alu1 36 36 36 36 6 b
rlabel alu1 44 36 44 36 6 b
rlabel alu1 52 36 52 36 6 b
rlabel alu1 76 6 76 6 6 vss
rlabel alu1 60 20 60 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 76 28 76 28 6 z
rlabel alu1 60 36 60 36 6 b
rlabel alu1 60 44 60 44 6 z
rlabel alu1 68 36 68 36 6 b
rlabel alu1 68 44 68 44 6 z
rlabel alu1 76 44 76 44 6 z
rlabel alu1 84 36 84 36 6 z
rlabel alu1 76 74 76 74 6 vdd
rlabel alu1 92 28 92 28 6 z
rlabel alu1 116 44 116 44 6 a1
rlabel alu1 132 28 132 28 6 a2
rlabel alu1 124 32 124 32 6 a2
rlabel alu1 124 44 124 44 6 a1
rlabel alu1 148 44 148 44 6 a1
rlabel alu1 132 44 132 44 6 a1
rlabel alu1 140 44 140 44 6 a1
<< end >>
