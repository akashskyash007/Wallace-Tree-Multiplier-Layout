magic
tech scmos
timestamp 1199201918
<< ab >>
rect 0 0 144 80
<< nwell >>
rect -5 36 149 88
<< pwell >>
rect -5 -8 149 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 99 70 101 74
rect 109 70 111 74
rect 119 70 121 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 31 39
rect 9 35 11 37
rect 13 35 21 37
rect 9 33 21 35
rect 19 27 21 33
rect 29 27 31 37
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 39 37 61 39
rect 39 35 45 37
rect 47 35 57 37
rect 59 35 61 37
rect 39 33 61 35
rect 39 30 41 33
rect 49 30 51 33
rect 59 30 61 33
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 69 37 91 39
rect 69 35 77 37
rect 79 35 85 37
rect 87 35 91 37
rect 69 33 91 35
rect 69 30 71 33
rect 79 30 81 33
rect 89 30 91 33
rect 99 39 101 42
rect 109 39 111 42
rect 119 39 121 42
rect 99 37 121 39
rect 99 30 101 37
rect 108 35 110 37
rect 112 35 117 37
rect 119 35 121 37
rect 108 33 121 35
rect 109 30 111 33
rect 119 30 121 33
rect 19 11 21 16
rect 29 11 31 16
rect 39 7 41 12
rect 49 7 51 12
rect 59 7 61 12
rect 69 7 71 12
rect 79 7 81 12
rect 89 7 91 12
rect 99 7 101 12
rect 109 7 111 12
rect 119 7 121 12
<< ndif >>
rect 34 27 39 30
rect 12 25 19 27
rect 12 23 14 25
rect 16 23 19 25
rect 12 21 19 23
rect 14 16 19 21
rect 21 20 29 27
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 31 25 39 27
rect 31 23 34 25
rect 36 23 39 25
rect 31 16 39 23
rect 34 12 39 16
rect 41 20 49 30
rect 41 18 44 20
rect 46 18 49 20
rect 41 12 49 18
rect 51 28 59 30
rect 51 26 54 28
rect 56 26 59 28
rect 51 12 59 26
rect 61 27 69 30
rect 61 25 64 27
rect 66 25 69 27
rect 61 20 69 25
rect 61 18 64 20
rect 66 18 69 20
rect 61 12 69 18
rect 71 28 79 30
rect 71 26 74 28
rect 76 26 79 28
rect 71 12 79 26
rect 81 20 89 30
rect 81 18 84 20
rect 86 18 89 20
rect 81 12 89 18
rect 91 28 99 30
rect 91 26 94 28
rect 96 26 99 28
rect 91 21 99 26
rect 91 19 94 21
rect 96 19 99 21
rect 91 12 99 19
rect 101 16 109 30
rect 101 14 104 16
rect 106 14 109 16
rect 101 12 109 14
rect 111 28 119 30
rect 111 26 114 28
rect 116 26 119 28
rect 111 21 119 26
rect 111 19 114 21
rect 116 19 119 21
rect 111 12 119 19
rect 121 24 128 30
rect 121 22 124 24
rect 126 22 128 24
rect 121 16 128 22
rect 121 14 124 16
rect 126 14 128 16
rect 121 12 128 14
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 42 39 52
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 61 49 66
rect 41 59 44 61
rect 46 59 49 61
rect 41 42 49 59
rect 51 53 59 70
rect 51 51 54 53
rect 56 51 59 53
rect 51 46 59 51
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 68 69 70
rect 61 66 64 68
rect 66 66 69 68
rect 61 61 69 66
rect 61 59 64 61
rect 66 59 69 61
rect 61 42 69 59
rect 71 53 79 70
rect 71 51 74 53
rect 76 51 79 53
rect 71 46 79 51
rect 71 44 74 46
rect 76 44 79 46
rect 71 42 79 44
rect 81 68 89 70
rect 81 66 84 68
rect 86 66 89 68
rect 81 61 89 66
rect 81 59 84 61
rect 86 59 89 61
rect 81 42 89 59
rect 91 53 99 70
rect 91 51 94 53
rect 96 51 99 53
rect 91 46 99 51
rect 91 44 94 46
rect 96 44 99 46
rect 91 42 99 44
rect 101 68 109 70
rect 101 66 104 68
rect 106 66 109 68
rect 101 61 109 66
rect 101 59 104 61
rect 106 59 109 61
rect 101 42 109 59
rect 111 61 119 70
rect 111 59 114 61
rect 116 59 119 61
rect 111 54 119 59
rect 111 52 114 54
rect 116 52 119 54
rect 111 42 119 52
rect 121 68 128 70
rect 121 66 124 68
rect 126 66 128 68
rect 121 61 128 66
rect 121 59 124 61
rect 126 59 128 61
rect 121 42 128 59
<< alu1 >>
rect -2 81 146 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 146 81
rect -2 68 146 79
rect 2 53 7 63
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 24 46
rect 26 44 30 46
rect 2 42 30 44
rect 2 37 15 38
rect 2 35 11 37
rect 13 35 15 37
rect 2 34 15 35
rect 2 17 6 34
rect 26 30 30 42
rect 41 38 47 46
rect 81 38 87 46
rect 122 38 127 55
rect 41 37 63 38
rect 41 35 45 37
rect 47 35 57 37
rect 59 35 63 37
rect 41 34 63 35
rect 73 37 95 38
rect 73 35 77 37
rect 79 35 85 37
rect 87 35 95 37
rect 73 34 95 35
rect 105 37 127 38
rect 105 35 110 37
rect 112 35 117 37
rect 119 35 127 37
rect 105 34 127 35
rect 13 28 58 30
rect 13 26 54 28
rect 56 26 58 28
rect 13 25 17 26
rect 13 23 14 25
rect 16 23 17 25
rect 13 21 17 23
rect 33 25 58 26
rect 33 23 34 25
rect 36 23 38 25
rect 33 17 38 23
rect -2 1 146 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 146 1
rect -2 -2 146 -1
<< ptie >>
rect 0 1 144 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 144 1
rect 0 -3 144 -1
<< ntie >>
rect 0 81 144 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 144 81
rect 0 77 144 79
<< nmos >>
rect 19 16 21 27
rect 29 16 31 27
rect 39 12 41 30
rect 49 12 51 30
rect 59 12 61 30
rect 69 12 71 30
rect 79 12 81 30
rect 89 12 91 30
rect 99 12 101 30
rect 109 12 111 30
rect 119 12 121 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 42 81 70
rect 89 42 91 70
rect 99 42 101 70
rect 109 42 111 70
rect 119 42 121 70
<< polyct1 >>
rect 11 35 13 37
rect 45 35 47 37
rect 57 35 59 37
rect 77 35 79 37
rect 85 35 87 37
rect 110 35 112 37
rect 117 35 119 37
<< ndifct0 >>
rect 24 18 26 20
rect 44 18 46 20
rect 64 25 66 27
rect 64 18 66 20
rect 74 26 76 28
rect 84 18 86 20
rect 94 26 96 28
rect 94 19 96 21
rect 104 14 106 16
rect 114 26 116 28
rect 114 19 116 21
rect 124 22 126 24
rect 124 14 126 16
<< ndifct1 >>
rect 14 23 16 25
rect 34 23 36 25
rect 54 26 56 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
<< pdifct0 >>
rect 14 59 16 61
rect 14 52 16 54
rect 24 51 26 53
rect 34 59 36 61
rect 34 52 36 54
rect 44 66 46 68
rect 44 59 46 61
rect 54 51 56 53
rect 54 44 56 46
rect 64 66 66 68
rect 64 59 66 61
rect 74 51 76 53
rect 74 44 76 46
rect 84 66 86 68
rect 84 59 86 61
rect 94 51 96 53
rect 94 44 96 46
rect 104 66 106 68
rect 104 59 106 61
rect 114 59 116 61
rect 114 52 116 54
rect 124 66 126 68
rect 124 59 126 61
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 44 26 46
<< alu0 >>
rect 42 66 44 68
rect 46 66 48 68
rect 12 61 38 62
rect 12 59 14 61
rect 16 59 34 61
rect 36 59 38 61
rect 12 58 38 59
rect 42 61 48 66
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 62 66 64 68
rect 66 66 68 68
rect 62 61 68 66
rect 62 59 64 61
rect 66 59 68 61
rect 62 58 68 59
rect 82 66 84 68
rect 86 66 88 68
rect 82 61 88 66
rect 82 59 84 61
rect 86 59 88 61
rect 82 58 88 59
rect 102 66 104 68
rect 106 66 108 68
rect 102 61 108 66
rect 122 66 124 68
rect 126 66 128 68
rect 102 59 104 61
rect 106 59 108 61
rect 102 58 108 59
rect 113 61 117 63
rect 113 59 114 61
rect 116 59 117 61
rect 12 54 18 58
rect 32 54 38 58
rect 113 54 117 59
rect 122 61 128 66
rect 122 59 124 61
rect 126 59 128 61
rect 122 58 128 59
rect 12 52 14 54
rect 16 52 18 54
rect 12 51 18 52
rect 22 53 28 54
rect 22 51 24 53
rect 26 51 28 53
rect 22 46 28 51
rect 32 52 34 54
rect 36 53 114 54
rect 36 52 54 53
rect 32 51 54 52
rect 56 51 74 53
rect 76 51 94 53
rect 96 52 114 53
rect 116 52 117 54
rect 96 51 117 52
rect 32 50 117 51
rect 53 46 57 50
rect 53 44 54 46
rect 56 44 57 46
rect 53 42 57 44
rect 73 46 77 50
rect 93 46 97 50
rect 73 44 74 46
rect 76 44 77 46
rect 73 42 77 44
rect 93 44 94 46
rect 96 44 97 46
rect 93 42 97 44
rect 63 27 67 29
rect 63 25 64 27
rect 66 25 67 27
rect 72 28 118 29
rect 72 26 74 28
rect 76 26 94 28
rect 96 26 114 28
rect 116 26 118 28
rect 72 25 118 26
rect 23 20 27 22
rect 23 18 24 20
rect 26 18 27 20
rect 23 12 27 18
rect 63 21 67 25
rect 93 21 97 25
rect 42 20 88 21
rect 42 18 44 20
rect 46 18 64 20
rect 66 18 84 20
rect 86 18 88 20
rect 42 17 88 18
rect 93 19 94 21
rect 96 19 97 21
rect 93 17 97 19
rect 113 21 118 25
rect 113 19 114 21
rect 116 19 118 21
rect 103 16 107 18
rect 113 17 118 19
rect 123 24 127 26
rect 123 22 124 24
rect 126 22 127 24
rect 103 14 104 16
rect 106 14 107 16
rect 103 12 107 14
rect 123 16 127 22
rect 123 14 124 16
rect 126 14 127 16
rect 123 12 127 14
<< labels >>
rlabel alu0 15 56 15 56 6 n3
rlabel alu0 55 48 55 48 6 n3
rlabel alu0 35 56 35 56 6 n3
rlabel alu0 65 23 65 23 6 n2
rlabel alu0 75 48 75 48 6 n3
rlabel ndifct0 65 19 65 19 6 n2
rlabel alu0 95 23 95 23 6 n1
rlabel alu0 95 48 95 48 6 n3
rlabel alu0 115 23 115 23 6 n1
rlabel ndifct0 95 27 95 27 6 n1
rlabel alu0 115 56 115 56 6 n3
rlabel alu0 74 52 74 52 6 n3
rlabel alu1 28 32 28 32 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 24 4 24 6 b
rlabel alu1 20 28 20 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 4 56 4 56 6 z
rlabel alu1 36 24 36 24 6 z
rlabel alu1 60 36 60 36 6 a3
rlabel alu1 52 36 52 36 6 a3
rlabel alu1 52 28 52 28 6 z
rlabel alu1 44 28 44 28 6 z
rlabel alu1 44 40 44 40 6 a3
rlabel alu1 72 6 72 6 6 vss
rlabel alu1 76 36 76 36 6 a2
rlabel alu1 92 36 92 36 6 a2
rlabel alu1 84 40 84 40 6 a2
rlabel alu1 72 74 72 74 6 vdd
rlabel alu1 108 36 108 36 6 a1
rlabel alu1 116 36 116 36 6 a1
rlabel alu1 124 44 124 44 6 a1
<< end >>
