magic
tech scmos
timestamp 1199201859
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 41 61 43 65
rect 9 33 11 50
rect 19 47 21 50
rect 29 47 31 50
rect 16 45 22 47
rect 16 43 18 45
rect 20 43 22 45
rect 16 41 22 43
rect 26 45 32 47
rect 26 43 28 45
rect 30 43 32 45
rect 26 41 32 43
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 9 27 15 29
rect 13 24 15 27
rect 20 24 22 41
rect 30 24 32 41
rect 41 39 43 45
rect 37 37 43 39
rect 37 35 39 37
rect 41 35 43 37
rect 37 33 43 35
rect 37 24 39 33
rect 13 12 15 17
rect 20 12 22 17
rect 30 12 32 17
rect 37 12 39 17
<< ndif >>
rect 4 17 13 24
rect 15 17 20 24
rect 22 21 30 24
rect 22 19 25 21
rect 27 19 30 21
rect 22 17 30 19
rect 32 17 37 24
rect 39 21 48 24
rect 39 19 43 21
rect 45 19 48 21
rect 39 17 48 19
rect 4 11 11 17
rect 4 9 7 11
rect 9 9 11 11
rect 4 7 11 9
<< pdif >>
rect 33 71 39 73
rect 33 69 35 71
rect 37 69 39 71
rect 33 66 39 69
rect 4 64 9 66
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 50 9 58
rect 11 54 19 66
rect 11 52 14 54
rect 16 52 19 54
rect 11 50 19 52
rect 21 62 29 66
rect 21 60 24 62
rect 26 60 29 62
rect 21 55 29 60
rect 21 53 24 55
rect 26 53 29 55
rect 21 50 29 53
rect 31 61 39 66
rect 31 50 41 61
rect 34 45 41 50
rect 43 59 50 61
rect 43 57 46 59
rect 48 57 50 59
rect 43 52 50 57
rect 43 50 46 52
rect 48 50 50 52
rect 43 48 50 50
rect 43 45 48 48
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 35 71
rect 37 69 58 71
rect -2 68 58 69
rect 2 54 18 55
rect 2 52 14 54
rect 16 52 18 54
rect 2 51 18 52
rect 2 22 6 51
rect 10 45 21 47
rect 34 46 38 55
rect 10 43 18 45
rect 20 43 21 45
rect 10 41 21 43
rect 25 45 47 46
rect 25 43 28 45
rect 30 43 47 45
rect 25 42 47 43
rect 17 38 21 41
rect 17 34 23 38
rect 27 37 47 38
rect 27 35 39 37
rect 41 35 47 37
rect 27 34 47 35
rect 10 29 11 30
rect 13 29 38 30
rect 10 26 38 29
rect 2 21 29 22
rect 2 19 25 21
rect 27 19 29 21
rect 2 17 29 19
rect 34 17 38 26
rect 42 25 47 34
rect -2 11 58 12
rect -2 9 7 11
rect 9 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 13 17 15 24
rect 20 17 22 24
rect 30 17 32 24
rect 37 17 39 24
<< pmos >>
rect 9 50 11 66
rect 19 50 21 66
rect 29 50 31 66
rect 41 45 43 61
<< polyct0 >>
rect 11 30 13 31
<< polyct1 >>
rect 18 43 20 45
rect 28 43 30 45
rect 11 29 13 30
rect 39 35 41 37
<< ndifct0 >>
rect 43 19 45 21
<< ndifct1 >>
rect 25 19 27 21
rect 7 9 9 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 60 6 62
rect 24 60 26 62
rect 24 53 26 55
rect 46 57 48 59
rect 46 50 48 52
<< pdifct1 >>
rect 35 69 37 71
rect 14 52 16 54
<< alu0 >>
rect 2 62 50 63
rect 2 60 4 62
rect 6 60 24 62
rect 26 60 50 62
rect 2 59 50 60
rect 23 55 27 59
rect 44 57 46 59
rect 48 57 50 59
rect 23 53 24 55
rect 26 53 27 55
rect 23 51 27 53
rect 44 52 50 57
rect 44 50 46 52
rect 48 50 50 52
rect 44 49 50 50
rect 10 31 14 33
rect 10 30 11 31
rect 13 30 14 31
rect 41 21 47 22
rect 41 19 43 21
rect 45 19 47 21
rect 41 12 47 19
<< labels >>
rlabel alu0 25 57 25 57 6 n3
rlabel alu0 47 56 47 56 6 n3
rlabel alu0 26 61 26 61 6 n3
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 28 20 28 6 b1
rlabel alu1 20 36 20 36 6 b2
rlabel alu1 12 44 12 44 6 b2
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 20 36 20 6 b1
rlabel alu1 28 28 28 28 6 b1
rlabel alu1 36 36 36 36 6 a1
rlabel alu1 28 44 28 44 6 a2
rlabel alu1 36 48 36 48 6 a2
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 44 44 44 44 6 a2
<< end >>
