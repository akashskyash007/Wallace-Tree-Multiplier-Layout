magic
tech scmos
timestamp 1684146972
<< ab >>
rect -35 6 45 77
rect 48 6 88 77
rect -44 5 88 6
rect -44 -66 52 5
<< nwell >>
rect -40 37 93 82
rect -49 -71 57 -26
<< pwell >>
rect -40 11 93 37
rect -49 0 93 11
rect -49 -26 57 0
<< poly >>
rect -26 62 -24 66
rect -16 64 -14 69
rect -6 64 -4 69
rect 14 62 16 66
rect 24 64 26 69
rect 34 64 36 69
rect -26 40 -24 44
rect -16 40 -14 51
rect -6 48 -4 51
rect -6 46 0 48
rect -6 44 -4 46
rect -2 44 0 46
rect 57 62 59 66
rect 67 64 69 69
rect 77 64 79 69
rect -6 42 0 44
rect -26 38 -20 40
rect -26 36 -24 38
rect -22 36 -20 38
rect -26 34 -20 36
rect -16 38 -10 40
rect -16 36 -14 38
rect -12 36 -10 38
rect -16 34 -10 36
rect -26 29 -24 34
rect -13 29 -11 34
rect -6 29 -4 42
rect 14 40 16 44
rect 24 40 26 51
rect 34 48 36 51
rect 34 46 40 48
rect 34 44 36 46
rect 38 44 40 46
rect 34 42 40 44
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 29 16 34
rect 27 29 29 34
rect 34 29 36 42
rect 57 40 59 44
rect 67 40 69 51
rect 77 48 79 51
rect 77 46 83 48
rect 77 44 79 46
rect 81 44 83 46
rect 77 42 83 44
rect 57 38 63 40
rect 57 36 59 38
rect 61 36 63 38
rect 57 34 63 36
rect 67 38 73 40
rect 67 36 69 38
rect 71 36 73 38
rect 67 34 73 36
rect 57 29 59 34
rect 70 29 72 34
rect 77 29 79 42
rect -26 16 -24 20
rect -13 13 -11 18
rect -6 13 -4 18
rect 14 16 16 20
rect 27 13 29 18
rect 34 13 36 18
rect 57 16 59 20
rect 70 13 72 18
rect 77 13 79 18
rect -27 0 -25 4
rect -16 0 -14 4
rect -9 0 -7 4
rect -27 -23 -25 -14
rect 11 -6 13 -1
rect 21 -6 23 -1
rect 31 -3 33 2
rect 41 0 43 4
rect -16 -23 -14 -20
rect -9 -23 -7 -20
rect 11 -23 13 -20
rect 21 -23 23 -20
rect -29 -25 -23 -23
rect -29 -27 -27 -25
rect -25 -27 -23 -25
rect -29 -29 -23 -27
rect -19 -25 -13 -23
rect -19 -27 -17 -25
rect -15 -27 -13 -25
rect -19 -29 -13 -27
rect -9 -25 13 -23
rect -9 -27 -7 -25
rect -5 -27 0 -25
rect 2 -27 13 -25
rect -9 -29 13 -27
rect 17 -25 23 -23
rect 17 -27 19 -25
rect 21 -27 23 -25
rect 17 -29 23 -27
rect 31 -26 33 -13
rect 41 -16 43 -13
rect 37 -18 43 -16
rect 37 -20 39 -18
rect 41 -20 43 -18
rect 37 -22 43 -20
rect 31 -28 37 -26
rect -27 -32 -25 -29
rect -17 -32 -15 -29
rect -7 -32 -5 -29
rect 11 -32 13 -29
rect 18 -32 20 -29
rect 31 -30 33 -28
rect 35 -30 37 -28
rect 28 -32 37 -30
rect 28 -35 30 -32
rect 41 -35 43 -22
rect 28 -53 30 -48
rect -27 -64 -25 -60
rect -17 -64 -15 -60
rect -7 -64 -5 -60
rect 11 -62 13 -57
rect 18 -62 20 -57
rect 41 -64 43 -60
<< ndif >>
rect -31 26 -26 29
rect -33 24 -26 26
rect -33 22 -31 24
rect -29 22 -26 24
rect -33 20 -26 22
rect -24 20 -13 29
rect -22 18 -13 20
rect -11 18 -6 29
rect -4 24 1 29
rect 9 26 14 29
rect 7 24 14 26
rect -4 22 3 24
rect -4 20 -1 22
rect 1 20 3 22
rect 7 22 9 24
rect 11 22 14 24
rect 7 20 14 22
rect 16 20 27 29
rect -4 18 3 20
rect -22 12 -15 18
rect 18 18 27 20
rect 29 18 34 29
rect 36 24 41 29
rect 52 26 57 29
rect 50 24 57 26
rect 36 22 43 24
rect 36 20 39 22
rect 41 20 43 22
rect 50 22 52 24
rect 54 22 57 24
rect 50 20 57 22
rect 59 20 70 29
rect 36 18 43 20
rect -22 10 -20 12
rect -18 10 -15 12
rect -22 8 -15 10
rect 18 12 25 18
rect 61 18 70 20
rect 72 18 77 29
rect 79 24 84 29
rect 79 22 86 24
rect 79 20 82 22
rect 84 20 86 22
rect 79 18 86 20
rect 18 10 20 12
rect 22 10 25 12
rect 18 8 25 10
rect 61 12 68 18
rect 61 10 63 12
rect 65 10 68 12
rect 61 8 68 10
rect -32 -7 -27 0
rect -34 -9 -27 -7
rect -34 -11 -32 -9
rect -30 -11 -27 -9
rect -34 -14 -27 -11
rect -25 -2 -16 0
rect -25 -4 -21 -2
rect -19 -4 -16 -2
rect -25 -14 -16 -4
rect -23 -20 -16 -14
rect -14 -20 -9 0
rect -7 -7 -2 0
rect 36 -3 41 0
rect 26 -6 31 -3
rect -7 -9 0 -7
rect -7 -11 -4 -9
rect -2 -11 0 -9
rect -7 -13 0 -11
rect 4 -9 11 -6
rect 4 -11 6 -9
rect 8 -11 11 -9
rect -7 -20 -2 -13
rect 4 -16 11 -11
rect 4 -18 6 -16
rect 8 -18 11 -16
rect 4 -20 11 -18
rect 13 -16 21 -6
rect 13 -18 16 -16
rect 18 -18 21 -16
rect 13 -20 21 -18
rect 23 -8 31 -6
rect 23 -10 26 -8
rect 28 -10 31 -8
rect 23 -13 31 -10
rect 33 -5 41 -3
rect 33 -7 36 -5
rect 38 -7 41 -5
rect 33 -13 41 -7
rect 43 -7 48 0
rect 43 -9 50 -7
rect 43 -11 46 -9
rect 48 -11 50 -9
rect 43 -13 50 -11
rect 23 -20 28 -13
<< pdif >>
rect -22 62 -16 64
rect -31 57 -26 62
rect -33 55 -26 57
rect -33 53 -31 55
rect -29 53 -26 55
rect -33 48 -26 53
rect -33 46 -31 48
rect -29 46 -26 48
rect -33 44 -26 46
rect -24 60 -16 62
rect -24 58 -21 60
rect -19 58 -16 60
rect -24 51 -16 58
rect -14 62 -6 64
rect -14 60 -11 62
rect -9 60 -6 62
rect -14 55 -6 60
rect -14 53 -11 55
rect -9 53 -6 55
rect -14 51 -6 53
rect -4 62 3 64
rect 18 62 24 64
rect -4 60 -1 62
rect 1 60 3 62
rect -4 51 3 60
rect 9 57 14 62
rect 7 55 14 57
rect 7 53 9 55
rect 11 53 14 55
rect -24 44 -18 51
rect 7 48 14 53
rect 7 46 9 48
rect 11 46 14 48
rect 7 44 14 46
rect 16 60 24 62
rect 16 58 19 60
rect 21 58 24 60
rect 16 51 24 58
rect 26 62 34 64
rect 26 60 29 62
rect 31 60 34 62
rect 26 55 34 60
rect 26 53 29 55
rect 31 53 34 55
rect 26 51 34 53
rect 36 62 43 64
rect 61 62 67 64
rect 36 60 39 62
rect 41 60 43 62
rect 36 51 43 60
rect 52 57 57 62
rect 50 55 57 57
rect 50 53 52 55
rect 54 53 57 55
rect 16 44 22 51
rect 50 48 57 53
rect 50 46 52 48
rect 54 46 57 48
rect 50 44 57 46
rect 59 60 67 62
rect 59 58 62 60
rect 64 58 67 60
rect 59 51 67 58
rect 69 62 77 64
rect 69 60 72 62
rect 74 60 77 62
rect 69 55 77 60
rect 69 53 72 55
rect 74 53 77 55
rect 69 51 77 53
rect 79 62 86 64
rect 79 60 82 62
rect 84 60 86 62
rect 79 51 86 60
rect 59 44 65 51
rect -34 -34 -27 -32
rect -34 -36 -32 -34
rect -30 -36 -27 -34
rect -34 -41 -27 -36
rect -34 -43 -32 -41
rect -30 -43 -27 -41
rect -34 -45 -27 -43
rect -32 -60 -27 -45
rect -25 -49 -17 -32
rect -25 -51 -22 -49
rect -20 -51 -17 -49
rect -25 -56 -17 -51
rect -25 -58 -22 -56
rect -20 -58 -17 -56
rect -25 -60 -17 -58
rect -15 -41 -7 -32
rect -15 -43 -12 -41
rect -10 -43 -7 -41
rect -15 -48 -7 -43
rect -15 -50 -12 -48
rect -10 -50 -7 -48
rect -15 -60 -7 -50
rect -5 -49 11 -32
rect -5 -51 0 -49
rect 2 -51 11 -49
rect -5 -56 11 -51
rect -5 -58 0 -56
rect 2 -57 11 -56
rect 13 -57 18 -32
rect 20 -35 25 -32
rect 20 -37 28 -35
rect 20 -39 23 -37
rect 25 -39 28 -37
rect 20 -48 28 -39
rect 30 -48 41 -35
rect 20 -57 25 -48
rect 32 -56 41 -48
rect 2 -58 9 -57
rect -5 -60 9 -58
rect 32 -58 35 -56
rect 37 -58 41 -56
rect 32 -60 41 -58
rect 43 -37 50 -35
rect 43 -39 46 -37
rect 48 -39 50 -37
rect 43 -44 50 -39
rect 43 -46 46 -44
rect 48 -46 50 -44
rect 43 -48 50 -46
rect 43 -60 48 -48
<< alu1 >>
rect -37 72 90 77
rect -37 70 -30 72
rect -28 70 10 72
rect 12 70 53 72
rect 55 70 90 72
rect -37 69 90 70
rect -33 55 -28 57
rect -33 53 -31 55
rect -29 53 -28 55
rect -33 48 -28 53
rect -33 46 -31 48
rect -29 46 -28 48
rect -33 44 -28 46
rect -1 55 3 56
rect -1 53 0 55
rect 2 53 3 55
rect -33 24 -29 44
rect -1 47 3 53
rect -10 46 3 47
rect -10 44 -4 46
rect -2 44 3 46
rect -10 43 3 44
rect 7 55 12 57
rect 7 53 9 55
rect 11 53 12 55
rect 7 48 12 53
rect 7 46 9 48
rect 11 46 12 48
rect 7 44 12 46
rect -18 38 -4 39
rect -18 36 -14 38
rect -12 36 -4 38
rect -18 35 -4 36
rect -33 22 -31 24
rect -29 22 -21 24
rect -33 21 -21 22
rect -33 19 -25 21
rect -23 19 -21 21
rect -9 26 -4 35
rect 7 24 11 44
rect 39 47 43 56
rect 30 46 43 47
rect 30 44 36 46
rect 38 44 43 46
rect 30 43 43 44
rect 50 55 55 57
rect 50 53 52 55
rect 54 53 55 55
rect 50 48 55 53
rect 50 46 52 48
rect 54 46 55 48
rect 50 44 55 46
rect 82 55 86 56
rect 82 53 83 55
rect 85 53 86 55
rect 22 38 36 39
rect 22 36 26 38
rect 28 36 36 38
rect 22 35 36 36
rect 7 22 9 24
rect 11 22 19 24
rect 7 21 19 22
rect 7 19 15 21
rect 17 19 19 21
rect 31 29 36 35
rect 31 27 33 29
rect 35 27 36 29
rect 31 26 36 27
rect 50 24 54 44
rect 82 47 86 53
rect 73 46 86 47
rect 73 44 79 46
rect 81 44 86 46
rect 73 43 86 44
rect 65 38 79 39
rect 65 36 69 38
rect 71 36 79 38
rect 65 35 79 36
rect 50 22 52 24
rect 54 22 62 24
rect -33 18 -21 19
rect 7 18 19 19
rect 50 18 62 22
rect 74 29 79 35
rect 74 27 76 29
rect 78 27 79 29
rect 74 26 79 27
rect -37 12 90 13
rect -37 10 -30 12
rect -28 10 -20 12
rect -18 10 10 12
rect 12 10 20 12
rect 22 10 53 12
rect 55 10 63 12
rect 65 10 90 12
rect -37 6 90 10
rect -46 5 90 6
rect -46 -2 54 5
rect -35 -9 -13 -8
rect -35 -11 -32 -9
rect -30 -11 -13 -9
rect -35 -12 -13 -11
rect 45 -9 50 -7
rect 45 -11 46 -9
rect 48 -11 50 -9
rect -35 -32 -31 -12
rect -2 -17 2 -15
rect -2 -19 -1 -17
rect 1 -19 2 -17
rect -35 -34 -29 -32
rect -35 -36 -32 -34
rect -30 -36 -29 -34
rect -35 -41 -29 -36
rect -35 -43 -32 -41
rect -30 -43 -29 -41
rect -35 -45 -29 -43
rect -2 -24 2 -19
rect 45 -13 50 -11
rect 14 -24 22 -23
rect -11 -25 4 -24
rect -11 -27 -7 -25
rect -5 -27 0 -25
rect 2 -27 4 -25
rect -11 -28 4 -27
rect 14 -26 15 -24
rect 17 -25 22 -24
rect 17 -26 19 -25
rect 14 -27 19 -26
rect 21 -27 22 -25
rect 14 -29 22 -27
rect 14 -32 19 -29
rect -19 -36 19 -32
rect 46 -35 50 -13
rect 45 -37 50 -35
rect 45 -39 46 -37
rect 48 -39 50 -37
rect 45 -44 50 -39
rect 45 -46 46 -44
rect 48 -46 50 -44
rect 45 -48 50 -46
rect 37 -52 50 -48
rect -46 -66 54 -58
<< alu2 >>
rect -1 60 3 61
rect -1 58 0 60
rect 2 58 3 60
rect -1 55 3 58
rect -1 53 0 55
rect 2 53 3 55
rect -1 52 3 53
rect 82 60 86 61
rect 82 58 83 60
rect 85 58 86 60
rect 82 55 86 58
rect 82 53 83 55
rect 85 53 86 55
rect 82 52 86 53
rect 32 29 36 31
rect 32 27 33 29
rect 35 27 36 29
rect 32 26 36 27
rect 32 24 33 26
rect 35 24 36 26
rect -26 21 -21 24
rect 32 23 36 24
rect 75 29 79 31
rect 75 27 76 29
rect 78 27 79 29
rect 75 26 79 27
rect 75 24 76 26
rect 78 24 79 26
rect 75 23 79 24
rect -26 19 -25 21
rect -23 19 -21 21
rect -26 -9 -21 19
rect 14 21 19 22
rect 14 19 15 21
rect 17 19 19 21
rect -26 -11 -25 -9
rect -23 -11 -21 -9
rect -26 -12 -21 -11
rect -2 -9 2 -8
rect -2 -11 -1 -9
rect 1 -11 2 -9
rect -2 -17 2 -11
rect -2 -19 -1 -17
rect 1 -19 2 -17
rect -2 -20 2 -19
rect 14 -24 19 19
rect 14 -26 15 -24
rect 17 -26 19 -24
rect 14 -27 19 -26
<< alu3 >>
rect -1 60 86 61
rect -1 58 0 60
rect 2 58 83 60
rect 85 58 86 60
rect -1 56 86 58
rect 32 26 79 27
rect 32 24 33 26
rect 35 24 76 26
rect 78 24 79 26
rect 32 23 79 24
rect -26 -9 2 -8
rect -26 -11 -25 -9
rect -23 -11 -1 -9
rect 1 -11 2 -9
rect -26 -12 2 -11
<< ptie >>
rect -32 12 -26 14
rect -32 10 -30 12
rect -28 10 -26 12
rect -32 8 -26 10
rect 8 12 14 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 51 12 57 14
rect 51 10 53 12
rect 55 10 57 12
rect 51 8 57 10
<< ntie >>
rect -32 72 -26 74
rect -32 70 -30 72
rect -28 70 -26 72
rect -32 68 -26 70
rect 8 72 14 74
rect 8 70 10 72
rect 12 70 14 72
rect 8 68 14 70
rect 51 72 57 74
rect 51 70 53 72
rect 55 70 57 72
rect 51 68 57 70
<< nmos >>
rect -26 20 -24 29
rect -13 18 -11 29
rect -6 18 -4 29
rect 14 20 16 29
rect 27 18 29 29
rect 34 18 36 29
rect 57 20 59 29
rect 70 18 72 29
rect 77 18 79 29
rect -27 -14 -25 0
rect -16 -20 -14 0
rect -9 -20 -7 0
rect 11 -20 13 -6
rect 21 -20 23 -6
rect 31 -13 33 -3
rect 41 -13 43 0
<< pmos >>
rect -26 44 -24 62
rect -16 51 -14 64
rect -6 51 -4 64
rect 14 44 16 62
rect 24 51 26 64
rect 34 51 36 64
rect 57 44 59 62
rect 67 51 69 64
rect 77 51 79 64
rect -27 -60 -25 -32
rect -17 -60 -15 -32
rect -7 -60 -5 -32
rect 11 -57 13 -32
rect 18 -57 20 -32
rect 28 -48 30 -35
rect 41 -60 43 -35
<< polyct0 >>
rect -24 36 -22 38
rect 16 36 18 38
rect 59 36 61 38
rect -27 -27 -25 -25
rect -17 -27 -15 -25
rect 39 -20 41 -18
rect 33 -30 35 -28
<< polyct1 >>
rect -4 44 -2 46
rect -14 36 -12 38
rect 36 44 38 46
rect 26 36 28 38
rect 79 44 81 46
rect 69 36 71 38
rect -7 -27 -5 -25
rect 0 -27 2 -25
rect 19 -27 21 -25
<< ndifct0 >>
rect -1 20 1 22
rect 39 20 41 22
rect 82 20 84 22
rect -21 -4 -19 -2
rect -4 -11 -2 -9
rect 6 -11 8 -9
rect 6 -18 8 -16
rect 16 -18 18 -16
rect 26 -10 28 -8
rect 36 -7 38 -5
<< ndifct1 >>
rect -31 22 -29 24
rect 9 22 11 24
rect 52 22 54 24
rect -20 10 -18 12
rect 20 10 22 12
rect 63 10 65 12
rect -32 -11 -30 -9
rect 46 -11 48 -9
<< ntiect1 >>
rect -30 70 -28 72
rect 10 70 12 72
rect 53 70 55 72
<< ptiect1 >>
rect -30 10 -28 12
rect 10 10 12 12
rect 53 10 55 12
<< pdifct0 >>
rect -21 58 -19 60
rect -11 60 -9 62
rect -11 53 -9 55
rect -1 60 1 62
rect 19 58 21 60
rect 29 60 31 62
rect 29 53 31 55
rect 39 60 41 62
rect 62 58 64 60
rect 72 60 74 62
rect 72 53 74 55
rect 82 60 84 62
rect -22 -51 -20 -49
rect -22 -58 -20 -56
rect -12 -43 -10 -41
rect -12 -50 -10 -48
rect 0 -51 2 -49
rect 0 -58 2 -56
rect 23 -39 25 -37
rect 35 -58 37 -56
<< pdifct1 >>
rect -31 53 -29 55
rect -31 46 -29 48
rect 9 53 11 55
rect 9 46 11 48
rect 52 53 54 55
rect 52 46 54 48
rect -32 -36 -30 -34
rect -32 -43 -30 -41
rect 46 -39 48 -37
rect 46 -46 48 -44
<< alu0 >>
rect -23 60 -17 69
rect -23 58 -21 60
rect -19 58 -17 60
rect -23 57 -17 58
rect -12 62 -8 64
rect -12 60 -11 62
rect -9 60 -8 62
rect -12 55 -8 60
rect -3 62 3 69
rect -3 60 -1 62
rect 1 60 3 62
rect -3 59 3 60
rect 17 60 23 69
rect 17 58 19 60
rect 21 58 23 60
rect 17 57 23 58
rect 28 62 32 64
rect 28 60 29 62
rect 31 60 32 62
rect -12 54 -11 55
rect -25 53 -11 54
rect -9 53 -8 55
rect -25 50 -8 53
rect -25 38 -21 50
rect 28 55 32 60
rect 37 62 43 69
rect 37 60 39 62
rect 41 60 43 62
rect 37 59 43 60
rect 60 60 66 69
rect 60 58 62 60
rect 64 58 66 60
rect 60 57 66 58
rect 71 62 75 64
rect 71 60 72 62
rect 74 60 75 62
rect 28 54 29 55
rect 15 53 29 54
rect 31 53 32 55
rect 15 50 32 53
rect -25 36 -24 38
rect -22 36 -21 38
rect -25 31 -21 36
rect -25 27 -13 31
rect -29 24 -28 26
rect -17 23 -13 27
rect 15 38 19 50
rect 71 55 75 60
rect 80 62 86 69
rect 80 60 82 62
rect 84 60 86 62
rect 80 59 86 60
rect 71 54 72 55
rect 58 53 72 54
rect 74 53 75 55
rect 58 50 75 53
rect 15 36 16 38
rect 18 36 19 38
rect 15 31 19 36
rect 15 27 27 31
rect 11 24 12 26
rect -17 22 3 23
rect -17 20 -1 22
rect 1 20 3 22
rect -17 19 3 20
rect 23 23 27 27
rect 58 38 62 50
rect 58 36 59 38
rect 61 36 62 38
rect 58 31 62 36
rect 58 27 70 31
rect 54 24 55 26
rect 23 22 43 23
rect 23 20 39 22
rect 41 20 43 22
rect 23 19 43 20
rect 66 23 70 27
rect 66 22 86 23
rect 66 20 82 22
rect 84 20 86 22
rect 66 19 86 20
rect -23 -4 -21 -2
rect -19 -4 -17 -2
rect -23 -5 -17 -4
rect 35 -5 39 -2
rect 35 -7 36 -5
rect 38 -7 39 -5
rect 5 -8 30 -7
rect -10 -9 0 -8
rect -10 -11 -4 -9
rect -2 -11 0 -9
rect -10 -12 0 -11
rect 5 -9 26 -8
rect 5 -11 6 -9
rect 8 -10 26 -9
rect 28 -10 30 -8
rect 35 -9 39 -7
rect 8 -11 30 -10
rect -10 -16 -6 -12
rect -26 -20 -6 -16
rect -26 -23 -22 -20
rect -28 -25 -22 -23
rect -28 -27 -27 -25
rect -25 -27 -22 -25
rect -28 -29 -22 -27
rect -26 -40 -22 -29
rect -18 -25 -14 -23
rect 5 -16 9 -11
rect 5 -18 6 -16
rect 8 -18 9 -16
rect 5 -20 9 -18
rect 14 -16 29 -15
rect 14 -18 16 -16
rect 18 -17 29 -16
rect 18 -18 43 -17
rect 14 -19 39 -18
rect 25 -20 39 -19
rect 41 -20 43 -18
rect 25 -21 43 -20
rect -18 -27 -17 -25
rect -15 -27 -14 -25
rect -18 -32 -14 -27
rect 25 -32 29 -21
rect 22 -36 29 -32
rect 32 -28 36 -26
rect 32 -30 33 -28
rect 35 -30 36 -28
rect 22 -37 26 -36
rect 22 -39 23 -37
rect 25 -39 26 -37
rect -26 -41 14 -40
rect 22 -41 26 -39
rect 32 -40 36 -30
rect -26 -43 -12 -41
rect -10 -43 14 -41
rect -26 -44 14 -43
rect 30 -44 36 -40
rect -13 -48 -9 -44
rect 10 -48 34 -44
rect -24 -49 -18 -48
rect -24 -51 -22 -49
rect -20 -51 -18 -49
rect -24 -56 -18 -51
rect -13 -50 -12 -48
rect -10 -50 -9 -48
rect -13 -52 -9 -50
rect -2 -49 4 -48
rect -2 -51 0 -49
rect 2 -51 4 -49
rect -24 -58 -22 -56
rect -20 -58 -18 -56
rect -2 -56 4 -51
rect -2 -58 0 -56
rect 2 -58 4 -56
rect 33 -56 39 -55
rect 33 -58 35 -56
rect 37 -58 39 -56
<< via1 >>
rect 0 53 2 55
rect -25 19 -23 21
rect 83 53 85 55
rect 15 19 17 21
rect 33 27 35 29
rect 76 27 78 29
rect -1 -19 1 -17
rect 15 -26 17 -24
<< via2 >>
rect 0 58 2 60
rect 83 58 85 60
rect 33 24 35 26
rect 76 24 78 26
rect -25 -11 -23 -9
rect -1 -11 1 -9
<< labels >>
rlabel alu1 25 9 25 9 6 vss
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 25 37 25 37 1 a0
rlabel alu1 33 33 33 33 1 a0
rlabel alu1 33 45 33 45 1 b1
rlabel alu1 41 53 41 53 1 b1
rlabel alu1 9 37 9 37 1 a0b1
rlabel alu1 17 21 17 21 1 a0b1
rlabel alu0 17 40 17 40 1 a0b1_inv
rlabel alu0 30 57 30 57 1 a0b1_inv
rlabel alu1 -15 9 -15 9 6 vss
rlabel alu1 -15 73 -15 73 6 vdd
rlabel alu1 -15 37 -15 37 1 a1
rlabel alu1 -7 33 -7 33 1 a1
rlabel alu1 -7 45 -7 45 1 b0
rlabel alu1 -31 37 -31 37 1 a1b0
rlabel alu1 -23 21 -23 21 1 a1b0
rlabel alu0 33 21 33 21 1 a0b1inv
rlabel alu0 -10 57 -10 57 1 a1b0inv
rlabel alu0 -23 40 -23 40 1 a1b0inv
rlabel alu0 -7 21 -7 21 1 a1b0inv
rlabel alu1 4 -62 4 -62 2 vdd
rlabel alu1 4 2 4 2 2 vss
rlabel ndifct1 -32 -10 -32 -10 1 c01
rlabel alu1 -24 -10 -24 -10 1 c01
rlabel alu1 -16 -10 -16 -10 1 c01
rlabel alu1 -32 -38 -32 -38 1 c01
rlabel alu0 -5 -10 -5 -10 1 c01_inv
rlabel alu0 -24 -30 -24 -30 1 c01_inv
rlabel alu0 -11 -46 -11 -46 1 c01_inv
rlabel alu0 -6 -42 -6 -42 1 c01_inv
rlabel alu1 48 -26 48 -26 1 res1
rlabel alu1 40 -50 40 -50 1 res1
rlabel alu0 34 -35 34 -35 1 c01_inv
rlabel alu0 34 -19 34 -19 1 res1_inv
rlabel alu0 24 -36 24 -36 1 res1_inv
rlabel alu0 22 -17 22 -17 1 res1_inv
rlabel alu0 7 -13 7 -13 1 ha01
rlabel alu0 18 -9 18 -9 1 ha01
rlabel alu1 0 -22 0 -22 1 a1b0
rlabel alu1 -8 -26 -8 -26 1 a1b0
rlabel alu1 -16 -34 -16 -34 1 a0b1
rlabel alu1 -8 -34 -8 -34 1 a0b1
rlabel alu1 0 -34 0 -34 1 a0b1
rlabel alu1 8 -34 8 -34 1 a0b1
rlabel alu1 16 -30 16 -30 1 a0b1
rlabel alu1 68 9 68 9 6 vss
rlabel alu1 68 73 68 73 6 vdd
rlabel alu1 68 37 68 37 1 a0
rlabel alu1 76 33 76 33 1 a0
rlabel alu1 76 45 76 45 1 b0
rlabel alu0 73 57 73 57 1 a0b0_inv
rlabel alu1 1 53 1 53 1 b0
rlabel alu1 84 53 84 53 1 b0
rlabel alu1 52 37 52 37 1 res0
rlabel alu1 60 21 60 21 1 res0
rlabel alu0 76 21 76 21 1 res0_inv
rlabel alu0 60 40 60 40 1 res0_inv
<< end >>
