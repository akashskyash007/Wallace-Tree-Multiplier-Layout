magic
tech scmos
timestamp 1199973079
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -5 40 101 97
<< pwell >>
rect -5 -9 101 40
<< poly >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 81 75 83
rect 66 79 71 81
rect 73 79 75 81
rect 66 77 75 79
rect 53 74 55 77
rect 73 74 75 77
rect 85 81 94 83
rect 85 79 87 81
rect 89 79 94 81
rect 85 77 94 79
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 41 14 43
rect 2 39 7 41
rect 9 39 14 41
rect 2 37 14 39
rect 18 41 30 43
rect 18 39 23 41
rect 25 39 30 41
rect 18 37 30 39
rect 34 41 46 43
rect 34 39 42 41
rect 44 39 46 41
rect 34 37 46 39
rect 50 41 62 43
rect 50 39 52 41
rect 54 39 62 41
rect 50 37 62 39
rect 66 41 78 43
rect 66 39 71 41
rect 73 39 78 41
rect 66 37 78 39
rect 82 37 94 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 5 62 11
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndif >>
rect 2 25 9 34
rect 2 23 4 25
rect 6 23 9 25
rect 2 18 9 23
rect 2 16 4 18
rect 6 16 9 18
rect 2 14 9 16
rect 11 28 21 34
rect 11 26 15 28
rect 17 26 21 28
rect 11 21 21 26
rect 11 19 15 21
rect 17 19 21 21
rect 11 14 21 19
rect 23 18 30 34
rect 23 16 26 18
rect 28 16 30 18
rect 23 14 30 16
rect 34 18 41 34
rect 34 16 36 18
rect 38 16 41 18
rect 34 14 41 16
rect 43 29 53 34
rect 43 27 47 29
rect 49 27 53 29
rect 43 22 53 27
rect 43 20 47 22
rect 49 20 53 22
rect 43 14 53 20
rect 55 18 62 34
rect 55 16 58 18
rect 60 16 62 18
rect 55 14 62 16
rect 66 18 73 34
rect 66 16 68 18
rect 70 16 73 18
rect 66 14 73 16
rect 75 32 85 34
rect 75 30 79 32
rect 81 30 85 32
rect 75 25 85 30
rect 75 23 79 25
rect 81 23 85 25
rect 75 14 85 23
rect 87 25 94 34
rect 87 23 90 25
rect 92 23 94 25
rect 87 18 94 23
rect 87 16 90 18
rect 92 16 94 18
rect 87 14 94 16
rect 13 2 19 14
rect 45 2 51 14
rect 77 2 83 14
<< pdif >>
rect 13 74 19 86
rect 45 77 51 86
rect 45 75 47 77
rect 49 75 51 77
rect 45 74 51 75
rect 77 74 83 86
rect 2 72 9 74
rect 2 70 4 72
rect 6 70 9 72
rect 2 65 9 70
rect 2 63 4 65
rect 6 63 9 65
rect 2 46 9 63
rect 11 58 21 74
rect 11 56 15 58
rect 17 56 21 58
rect 11 51 21 56
rect 11 49 15 51
rect 17 49 21 51
rect 11 46 21 49
rect 23 72 30 74
rect 23 70 26 72
rect 28 70 30 72
rect 23 65 30 70
rect 23 63 26 65
rect 28 63 30 65
rect 23 46 30 63
rect 34 60 41 74
rect 34 58 36 60
rect 38 58 41 60
rect 34 51 41 58
rect 34 49 36 51
rect 38 49 41 51
rect 34 46 41 49
rect 43 70 53 74
rect 43 68 47 70
rect 49 68 53 70
rect 43 46 53 68
rect 55 60 62 74
rect 55 58 58 60
rect 60 58 62 60
rect 55 53 62 58
rect 55 51 58 53
rect 60 51 62 53
rect 55 46 62 51
rect 66 69 73 74
rect 66 67 68 69
rect 70 67 73 69
rect 66 46 73 67
rect 75 57 85 74
rect 75 55 79 57
rect 81 55 85 57
rect 75 50 85 55
rect 75 48 79 50
rect 81 48 85 50
rect 75 46 85 48
rect 87 68 94 74
rect 87 66 90 68
rect 92 66 94 68
rect 87 61 94 66
rect 87 59 90 61
rect 92 59 94 61
rect 87 46 94 59
<< alu1 >>
rect -2 89 98 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 73 87 87 89
rect 89 87 91 89
rect 93 87 98 89
rect -2 86 98 87
rect 3 81 7 86
rect 3 79 4 81
rect 6 79 7 81
rect 3 72 7 79
rect 3 70 4 72
rect 6 70 7 72
rect 3 65 7 70
rect 3 63 4 65
rect 6 63 7 65
rect 3 61 7 63
rect 25 81 29 86
rect 25 79 26 81
rect 28 79 29 81
rect 25 72 29 79
rect 25 70 26 72
rect 28 70 29 72
rect 25 65 29 70
rect 25 63 26 65
rect 28 63 29 65
rect 25 61 29 63
rect 6 41 10 55
rect 6 39 7 41
rect 9 39 10 41
rect 6 38 10 39
rect 21 41 27 46
rect 45 42 51 54
rect 21 39 23 41
rect 25 39 27 41
rect 21 38 27 39
rect 40 41 56 42
rect 40 39 42 41
rect 44 39 52 41
rect 54 39 56 41
rect 40 38 56 39
rect 70 41 74 63
rect 70 39 71 41
rect 73 39 74 41
rect 70 38 74 39
rect 6 34 27 38
rect 45 34 51 38
rect 61 34 74 38
rect 78 57 82 63
rect 78 55 79 57
rect 81 55 82 57
rect 78 50 82 55
rect 78 48 79 50
rect 81 48 82 50
rect 6 33 10 34
rect 78 32 82 48
rect 78 30 79 32
rect 81 30 82 32
rect 14 29 82 30
rect 14 28 47 29
rect 3 25 7 27
rect 3 23 4 25
rect 6 23 7 25
rect 3 18 7 23
rect 3 16 4 18
rect 6 16 7 18
rect 14 26 15 28
rect 17 27 47 28
rect 49 27 82 29
rect 17 26 82 27
rect 14 21 18 26
rect 14 19 15 21
rect 17 19 18 21
rect 46 22 50 26
rect 46 20 47 22
rect 49 20 50 22
rect 78 25 82 26
rect 78 23 79 25
rect 81 23 82 25
rect 14 17 18 19
rect 25 18 29 20
rect 3 9 7 16
rect 3 7 4 9
rect 6 7 7 9
rect 3 2 7 7
rect 25 16 26 18
rect 28 16 29 18
rect 25 9 29 16
rect 25 7 26 9
rect 28 7 29 9
rect 25 2 29 7
rect 35 18 39 20
rect 35 16 36 18
rect 38 16 39 18
rect 46 17 50 20
rect 57 18 61 20
rect 35 9 39 16
rect 35 7 36 9
rect 38 7 39 9
rect 35 2 39 7
rect 57 16 58 18
rect 60 16 61 18
rect 57 9 61 16
rect 57 7 58 9
rect 60 7 61 9
rect 57 2 61 7
rect 67 18 71 20
rect 67 16 68 18
rect 70 16 71 18
rect 78 17 82 23
rect 89 25 93 27
rect 89 23 90 25
rect 92 23 93 25
rect 89 18 93 23
rect 67 9 71 16
rect 67 7 68 9
rect 70 7 71 9
rect 67 2 71 7
rect 89 16 90 18
rect 92 16 93 18
rect 89 9 93 16
rect 89 7 90 9
rect 92 7 93 9
rect 89 2 93 7
rect -2 1 98 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 73 -1 87 1
rect 89 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< alu2 >>
rect -2 89 98 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 71 89
rect 73 87 87 89
rect 89 87 98 89
rect -2 81 98 87
rect -2 79 4 81
rect 6 79 26 81
rect 28 79 98 81
rect -2 76 98 79
rect -2 9 98 12
rect -2 7 4 9
rect 6 7 26 9
rect 28 7 36 9
rect 38 7 58 9
rect 60 7 68 9
rect 70 7 90 9
rect 92 7 98 9
rect -2 1 98 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 71 1
rect 73 -1 87 1
rect 89 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 71 3
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 57 -3 71 -1
rect 89 1 96 3
rect 89 -1 91 1
rect 93 -1 96 1
rect 89 -3 96 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 71 91
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 57 85 71 87
rect 89 89 96 91
rect 89 87 91 89
rect 93 87 96 89
rect 89 85 96 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polyct0 >>
rect 71 79 73 81
rect 87 79 89 81
<< polyct1 >>
rect 7 39 9 41
rect 23 39 25 41
rect 42 39 44 41
rect 52 39 54 41
rect 71 39 73 41
<< ndifct1 >>
rect 4 23 6 25
rect 4 16 6 18
rect 15 26 17 28
rect 15 19 17 21
rect 26 16 28 18
rect 36 16 38 18
rect 47 27 49 29
rect 47 20 49 22
rect 58 16 60 18
rect 68 16 70 18
rect 79 30 81 32
rect 79 23 81 25
rect 90 23 92 25
rect 90 16 92 18
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
rect 67 87 69 89
rect 91 87 93 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 91 -1 93 1
<< pdifct0 >>
rect 47 75 49 77
rect 15 56 17 58
rect 15 49 17 51
rect 36 58 38 60
rect 36 49 38 51
rect 47 68 49 70
rect 58 58 60 60
rect 58 51 60 53
rect 68 67 70 69
rect 90 66 92 68
rect 90 59 92 61
<< pdifct1 >>
rect 4 70 6 72
rect 4 63 6 65
rect 26 70 28 72
rect 26 63 28 65
rect 79 55 81 57
rect 79 48 81 50
<< alu0 >>
rect 69 81 91 82
rect 69 79 71 81
rect 73 79 87 81
rect 89 79 91 81
rect 46 77 50 79
rect 69 78 91 79
rect 46 75 47 77
rect 49 75 50 77
rect 46 70 50 75
rect 46 68 47 70
rect 49 69 93 70
rect 49 68 68 69
rect 46 67 68 68
rect 70 68 93 69
rect 70 67 90 68
rect 46 66 90 67
rect 92 66 93 68
rect 35 60 61 62
rect 14 58 18 60
rect 14 56 15 58
rect 17 56 18 58
rect 14 55 18 56
rect 35 58 36 60
rect 38 58 58 60
rect 60 58 61 60
rect 35 55 39 58
rect 14 51 39 55
rect 14 49 15 51
rect 17 49 18 51
rect 14 47 18 49
rect 35 49 36 51
rect 38 49 39 51
rect 35 47 39 49
rect 57 53 61 58
rect 57 51 58 53
rect 60 51 61 53
rect 57 49 61 51
rect 89 61 93 66
rect 89 59 90 61
rect 92 59 93 61
rect 89 57 93 59
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 71 87 73 89
rect 87 87 89 89
rect 4 79 6 81
rect 26 79 28 81
rect 4 7 6 9
rect 26 7 28 9
rect 36 7 38 9
rect 58 7 60 9
rect 68 7 70 9
rect 90 7 92 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
rect 71 -1 73 1
rect 87 -1 89 1
<< labels >>
rlabel ndifct1 16 20 16 20 6 z
rlabel alu1 16 36 16 36 6 a
rlabel alu1 8 44 8 44 6 a
rlabel alu1 24 28 24 28 6 z
rlabel polyct1 24 40 24 40 6 a
rlabel alu1 40 28 40 28 6 z
rlabel alu1 32 28 32 28 6 z
rlabel alu1 48 24 48 24 6 z
rlabel alu1 64 36 64 36 6 c
rlabel alu1 64 28 64 28 6 z
rlabel alu1 56 28 56 28 6 z
rlabel alu1 48 44 48 44 6 b
rlabel alu1 72 28 72 28 6 z
rlabel alu1 80 40 80 40 6 z
rlabel alu1 72 52 72 52 6 c
rlabel alu2 48 6 48 6 6 vss
rlabel alu2 48 82 48 82 6 vdd
<< end >>
