magic
tech scmos
timestamp 1199203384
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< alu1 >>
rect -2 67 58 72
rect -2 65 8 67
rect 10 65 15 67
rect 17 65 23 67
rect 25 65 31 67
rect 33 65 39 67
rect 41 65 46 67
rect 48 65 58 67
rect -2 64 58 65
rect -2 7 58 8
rect -2 5 8 7
rect 10 5 15 7
rect 17 5 23 7
rect 25 5 31 7
rect 33 5 39 7
rect 41 5 46 7
rect 48 5 58 7
rect -2 0 58 5
<< ptie >>
rect 6 7 50 26
rect 6 5 8 7
rect 10 5 15 7
rect 17 5 23 7
rect 25 5 31 7
rect 33 5 39 7
rect 41 5 46 7
rect 48 5 50 7
rect 6 3 50 5
<< ntie >>
rect 6 67 50 69
rect 6 65 8 67
rect 10 65 15 67
rect 17 65 23 67
rect 25 65 31 67
rect 33 65 39 67
rect 41 65 46 67
rect 48 65 50 67
rect 6 38 50 65
<< ntiect1 >>
rect 8 65 10 67
rect 15 65 17 67
rect 23 65 25 67
rect 31 65 33 67
rect 39 65 41 67
rect 46 65 48 67
<< ptiect1 >>
rect 8 5 10 7
rect 15 5 17 7
rect 23 5 25 7
rect 31 5 33 7
rect 39 5 41 7
rect 46 5 48 7
<< labels >>
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 68 28 68 6 vdd
<< end >>
