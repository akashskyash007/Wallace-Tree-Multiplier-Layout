magic
tech scmos
timestamp 1199202317
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 63 11 67
rect 19 61 21 65
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 21 39
rect 9 35 16 37
rect 18 35 21 37
rect 9 33 21 35
rect 9 30 11 33
rect 19 30 21 33
rect 9 6 11 10
rect 19 6 21 10
<< ndif >>
rect 2 21 9 30
rect 2 19 4 21
rect 6 19 9 21
rect 2 14 9 19
rect 2 12 4 14
rect 6 12 9 14
rect 2 10 9 12
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 10 19 19
rect 21 21 28 30
rect 21 19 24 21
rect 26 19 28 21
rect 21 14 28 19
rect 21 12 24 14
rect 26 12 28 14
rect 21 10 28 12
<< pdif >>
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 16 63
rect 11 59 19 61
rect 11 57 14 59
rect 16 57 19 59
rect 11 52 19 57
rect 11 50 14 52
rect 16 50 19 52
rect 11 42 19 50
rect 21 59 28 61
rect 21 57 24 59
rect 26 57 28 59
rect 21 52 28 57
rect 21 50 24 52
rect 26 50 28 52
rect 21 42 28 50
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 12 59 18 60
rect 12 57 14 59
rect 16 57 18 59
rect 12 55 18 57
rect 2 52 18 55
rect 2 50 14 52
rect 16 50 18 52
rect 2 29 6 50
rect 17 39 23 46
rect 10 37 23 39
rect 10 35 16 37
rect 18 35 23 37
rect 10 33 23 35
rect 2 28 18 29
rect 2 26 14 28
rect 16 26 18 28
rect 2 25 18 26
rect 13 21 18 25
rect 13 19 14 21
rect 16 19 18 21
rect 13 17 18 19
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 10 11 30
rect 19 10 21 30
<< pmos >>
rect 9 42 11 63
rect 19 42 21 61
<< polyct1 >>
rect 16 35 18 37
<< ndifct0 >>
rect 4 19 6 21
rect 4 12 6 14
rect 24 19 26 21
rect 24 12 26 14
<< ndifct1 >>
rect 14 26 16 28
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 59 6 61
rect 24 57 26 59
rect 24 50 26 52
<< pdifct1 >>
rect 14 57 16 59
rect 14 50 16 52
<< alu0 >>
rect 2 61 8 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 6 49 18 50
rect 22 59 28 68
rect 22 57 24 59
rect 26 57 28 59
rect 22 52 28 57
rect 22 50 24 52
rect 26 50 28 52
rect 22 49 28 50
rect 2 21 8 22
rect 2 19 4 21
rect 6 19 8 21
rect 2 14 8 19
rect 22 21 28 22
rect 22 19 24 21
rect 26 19 28 21
rect 2 12 4 14
rect 6 12 8 14
rect 22 14 28 19
rect 22 12 24 14
rect 26 12 28 14
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 36 12 36 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 40 20 40 6 a
rlabel alu1 16 74 16 74 6 vdd
<< end >>
