magic
tech scmos
timestamp 1199201764
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 41 70 43 74
rect 51 70 53 74
rect 9 34 11 42
rect 19 39 21 53
rect 29 47 31 53
rect 41 50 43 53
rect 41 48 47 50
rect 29 45 37 47
rect 29 43 32 45
rect 34 43 37 45
rect 41 46 43 48
rect 45 46 47 48
rect 41 44 47 46
rect 29 41 37 43
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 9 32 15 34
rect 19 33 30 35
rect 9 30 11 32
rect 13 30 15 32
rect 28 30 30 33
rect 35 30 37 41
rect 42 30 44 44
rect 51 39 53 53
rect 49 37 62 39
rect 49 35 58 37
rect 60 35 62 37
rect 49 33 62 35
rect 49 30 51 33
rect 9 28 15 30
rect 9 25 11 28
rect 9 6 11 11
rect 28 6 30 10
rect 35 6 37 10
rect 42 6 44 10
rect 49 6 51 10
<< ndif >>
rect 21 28 28 30
rect 21 26 23 28
rect 25 26 28 28
rect 4 23 9 25
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 11 9 17
rect 11 20 17 25
rect 21 24 28 26
rect 11 11 19 20
rect 13 9 15 11
rect 17 9 19 11
rect 23 10 28 24
rect 30 10 35 30
rect 37 10 42 30
rect 44 10 49 30
rect 51 21 58 30
rect 51 19 54 21
rect 56 19 58 21
rect 51 14 58 19
rect 51 12 54 14
rect 56 12 58 14
rect 51 10 58 12
rect 13 7 19 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 53 19 59
rect 21 61 29 70
rect 21 59 24 61
rect 26 59 29 61
rect 21 53 29 59
rect 31 68 41 70
rect 31 66 35 68
rect 37 66 41 68
rect 31 53 41 66
rect 43 61 51 70
rect 43 59 46 61
rect 48 59 51 61
rect 43 53 51 59
rect 53 68 60 70
rect 53 66 56 68
rect 58 66 60 68
rect 53 60 60 66
rect 53 58 56 60
rect 58 58 60 60
rect 53 53 60 58
rect 11 42 17 53
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 53 7 63
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 2 23 6 42
rect 34 46 38 55
rect 17 45 38 46
rect 17 43 32 45
rect 34 43 38 45
rect 17 42 38 43
rect 42 48 46 55
rect 42 46 43 48
rect 45 47 46 48
rect 45 46 54 47
rect 42 41 54 46
rect 17 37 38 38
rect 17 35 21 37
rect 23 35 38 37
rect 17 34 38 35
rect 2 21 14 23
rect 2 19 4 21
rect 6 19 14 21
rect 2 17 14 19
rect 34 17 38 34
rect 42 33 46 41
rect 58 37 62 39
rect 60 35 62 37
rect 58 31 62 35
rect 50 29 62 31
rect 42 25 62 29
rect 42 17 46 25
rect -2 11 66 12
rect -2 9 15 11
rect 17 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 11 11 25
rect 28 10 30 30
rect 35 10 37 30
rect 42 10 44 30
rect 49 10 51 30
<< pmos >>
rect 9 42 11 70
rect 19 53 21 70
rect 29 53 31 70
rect 41 53 43 70
rect 51 53 53 70
<< polyct0 >>
rect 11 30 13 32
<< polyct1 >>
rect 32 43 34 45
rect 43 46 45 48
rect 21 35 23 37
rect 58 35 60 37
<< ndifct0 >>
rect 23 26 25 28
rect 54 19 56 21
rect 54 12 56 14
<< ndifct1 >>
rect 4 19 6 21
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 14 66 16 68
rect 14 59 16 61
rect 24 59 26 61
rect 35 66 37 68
rect 46 59 48 61
rect 56 66 58 68
rect 56 58 58 60
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 61 18 66
rect 33 66 35 68
rect 37 66 39 68
rect 33 65 39 66
rect 55 66 56 68
rect 58 66 59 68
rect 12 59 14 61
rect 16 59 18 61
rect 12 58 18 59
rect 22 61 50 62
rect 22 59 24 61
rect 26 59 46 61
rect 48 59 50 61
rect 22 58 50 59
rect 55 60 59 66
rect 55 58 56 60
rect 58 58 59 60
rect 22 54 26 58
rect 55 56 59 58
rect 10 50 26 54
rect 10 32 14 50
rect 10 30 11 32
rect 13 30 14 32
rect 10 28 27 30
rect 10 26 23 28
rect 25 26 27 28
rect 21 25 27 26
rect 56 31 58 38
rect 52 21 58 22
rect 52 19 54 21
rect 56 19 58 21
rect 52 14 58 19
rect 52 12 54 14
rect 56 12 58 14
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel ndifct0 24 27 24 27 6 zn
rlabel alu0 36 60 36 60 6 zn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 36 20 36 6 d
rlabel alu1 28 36 28 36 6 d
rlabel alu1 20 44 20 44 6 c
rlabel alu1 28 44 28 44 6 c
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 20 44 20 6 a
rlabel alu1 36 24 36 24 6 d
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 52 36 52 6 c
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 a
rlabel alu1 60 32 60 32 6 a
rlabel alu1 52 44 52 44 6 b
<< end >>
