magic
tech scmos
timestamp 1199202900
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 12 47 14 50
rect 9 45 15 47
rect 9 43 11 45
rect 13 43 15 45
rect 9 41 15 43
rect 10 29 12 41
rect 19 38 21 50
rect 19 36 25 38
rect 19 34 21 36
rect 23 34 25 36
rect 19 32 25 34
rect 20 29 22 32
rect 10 18 12 23
rect 20 18 22 23
<< ndif >>
rect 2 27 10 29
rect 2 25 4 27
rect 6 25 10 27
rect 2 23 10 25
rect 12 27 20 29
rect 12 25 15 27
rect 17 25 20 27
rect 12 23 20 25
rect 22 27 30 29
rect 22 25 26 27
rect 28 25 30 27
rect 22 23 30 25
<< pdif >>
rect 7 64 12 70
rect 5 62 12 64
rect 5 60 7 62
rect 9 60 12 62
rect 5 58 12 60
rect 7 50 12 58
rect 14 50 19 70
rect 21 68 30 70
rect 21 66 26 68
rect 28 66 30 68
rect 21 61 30 66
rect 21 59 26 61
rect 28 59 30 61
rect 21 50 30 59
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 62 11 63
rect 2 60 7 62
rect 9 60 11 62
rect 2 59 11 60
rect 2 37 6 59
rect 18 50 22 55
rect 10 46 22 50
rect 10 45 14 46
rect 10 43 11 45
rect 13 43 14 45
rect 10 41 14 43
rect 26 39 30 47
rect 2 33 14 37
rect 18 36 30 39
rect 18 34 21 36
rect 23 34 30 36
rect 18 33 30 34
rect 10 28 14 33
rect 10 27 19 28
rect 10 25 15 27
rect 17 25 19 27
rect 10 24 19 25
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 10 23 12 29
rect 20 23 22 29
<< pmos >>
rect 12 50 14 70
rect 19 50 21 70
<< polyct1 >>
rect 11 43 13 45
rect 21 34 23 36
<< ndifct0 >>
rect 4 25 6 27
rect 26 25 28 27
<< ndifct1 >>
rect 15 25 17 27
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 26 66 28 68
rect 26 59 28 61
<< pdifct1 >>
rect 7 60 9 62
<< alu0 >>
rect 25 66 26 68
rect 28 66 29 68
rect 25 61 29 66
rect 25 59 26 61
rect 28 59 29 61
rect 25 57 29 59
rect 3 27 7 29
rect 3 25 4 27
rect 6 25 7 27
rect 3 12 7 25
rect 25 27 29 29
rect 25 25 26 27
rect 28 25 29 27
rect 25 12 29 25
<< labels >>
rlabel alu1 4 48 4 48 6 z
rlabel alu1 12 28 12 28 6 z
rlabel polyct1 12 44 12 44 6 b
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 20 52 20 52 6 b
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 40 28 40 6 a
<< end >>
