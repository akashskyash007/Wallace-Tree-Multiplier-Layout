magic
tech scmos
timestamp 1199201687
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 9 66 11 70
rect 20 54 22 59
rect 30 54 32 59
rect 9 35 11 38
rect 20 35 22 46
rect 30 43 32 46
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 29 37 35 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 9 26 11 29
rect 22 21 24 29
rect 29 21 31 37
rect 9 7 11 12
rect 22 9 24 14
rect 29 9 31 14
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 16 9 22
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 21 19 26
rect 11 14 22 21
rect 24 14 29 21
rect 31 18 38 21
rect 31 16 34 18
rect 36 16 38 18
rect 31 14 38 16
rect 11 12 19 14
rect 13 7 19 12
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 18 66
rect 11 62 14 64
rect 16 62 18 64
rect 11 57 18 62
rect 32 65 38 67
rect 32 63 34 65
rect 36 63 38 65
rect 32 61 38 63
rect 11 55 14 57
rect 16 55 18 57
rect 11 54 18 55
rect 34 54 38 61
rect 11 46 20 54
rect 22 50 30 54
rect 22 48 25 50
rect 27 48 30 50
rect 22 46 30 48
rect 32 46 38 54
rect 11 38 18 46
<< alu1 >>
rect -2 67 42 72
rect -2 65 24 67
rect 26 65 42 67
rect -2 64 34 65
rect 36 64 42 65
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 2 40 4 42
rect 6 40 7 42
rect 2 38 7 40
rect 2 24 6 38
rect 34 42 38 51
rect 25 41 38 42
rect 25 39 31 41
rect 33 39 38 41
rect 25 38 38 39
rect 17 33 31 34
rect 17 31 21 33
rect 23 31 31 33
rect 17 30 31 31
rect 2 22 4 24
rect 2 19 6 22
rect 25 22 31 30
rect 2 16 14 19
rect 2 14 4 16
rect 6 14 14 16
rect 2 13 14 14
rect -2 7 42 8
rect -2 5 15 7
rect 17 5 42 7
rect -2 0 42 5
<< ntie >>
rect 22 67 28 69
rect 22 65 24 67
rect 26 65 28 67
rect 22 61 28 65
<< nmos >>
rect 9 12 11 26
rect 22 14 24 21
rect 29 14 31 21
<< pmos >>
rect 9 38 11 66
rect 20 46 22 54
rect 30 46 32 54
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 31 39 33 41
rect 21 31 23 33
<< ndifct0 >>
rect 34 16 36 18
<< ndifct1 >>
rect 4 22 6 24
rect 4 14 6 16
rect 15 5 17 7
<< ntiect1 >>
rect 24 65 26 67
<< pdifct0 >>
rect 14 62 16 64
rect 34 63 36 64
rect 14 55 16 57
rect 25 48 27 50
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 34 64 36 65
<< alu0 >>
rect 12 62 14 64
rect 16 62 18 64
rect 32 63 34 64
rect 36 63 38 64
rect 32 62 38 63
rect 12 57 18 62
rect 12 55 14 57
rect 16 55 18 57
rect 12 54 18 55
rect 10 50 29 51
rect 10 48 25 50
rect 27 48 29 50
rect 10 47 29 48
rect 10 33 14 47
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 6 19 7 26
rect 10 22 22 26
rect 18 19 22 22
rect 18 18 38 19
rect 18 16 34 18
rect 36 16 38 18
rect 18 15 38 16
<< labels >>
rlabel alu0 12 36 12 36 6 zn
rlabel alu0 28 17 28 17 6 zn
rlabel alu0 19 49 19 49 6 zn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 20 32 20 32 6 a
rlabel alu1 28 28 28 28 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 36 48 36 48 6 b
<< end >>
