magic
tech scmos
timestamp 1199202759
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 60 11 65
rect 21 60 23 65
rect 31 60 33 65
rect 45 64 47 69
rect 9 32 11 50
rect 21 39 23 50
rect 31 39 33 50
rect 45 49 47 52
rect 41 47 47 49
rect 41 45 43 47
rect 45 45 47 47
rect 41 43 47 45
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 31 37 41 39
rect 31 35 37 37
rect 39 35 41 37
rect 31 33 41 35
rect 9 30 15 32
rect 9 28 11 30
rect 13 29 15 30
rect 13 28 17 29
rect 9 26 17 28
rect 15 23 17 26
rect 22 23 24 33
rect 31 29 33 33
rect 45 30 47 43
rect 29 26 33 29
rect 29 23 31 26
rect 45 19 47 24
rect 15 8 17 13
rect 22 8 24 13
rect 29 8 31 13
<< ndif >>
rect 35 24 45 30
rect 47 28 54 30
rect 47 26 50 28
rect 52 26 54 28
rect 47 24 54 26
rect 35 23 43 24
rect 8 20 15 23
rect 8 18 10 20
rect 12 18 15 20
rect 8 16 15 18
rect 10 13 15 16
rect 17 13 22 23
rect 24 13 29 23
rect 31 19 43 23
rect 31 17 37 19
rect 39 17 43 19
rect 31 13 43 17
<< pdif >>
rect 35 60 45 64
rect 4 56 9 60
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 11 58 21 60
rect 11 56 15 58
rect 17 56 21 58
rect 11 50 21 56
rect 23 54 31 60
rect 23 52 26 54
rect 28 52 31 54
rect 23 50 31 52
rect 33 58 45 60
rect 33 56 36 58
rect 38 56 45 58
rect 33 52 45 56
rect 47 58 52 64
rect 47 56 54 58
rect 47 54 50 56
rect 52 54 54 56
rect 47 52 54 54
rect 33 50 39 52
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 54 7 56
rect 25 54 29 56
rect 2 52 4 54
rect 6 52 7 54
rect 2 46 7 52
rect 25 52 26 54
rect 28 52 29 54
rect 25 46 29 52
rect 42 47 46 63
rect 42 46 43 47
rect 2 42 29 46
rect 33 45 43 46
rect 45 45 46 47
rect 33 42 46 45
rect 2 21 6 42
rect 19 37 31 38
rect 19 35 21 37
rect 23 35 31 37
rect 19 34 31 35
rect 10 30 14 32
rect 10 28 11 30
rect 13 29 14 30
rect 26 31 31 34
rect 13 28 22 29
rect 10 25 22 28
rect 26 25 38 31
rect 2 20 14 21
rect 2 18 10 20
rect 12 18 14 20
rect 2 17 14 18
rect 18 17 22 25
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 45 24 47 30
rect 15 13 17 23
rect 22 13 24 23
rect 29 13 31 23
<< pmos >>
rect 9 50 11 60
rect 21 50 23 60
rect 31 50 33 60
rect 45 52 47 64
<< polyct0 >>
rect 37 35 39 37
<< polyct1 >>
rect 43 45 45 47
rect 21 35 23 37
rect 11 28 13 30
<< ndifct0 >>
rect 50 26 52 28
rect 37 17 39 19
<< ndifct1 >>
rect 10 18 12 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 15 56 17 58
rect 36 56 38 58
rect 50 54 52 56
<< pdifct1 >>
rect 4 52 6 54
rect 26 52 28 54
<< alu0 >>
rect 14 58 18 68
rect 14 56 15 58
rect 17 56 18 58
rect 35 58 39 68
rect 35 56 36 58
rect 38 56 39 58
rect 14 54 18 56
rect 35 54 39 56
rect 49 56 53 58
rect 49 54 50 56
rect 52 54 53 56
rect 49 38 53 54
rect 35 37 53 38
rect 35 35 37 37
rect 39 35 53 37
rect 35 34 53 35
rect 49 28 53 34
rect 49 26 50 28
rect 52 26 53 28
rect 49 24 53 26
rect 36 19 40 21
rect 36 17 37 19
rect 39 17 40 19
rect 36 12 40 17
<< labels >>
rlabel alu0 44 36 44 36 6 an
rlabel alu0 51 41 51 41 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 c
rlabel alu1 12 28 12 28 6 c
rlabel alu1 20 44 20 44 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 32 28 32 6 b
rlabel alu1 36 28 36 28 6 b
rlabel alu1 36 44 36 44 6 a
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 56 44 56 6 a
<< end >>
