magic
tech scmos
timestamp 1199203349
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 12 61 14 65
rect 12 38 14 42
rect 4 36 14 38
rect 4 34 6 36
rect 8 34 14 36
rect 4 32 14 34
rect 12 29 14 32
rect 12 15 14 19
<< ndif >>
rect 3 27 12 29
rect 3 25 6 27
rect 8 25 12 27
rect 3 19 12 25
rect 14 27 22 29
rect 14 25 18 27
rect 20 25 22 27
rect 14 19 22 25
rect 3 17 6 19
rect 8 17 10 19
rect 3 11 10 17
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
<< pdif >>
rect 3 69 10 72
rect 3 67 6 69
rect 8 67 10 69
rect 3 62 10 67
rect 3 60 6 62
rect 8 61 10 62
rect 8 60 12 61
rect 3 55 12 60
rect 3 53 6 55
rect 8 53 12 55
rect 3 42 12 53
rect 14 53 22 61
rect 14 51 18 53
rect 20 51 22 53
rect 14 46 22 51
rect 14 44 18 46
rect 20 44 22 46
rect 14 42 22 44
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 69 26 79
rect -2 68 6 69
rect 8 68 26 69
rect 17 53 22 63
rect 17 51 18 53
rect 20 51 22 53
rect 17 47 22 51
rect 2 46 22 47
rect 2 44 18 46
rect 20 44 22 46
rect 2 41 22 44
rect 17 27 22 41
rect 17 25 18 27
rect 20 25 22 27
rect 17 17 22 25
rect -2 11 26 12
rect -2 9 6 11
rect 8 9 26 11
rect -2 1 26 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 12 19 14 29
<< pmos >>
rect 12 42 14 61
<< polyct0 >>
rect 6 34 8 36
<< ndifct0 >>
rect 6 25 8 27
rect 6 17 8 19
<< ndifct1 >>
rect 18 25 20 27
rect 6 9 8 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct0 >>
rect 6 67 8 68
rect 6 60 8 62
rect 6 53 8 55
<< pdifct1 >>
rect 6 68 8 69
rect 18 51 20 53
rect 18 44 20 46
<< alu0 >>
rect 5 67 6 68
rect 8 67 9 68
rect 5 62 9 67
rect 5 60 6 62
rect 8 60 9 62
rect 5 55 9 60
rect 5 53 6 55
rect 8 53 9 55
rect 5 51 9 53
rect 4 36 10 37
rect 4 34 6 36
rect 8 34 10 36
rect 4 27 10 34
rect 4 25 6 27
rect 8 25 10 27
rect 4 19 10 25
rect 4 17 6 19
rect 8 17 10 19
rect 4 12 10 17
<< labels >>
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 44 12 44 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 40 20 40 6 z
<< end >>
