magic
tech scmos
timestamp 1199203473
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 13 69 35 71
rect 43 70 45 74
rect 50 70 52 74
rect 13 61 15 69
rect 23 61 25 65
rect 33 61 35 69
rect 13 40 15 43
rect 9 38 17 40
rect 23 39 25 43
rect 9 36 11 38
rect 13 36 17 38
rect 9 34 17 36
rect 2 28 8 30
rect 2 26 4 28
rect 6 26 8 28
rect 2 24 8 26
rect 15 25 17 34
rect 22 37 28 39
rect 33 38 35 43
rect 43 39 45 42
rect 50 39 52 42
rect 22 35 24 37
rect 26 35 28 37
rect 22 33 28 35
rect 39 37 45 39
rect 49 37 55 39
rect 25 25 27 33
rect 39 30 41 37
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 49 30 51 33
rect 35 28 41 30
rect 45 28 51 30
rect 35 25 37 28
rect 45 25 47 28
rect 4 8 6 24
rect 56 20 62 22
rect 56 18 58 20
rect 60 18 62 20
rect 56 16 62 18
rect 15 12 17 16
rect 25 12 27 16
rect 35 8 37 16
rect 45 12 47 16
rect 56 8 58 16
rect 4 6 58 8
<< ndif >>
rect 10 22 15 25
rect 8 20 15 22
rect 8 18 10 20
rect 12 18 15 20
rect 8 16 15 18
rect 17 20 25 25
rect 17 18 20 20
rect 22 18 25 20
rect 17 16 25 18
rect 27 23 35 25
rect 27 21 30 23
rect 32 21 35 23
rect 27 16 35 21
rect 37 21 45 25
rect 37 19 40 21
rect 42 19 45 21
rect 37 16 45 19
rect 47 22 52 25
rect 47 20 54 22
rect 47 18 50 20
rect 52 18 54 20
rect 47 16 54 18
<< pdif >>
rect 38 61 43 70
rect 8 55 13 61
rect 6 53 13 55
rect 6 51 8 53
rect 10 51 13 53
rect 6 49 13 51
rect 8 43 13 49
rect 15 59 23 61
rect 15 57 18 59
rect 20 57 23 59
rect 15 52 23 57
rect 15 50 18 52
rect 20 50 23 52
rect 15 43 23 50
rect 25 54 33 61
rect 25 52 28 54
rect 30 52 33 54
rect 25 47 33 52
rect 25 45 28 47
rect 30 45 33 47
rect 25 43 33 45
rect 35 53 43 61
rect 35 51 38 53
rect 40 51 43 53
rect 35 43 43 51
rect 38 42 43 43
rect 45 42 50 70
rect 52 68 60 70
rect 52 66 55 68
rect 57 66 60 68
rect 52 61 60 66
rect 52 59 55 61
rect 57 59 60 61
rect 52 42 60 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 36 53 62 54
rect 36 51 38 53
rect 40 51 62 53
rect 36 50 62 51
rect 10 42 23 46
rect 10 38 14 42
rect 10 36 11 38
rect 13 36 14 38
rect 10 33 14 36
rect 18 37 31 38
rect 18 35 24 37
rect 26 35 31 37
rect 18 34 31 35
rect 18 25 22 34
rect 58 30 62 50
rect 41 26 62 30
rect 41 22 45 26
rect 38 21 45 22
rect 38 19 40 21
rect 42 19 45 21
rect 38 18 45 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 15 16 17 25
rect 25 16 27 25
rect 35 16 37 25
rect 45 16 47 25
<< pmos >>
rect 13 43 15 61
rect 23 43 25 61
rect 33 43 35 61
rect 43 42 45 70
rect 50 42 52 70
<< polyct0 >>
rect 4 26 6 28
rect 51 35 53 37
rect 58 18 60 20
<< polyct1 >>
rect 11 36 13 38
rect 24 35 26 37
<< ndifct0 >>
rect 10 18 12 20
rect 20 18 22 20
rect 30 21 32 23
rect 50 18 52 20
<< ndifct1 >>
rect 40 19 42 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 8 51 10 53
rect 18 57 20 59
rect 18 50 20 52
rect 28 52 30 54
rect 28 45 30 47
rect 55 66 57 68
rect 55 59 57 61
<< pdifct1 >>
rect 38 51 40 53
<< alu0 >>
rect 16 59 22 68
rect 16 57 18 59
rect 20 57 22 59
rect 53 66 55 68
rect 57 66 59 68
rect 53 61 59 66
rect 53 59 55 61
rect 57 59 59 61
rect 53 58 59 59
rect 2 53 12 54
rect 2 51 8 53
rect 10 51 12 53
rect 2 50 12 51
rect 16 52 22 57
rect 16 50 18 52
rect 20 50 22 52
rect 2 30 6 50
rect 16 49 22 50
rect 27 54 31 56
rect 27 52 28 54
rect 30 52 31 54
rect 27 47 31 52
rect 27 45 28 47
rect 30 46 31 47
rect 30 45 38 46
rect 27 42 38 45
rect 34 38 38 42
rect 34 37 55 38
rect 34 35 51 37
rect 53 35 55 37
rect 34 34 55 35
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 34 30 38 34
rect 29 26 38 30
rect 29 23 33 26
rect 2 20 14 21
rect 2 18 10 20
rect 12 18 14 20
rect 2 17 14 18
rect 19 20 23 22
rect 19 18 20 20
rect 22 18 23 20
rect 29 21 30 23
rect 32 21 33 23
rect 29 19 33 21
rect 48 20 62 21
rect 48 18 50 20
rect 52 18 58 20
rect 60 18 62 20
rect 19 12 23 18
rect 48 17 62 18
<< labels >>
rlabel alu0 8 19 8 19 6 bn
rlabel alu0 4 35 4 35 6 bn
rlabel alu0 7 52 7 52 6 bn
rlabel alu0 29 49 29 49 6 an
rlabel alu0 31 24 31 24 6 an
rlabel alu0 55 19 55 19 6 bn
rlabel alu0 44 36 44 36 6 an
rlabel alu1 12 36 12 36 6 b
rlabel alu1 28 36 28 36 6 a
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 44 20 44 6 b
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 28 44 28 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 z
rlabel alu1 60 40 60 40 6 z
rlabel alu1 52 52 52 52 6 z
<< end >>
