magic
tech scmos
timestamp 1199469801
<< ab >>
rect 0 0 40 100
<< nwell >>
rect -2 48 42 104
<< pwell >>
rect -2 -4 42 48
<< poly >>
rect 13 76 15 81
rect 25 76 27 81
rect 13 53 15 56
rect 13 51 21 53
rect 13 49 17 51
rect 19 49 21 51
rect 13 47 21 49
rect 15 33 17 47
rect 25 43 27 56
rect 23 41 33 43
rect 23 39 29 41
rect 31 39 33 41
rect 23 37 33 39
rect 23 33 25 37
rect 15 11 17 16
rect 23 11 25 16
<< ndif >>
rect 7 31 15 33
rect 7 29 9 31
rect 11 29 15 31
rect 7 23 15 29
rect 7 21 9 23
rect 11 21 15 23
rect 7 19 15 21
rect 10 16 15 19
rect 17 16 23 33
rect 25 21 34 33
rect 25 19 29 21
rect 31 19 34 21
rect 25 16 34 19
<< pdif >>
rect 4 71 13 76
rect 4 69 7 71
rect 9 69 13 71
rect 4 56 13 69
rect 15 71 25 76
rect 15 69 19 71
rect 21 69 25 71
rect 15 61 25 69
rect 15 59 19 61
rect 21 59 25 61
rect 15 56 25 59
rect 27 71 36 76
rect 27 69 31 71
rect 33 69 36 71
rect 27 61 36 69
rect 27 59 31 61
rect 33 59 36 61
rect 27 56 36 59
<< alu1 >>
rect -2 95 42 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 42 95
rect -2 88 42 93
rect 6 71 10 88
rect 6 69 7 71
rect 9 69 10 71
rect 6 67 10 69
rect 18 71 22 73
rect 18 69 19 71
rect 21 69 22 71
rect 18 63 22 69
rect 8 61 22 63
rect 8 59 19 61
rect 21 59 22 61
rect 8 57 22 59
rect 30 71 34 88
rect 30 69 31 71
rect 33 69 34 71
rect 30 61 34 69
rect 30 59 31 61
rect 33 59 34 61
rect 30 57 34 59
rect 8 31 12 57
rect 16 51 32 53
rect 16 49 17 51
rect 19 49 32 51
rect 16 47 32 49
rect 18 37 22 47
rect 28 41 32 43
rect 28 39 29 41
rect 31 39 32 41
rect 28 33 32 39
rect 8 29 9 31
rect 11 29 12 31
rect 8 23 12 29
rect 18 27 32 33
rect 8 21 9 23
rect 11 21 12 23
rect 8 17 12 21
rect 28 21 32 23
rect 28 19 29 21
rect 31 19 32 21
rect 28 12 32 19
rect -2 7 42 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 42 7
rect -2 0 42 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 15 16 17 33
rect 23 16 25 33
<< pmos >>
rect 13 56 15 76
rect 25 56 27 76
<< polyct1 >>
rect 17 49 19 51
rect 29 39 31 41
<< ndifct1 >>
rect 9 29 11 31
rect 9 21 11 23
rect 29 19 31 21
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 7 69 9 71
rect 19 69 21 71
rect 19 59 21 61
rect 31 69 33 71
rect 31 59 33 61
<< labels >>
rlabel alu1 10 40 10 40 6 z
rlabel ptiect1 20 6 20 6 6 vss
rlabel alu1 20 30 20 30 6 a
rlabel alu1 20 45 20 45 6 b
rlabel alu1 20 65 20 65 6 z
rlabel ntiect1 20 94 20 94 6 vdd
rlabel alu1 30 35 30 35 6 a
rlabel alu1 30 50 30 50 6 b
<< end >>
