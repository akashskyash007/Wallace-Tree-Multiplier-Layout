magic
tech scmos
timestamp 1199202992
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 9 69 11 74
rect 16 69 18 74
rect 27 61 29 65
rect 37 61 39 65
rect 9 36 11 49
rect 16 46 18 49
rect 16 44 23 46
rect 16 42 19 44
rect 21 42 23 44
rect 16 40 23 42
rect 9 34 15 36
rect 9 32 11 34
rect 13 32 15 34
rect 9 30 15 32
rect 10 22 12 30
rect 20 22 22 40
rect 27 36 29 49
rect 37 46 39 49
rect 37 44 46 46
rect 37 42 42 44
rect 44 42 46 44
rect 37 40 46 42
rect 26 34 32 36
rect 26 32 28 34
rect 30 32 32 34
rect 26 30 32 32
rect 30 26 32 30
rect 37 26 39 40
rect 10 11 12 16
rect 20 11 22 16
rect 30 11 32 16
rect 37 11 39 16
<< ndif >>
rect 24 22 30 26
rect 2 16 10 22
rect 12 20 20 22
rect 12 18 15 20
rect 17 18 20 20
rect 12 16 20 18
rect 22 20 30 22
rect 22 18 25 20
rect 27 18 30 20
rect 22 16 30 18
rect 32 16 37 26
rect 39 24 46 26
rect 39 22 42 24
rect 44 22 46 24
rect 39 20 46 22
rect 39 16 44 20
rect 2 11 8 16
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
<< pdif >>
rect 40 71 46 73
rect 40 69 42 71
rect 44 69 46 71
rect 4 62 9 69
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 53 9 58
rect 2 51 4 53
rect 6 51 9 53
rect 2 49 9 51
rect 11 49 16 69
rect 18 61 25 69
rect 40 67 46 69
rect 41 61 46 67
rect 18 59 21 61
rect 23 59 27 61
rect 18 49 27 59
rect 29 53 37 61
rect 29 51 32 53
rect 34 51 37 53
rect 29 49 37 51
rect 39 49 46 61
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 71 50 79
rect -2 69 42 71
rect 44 69 50 71
rect -2 68 50 69
rect 2 60 6 63
rect 2 58 4 60
rect 2 53 6 58
rect 2 51 4 53
rect 2 23 6 51
rect 33 58 46 63
rect 10 50 23 54
rect 10 34 14 50
rect 42 46 46 58
rect 10 32 11 34
rect 13 32 14 34
rect 10 30 14 32
rect 25 34 31 38
rect 25 32 28 34
rect 30 32 31 34
rect 41 44 46 46
rect 41 42 42 44
rect 44 42 46 44
rect 41 40 46 42
rect 25 31 31 32
rect 18 25 31 31
rect 2 21 14 23
rect 2 20 19 21
rect 2 18 15 20
rect 17 18 19 20
rect 2 17 19 18
rect -2 11 50 12
rect -2 9 4 11
rect 6 9 50 11
rect -2 1 50 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 10 16 12 22
rect 20 16 22 22
rect 30 16 32 26
rect 37 16 39 26
<< pmos >>
rect 9 49 11 69
rect 16 49 18 69
rect 27 49 29 61
rect 37 49 39 61
<< polyct0 >>
rect 19 42 21 44
<< polyct1 >>
rect 11 32 13 34
rect 42 42 44 44
rect 28 32 30 34
<< ndifct0 >>
rect 25 18 27 20
rect 42 22 44 24
<< ndifct1 >>
rect 15 18 17 20
rect 4 9 6 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 21 59 23 61
rect 32 51 34 53
<< pdifct1 >>
rect 42 69 44 71
rect 4 58 6 60
rect 4 51 6 53
<< alu0 >>
rect 6 50 7 62
rect 19 61 25 68
rect 19 59 21 61
rect 23 59 25 61
rect 19 58 25 59
rect 31 53 35 55
rect 31 51 32 53
rect 34 51 35 53
rect 31 45 35 51
rect 17 44 38 45
rect 17 42 19 44
rect 21 42 38 44
rect 17 41 38 42
rect 34 36 38 41
rect 34 32 45 36
rect 41 24 45 32
rect 41 22 42 24
rect 44 22 45 24
rect 23 20 29 21
rect 41 20 45 22
rect 23 18 25 20
rect 27 18 29 20
rect 23 12 29 18
<< labels >>
rlabel alu0 33 48 33 48 6 nd
rlabel alu0 43 28 43 28 6 nd
rlabel alu0 27 43 27 43 6 nd
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel alu1 12 40 12 40 6 c
rlabel alu1 20 52 20 52 6 c
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 32 28 32 6 a
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 44 52 44 52 6 b
rlabel alu1 36 60 36 60 6 b
<< end >>
