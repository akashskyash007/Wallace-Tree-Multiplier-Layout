magic
tech scmos
timestamp 1199202875
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 27 70 29 74
rect 34 70 36 74
rect 44 70 46 74
rect 51 70 53 74
rect 61 70 63 74
rect 9 39 11 45
rect 2 37 12 39
rect 2 35 4 37
rect 6 35 12 37
rect 2 33 12 35
rect 16 35 18 45
rect 27 35 29 45
rect 34 42 36 45
rect 44 42 46 45
rect 34 40 46 42
rect 40 38 46 40
rect 40 36 42 38
rect 44 36 46 38
rect 16 33 36 35
rect 40 34 46 36
rect 10 30 12 33
rect 20 30 22 33
rect 34 30 36 33
rect 51 30 53 45
rect 61 39 63 42
rect 57 37 63 39
rect 57 35 59 37
rect 61 35 63 37
rect 57 33 63 35
rect 61 30 63 33
rect 34 28 53 30
rect 44 26 46 28
rect 48 26 50 28
rect 44 24 50 26
rect 61 11 63 16
rect 10 6 12 10
rect 20 6 22 10
<< ndif >>
rect 2 11 10 30
rect 2 9 4 11
rect 6 10 10 11
rect 12 28 20 30
rect 12 26 15 28
rect 17 26 20 28
rect 12 10 20 26
rect 22 11 31 30
rect 56 26 61 30
rect 53 20 61 26
rect 53 18 56 20
rect 58 18 61 20
rect 53 16 61 18
rect 63 28 70 30
rect 63 26 66 28
rect 68 26 70 28
rect 63 21 70 26
rect 63 19 66 21
rect 68 19 70 21
rect 63 16 70 19
rect 22 10 26 11
rect 6 9 8 10
rect 2 7 8 9
rect 24 9 26 10
rect 28 9 31 11
rect 24 7 31 9
<< pdif >>
rect 4 62 9 70
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 53 9 58
rect 2 51 4 53
rect 6 51 9 53
rect 2 49 9 51
rect 4 45 9 49
rect 11 45 16 70
rect 18 68 27 70
rect 18 66 22 68
rect 24 66 27 68
rect 18 61 27 66
rect 18 59 22 61
rect 24 59 27 61
rect 18 45 27 59
rect 29 45 34 70
rect 36 61 44 70
rect 36 59 39 61
rect 41 59 44 61
rect 36 54 44 59
rect 36 52 39 54
rect 41 52 44 54
rect 36 45 44 52
rect 46 45 51 70
rect 53 68 61 70
rect 53 66 56 68
rect 58 66 61 68
rect 53 61 61 66
rect 53 59 56 61
rect 58 59 61 61
rect 53 45 61 59
rect 56 42 61 45
rect 63 55 68 70
rect 63 53 70 55
rect 63 51 66 53
rect 68 51 70 53
rect 63 46 70 51
rect 63 44 66 46
rect 68 44 70 46
rect 63 42 70 44
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 60 7 63
rect 2 58 4 60
rect 6 58 7 60
rect 38 61 46 63
rect 38 59 39 61
rect 41 59 46 61
rect 2 54 7 58
rect 38 57 46 59
rect 38 54 42 57
rect 2 53 39 54
rect 2 51 4 53
rect 6 52 39 53
rect 41 52 42 54
rect 6 51 42 52
rect 2 50 42 51
rect 2 37 7 39
rect 2 35 4 37
rect 6 35 7 37
rect 2 21 7 35
rect 18 29 22 50
rect 50 39 54 47
rect 13 28 22 29
rect 13 26 15 28
rect 17 26 22 28
rect 13 25 22 26
rect 26 38 46 39
rect 26 36 42 38
rect 44 36 46 38
rect 26 33 46 36
rect 50 37 62 39
rect 50 35 59 37
rect 61 35 62 37
rect 50 33 62 35
rect 26 21 30 33
rect 2 17 30 21
rect -2 11 74 12
rect -2 9 4 11
rect 6 9 26 11
rect 28 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 10 10 12 30
rect 20 10 22 30
rect 61 16 63 30
<< pmos >>
rect 9 45 11 70
rect 16 45 18 70
rect 27 45 29 70
rect 34 45 36 70
rect 44 45 46 70
rect 51 45 53 70
rect 61 42 63 70
<< polyct0 >>
rect 46 26 48 28
<< polyct1 >>
rect 4 35 6 37
rect 42 36 44 38
rect 59 35 61 37
<< ndifct0 >>
rect 56 18 58 20
rect 66 26 68 28
rect 66 19 68 21
<< ndifct1 >>
rect 4 9 6 11
rect 15 26 17 28
rect 26 9 28 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 22 66 24 68
rect 22 59 24 61
rect 56 66 58 68
rect 56 59 58 61
rect 66 51 68 53
rect 66 44 68 46
<< pdifct1 >>
rect 4 58 6 60
rect 4 51 6 53
rect 39 59 41 61
rect 39 52 41 54
<< alu0 >>
rect 20 66 22 68
rect 24 66 26 68
rect 20 61 26 66
rect 54 66 56 68
rect 58 66 60 68
rect 20 59 22 61
rect 24 59 26 61
rect 20 58 26 59
rect 54 61 60 66
rect 54 59 56 61
rect 58 59 60 61
rect 54 58 60 59
rect 65 53 69 55
rect 65 51 66 53
rect 68 51 69 53
rect 65 46 69 51
rect 65 44 66 46
rect 68 44 69 46
rect 65 29 69 44
rect 44 28 69 29
rect 44 26 46 28
rect 48 26 66 28
rect 68 26 69 28
rect 44 25 69 26
rect 65 21 69 25
rect 54 20 60 21
rect 54 18 56 20
rect 58 18 60 20
rect 54 12 60 18
rect 65 19 66 21
rect 68 19 69 21
rect 65 17 69 19
<< labels >>
rlabel alu0 56 27 56 27 6 an
rlabel alu0 67 36 67 36 6 an
rlabel alu1 4 28 4 28 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 4 60 4 60 6 z
rlabel alu1 28 28 28 28 6 b
rlabel alu1 20 40 20 40 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 36 36 36 6 b
rlabel alu1 44 36 44 36 6 b
rlabel alu1 52 40 52 40 6 a
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel polyct1 60 36 60 36 6 a
<< end >>
