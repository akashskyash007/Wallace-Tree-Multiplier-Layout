magic
tech scmos
timestamp 1199203442
<< ab >>
rect 0 0 176 80
<< nwell >>
rect -5 36 181 88
<< pwell >>
rect -5 -8 181 36
<< poly >>
rect 22 70 24 74
rect 32 70 34 74
rect 42 70 44 74
rect 52 70 54 74
rect 62 70 64 74
rect 72 70 74 74
rect 82 70 84 74
rect 92 70 94 74
rect 102 70 104 74
rect 112 70 114 74
rect 122 70 124 74
rect 132 70 134 74
rect 142 70 144 74
rect 152 70 154 74
rect 162 70 164 74
rect 22 35 24 42
rect 32 39 34 42
rect 42 39 44 42
rect 32 37 44 39
rect 52 39 54 42
rect 62 39 64 42
rect 72 39 74 42
rect 82 39 84 42
rect 92 39 94 42
rect 102 39 104 42
rect 112 39 114 42
rect 122 39 124 42
rect 132 39 134 42
rect 52 37 58 39
rect 62 37 74 39
rect 32 35 35 37
rect 37 35 40 37
rect 9 33 40 35
rect 56 33 58 37
rect 68 35 70 37
rect 72 35 74 37
rect 68 33 74 35
rect 78 37 94 39
rect 98 37 104 39
rect 110 37 116 39
rect 78 35 80 37
rect 82 35 90 37
rect 78 33 90 35
rect 98 33 100 37
rect 110 35 112 37
rect 114 35 116 37
rect 110 33 116 35
rect 9 30 11 33
rect 19 30 21 33
rect 38 30 40 33
rect 49 29 51 33
rect 56 31 64 33
rect 58 29 60 31
rect 62 29 64 31
rect 71 30 73 33
rect 78 30 80 33
rect 58 27 64 29
rect 9 6 11 10
rect 19 6 21 10
rect 38 8 40 11
rect 49 8 51 11
rect 88 24 90 33
rect 94 31 100 33
rect 94 29 96 31
rect 98 29 100 31
rect 114 30 116 33
rect 121 37 134 39
rect 121 35 127 37
rect 129 35 134 37
rect 142 39 144 42
rect 152 39 154 42
rect 142 37 154 39
rect 162 37 164 42
rect 142 35 145 37
rect 147 35 150 37
rect 121 33 134 35
rect 138 33 150 35
rect 161 35 167 37
rect 161 33 163 35
rect 165 33 167 35
rect 121 30 123 33
rect 131 30 133 33
rect 138 30 140 33
rect 94 27 100 29
rect 95 24 97 27
rect 148 28 150 33
rect 155 31 167 33
rect 155 28 157 31
rect 38 6 51 8
rect 71 6 73 10
rect 78 6 80 10
rect 88 6 90 10
rect 95 6 97 10
rect 114 6 116 10
rect 121 6 123 10
rect 131 6 133 10
rect 138 6 140 10
rect 148 6 150 10
rect 155 6 157 10
<< ndif >>
rect 4 22 9 30
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 4 10 9 16
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 10 19 26
rect 21 28 28 30
rect 21 26 24 28
rect 26 26 28 28
rect 21 24 28 26
rect 21 10 26 24
rect 32 20 38 30
rect 30 13 38 20
rect 30 11 32 13
rect 34 11 38 13
rect 40 29 47 30
rect 40 28 49 29
rect 40 26 43 28
rect 45 26 49 28
rect 40 11 49 26
rect 51 24 56 29
rect 66 24 71 30
rect 51 21 71 24
rect 51 19 60 21
rect 62 19 71 21
rect 51 14 71 19
rect 51 12 60 14
rect 62 12 71 14
rect 51 11 71 12
rect 30 9 36 11
rect 53 10 71 11
rect 73 10 78 30
rect 80 24 85 30
rect 102 24 114 30
rect 80 21 88 24
rect 80 19 83 21
rect 85 19 88 21
rect 80 10 88 19
rect 90 10 95 24
rect 97 14 114 24
rect 97 12 100 14
rect 102 12 109 14
rect 111 12 114 14
rect 97 10 114 12
rect 116 10 121 30
rect 123 21 131 30
rect 123 19 126 21
rect 128 19 131 21
rect 123 10 131 19
rect 133 10 138 30
rect 140 28 145 30
rect 140 14 148 28
rect 140 12 143 14
rect 145 12 148 14
rect 140 10 148 12
rect 150 10 155 28
rect 157 23 162 28
rect 157 21 164 23
rect 157 19 160 21
rect 162 19 164 21
rect 157 17 164 19
rect 157 10 162 17
<< pdif >>
rect 14 68 22 70
rect 14 66 17 68
rect 19 66 22 68
rect 14 42 22 66
rect 24 46 32 70
rect 24 44 27 46
rect 29 44 32 46
rect 24 42 32 44
rect 34 68 42 70
rect 34 66 37 68
rect 39 66 42 68
rect 34 42 42 66
rect 44 46 52 70
rect 44 44 47 46
rect 49 44 52 46
rect 44 42 52 44
rect 54 53 62 70
rect 54 51 57 53
rect 59 51 62 53
rect 54 42 62 51
rect 64 61 72 70
rect 64 59 67 61
rect 69 59 72 61
rect 64 42 72 59
rect 74 53 82 70
rect 74 51 77 53
rect 79 51 82 53
rect 74 42 82 51
rect 84 46 92 70
rect 84 44 87 46
rect 89 44 92 46
rect 84 42 92 44
rect 94 53 102 70
rect 94 51 97 53
rect 99 51 102 53
rect 94 46 102 51
rect 94 44 97 46
rect 99 44 102 46
rect 94 42 102 44
rect 104 61 112 70
rect 104 59 107 61
rect 109 59 112 61
rect 104 54 112 59
rect 104 52 107 54
rect 109 52 112 54
rect 104 42 112 52
rect 114 68 122 70
rect 114 66 117 68
rect 119 66 122 68
rect 114 61 122 66
rect 114 59 117 61
rect 119 59 122 61
rect 114 42 122 59
rect 124 60 132 70
rect 124 58 127 60
rect 129 58 132 60
rect 124 53 132 58
rect 124 51 127 53
rect 129 51 132 53
rect 124 42 132 51
rect 134 68 142 70
rect 134 66 137 68
rect 139 66 142 68
rect 134 61 142 66
rect 134 59 137 61
rect 139 59 142 61
rect 134 42 142 59
rect 144 60 152 70
rect 144 58 147 60
rect 149 58 152 60
rect 144 53 152 58
rect 144 51 147 53
rect 149 51 152 53
rect 144 42 152 51
rect 154 68 162 70
rect 154 66 157 68
rect 159 66 162 68
rect 154 61 162 66
rect 154 59 157 61
rect 159 59 162 61
rect 154 42 162 59
rect 164 62 169 70
rect 164 60 171 62
rect 164 58 167 60
rect 169 58 171 60
rect 164 53 171 58
rect 164 51 167 53
rect 169 51 171 53
rect 164 49 171 51
rect 164 42 169 49
<< alu1 >>
rect -2 81 178 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 178 81
rect -2 68 178 79
rect 10 53 101 54
rect 10 51 57 53
rect 59 51 77 53
rect 79 51 97 53
rect 99 51 101 53
rect 10 50 101 51
rect 10 29 14 50
rect 26 37 38 39
rect 26 35 35 37
rect 37 35 38 37
rect 26 33 38 35
rect 10 28 18 29
rect 10 26 14 28
rect 16 26 18 28
rect 10 25 18 26
rect 34 25 38 33
rect 96 46 101 50
rect 96 44 97 46
rect 99 44 107 46
rect 96 42 107 44
rect 103 22 107 42
rect 113 37 119 46
rect 129 42 166 46
rect 129 38 135 42
rect 114 35 119 37
rect 113 30 119 35
rect 125 37 135 38
rect 125 35 127 37
rect 129 35 135 37
rect 125 34 135 35
rect 139 37 151 38
rect 139 35 145 37
rect 147 35 151 37
rect 139 34 151 35
rect 162 35 166 42
rect 139 30 143 34
rect 113 26 143 30
rect 162 33 163 35
rect 165 33 166 35
rect 162 25 166 33
rect 81 21 111 22
rect 81 19 83 21
rect 85 19 111 21
rect 81 18 111 19
rect -2 11 32 12
rect 34 11 178 12
rect -2 1 178 11
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 178 1
rect -2 -2 178 -1
<< ptie >>
rect 0 1 176 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 176 1
rect 0 -3 176 -1
<< ntie >>
rect 0 81 176 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 176 81
rect 0 77 176 79
<< nmos >>
rect 9 10 11 30
rect 19 10 21 30
rect 38 11 40 30
rect 49 11 51 29
rect 71 10 73 30
rect 78 10 80 30
rect 88 10 90 24
rect 95 10 97 24
rect 114 10 116 30
rect 121 10 123 30
rect 131 10 133 30
rect 138 10 140 30
rect 148 10 150 28
rect 155 10 157 28
<< pmos >>
rect 22 42 24 70
rect 32 42 34 70
rect 42 42 44 70
rect 52 42 54 70
rect 62 42 64 70
rect 72 42 74 70
rect 82 42 84 70
rect 92 42 94 70
rect 102 42 104 70
rect 112 42 114 70
rect 122 42 124 70
rect 132 42 134 70
rect 142 42 144 70
rect 152 42 154 70
rect 162 42 164 70
<< polyct0 >>
rect 70 35 72 37
rect 80 35 82 37
rect 112 35 113 37
rect 60 29 62 31
rect 96 29 98 31
<< polyct1 >>
rect 35 35 37 37
rect 113 35 114 37
rect 127 35 129 37
rect 145 35 147 37
rect 163 33 165 35
<< ndifct0 >>
rect 4 18 6 20
rect 24 26 26 28
rect 32 12 34 13
rect 43 26 45 28
rect 60 19 62 21
rect 60 12 62 14
rect 100 12 102 14
rect 109 12 111 14
rect 126 19 128 21
rect 143 12 145 14
rect 160 19 162 21
<< ndifct1 >>
rect 14 26 16 28
rect 32 11 34 12
rect 83 19 85 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
rect 171 79 173 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
rect 171 -1 173 1
<< pdifct0 >>
rect 17 66 19 68
rect 27 44 29 46
rect 37 66 39 68
rect 47 44 49 46
rect 67 59 69 61
rect 87 44 89 46
rect 107 59 109 61
rect 107 52 109 54
rect 117 66 119 68
rect 117 59 119 61
rect 127 58 129 60
rect 127 51 129 53
rect 137 66 139 68
rect 137 59 139 61
rect 147 58 149 60
rect 147 51 149 53
rect 157 66 159 68
rect 157 59 159 61
rect 167 58 169 60
rect 167 51 169 53
<< pdifct1 >>
rect 57 51 59 53
rect 77 51 79 53
rect 97 51 99 53
rect 97 44 99 46
<< alu0 >>
rect 15 66 17 68
rect 19 66 21 68
rect 15 65 21 66
rect 35 66 37 68
rect 39 66 41 68
rect 35 65 41 66
rect 115 66 117 68
rect 119 66 121 68
rect 2 61 111 62
rect 2 59 67 61
rect 69 59 107 61
rect 109 59 111 61
rect 2 58 111 59
rect 115 61 121 66
rect 135 66 137 68
rect 139 66 141 68
rect 115 59 117 61
rect 119 59 121 61
rect 115 58 121 59
rect 126 60 130 62
rect 126 58 127 60
rect 129 58 130 60
rect 135 61 141 66
rect 155 66 157 68
rect 159 66 161 68
rect 135 59 137 61
rect 139 59 141 61
rect 135 58 141 59
rect 146 60 150 62
rect 146 58 147 60
rect 149 58 150 60
rect 155 61 161 66
rect 155 59 157 61
rect 159 59 161 61
rect 155 58 161 59
rect 166 60 170 62
rect 166 58 167 60
rect 169 58 170 60
rect 2 21 6 58
rect 106 54 111 58
rect 126 54 130 58
rect 146 54 150 58
rect 166 54 170 58
rect 106 52 107 54
rect 109 53 174 54
rect 109 52 127 53
rect 106 51 127 52
rect 129 51 147 53
rect 149 51 167 53
rect 169 51 174 53
rect 106 50 174 51
rect 25 46 92 47
rect 25 44 27 46
rect 29 44 47 46
rect 49 44 87 46
rect 89 44 92 46
rect 25 43 92 44
rect 23 28 27 30
rect 23 26 24 28
rect 26 26 27 28
rect 23 21 27 26
rect 42 28 46 43
rect 68 37 74 43
rect 68 35 70 37
rect 72 35 74 37
rect 68 34 74 35
rect 78 37 84 38
rect 78 35 80 37
rect 82 35 84 37
rect 59 31 63 33
rect 59 30 60 31
rect 42 26 43 28
rect 45 26 46 28
rect 42 24 46 26
rect 49 29 60 30
rect 62 30 63 31
rect 78 30 84 35
rect 62 29 84 30
rect 49 26 84 29
rect 88 33 92 43
rect 88 31 99 33
rect 88 29 96 31
rect 98 29 99 31
rect 88 27 99 29
rect 49 21 53 26
rect 111 37 113 39
rect 111 35 112 37
rect 111 33 113 35
rect 170 22 174 50
rect 2 20 53 21
rect 2 18 4 20
rect 6 18 53 20
rect 2 17 53 18
rect 58 21 64 22
rect 58 19 60 21
rect 62 19 64 21
rect 58 14 64 19
rect 124 21 174 22
rect 124 19 126 21
rect 128 19 160 21
rect 162 19 174 21
rect 124 18 174 19
rect 30 13 36 14
rect 30 12 32 13
rect 34 12 36 13
rect 58 12 60 14
rect 62 12 64 14
rect 97 14 113 15
rect 97 12 100 14
rect 102 12 109 14
rect 111 12 113 14
rect 141 14 147 15
rect 141 12 143 14
rect 145 12 147 14
<< labels >>
rlabel alu0 25 23 25 23 6 an
rlabel alu0 27 19 27 19 6 an
rlabel alu0 44 35 44 35 6 bn
rlabel alu0 66 28 66 28 6 an
rlabel alu0 81 32 81 32 6 an
rlabel alu0 93 30 93 30 6 bn
rlabel alu0 71 40 71 40 6 bn
rlabel alu0 58 45 58 45 6 bn
rlabel alu0 128 56 128 56 6 an
rlabel alu0 108 56 108 56 6 an
rlabel alu0 56 60 56 60 6 an
rlabel alu0 149 20 149 20 6 an
rlabel alu0 148 56 148 56 6 an
rlabel alu0 168 56 168 56 6 an
rlabel alu0 140 52 140 52 6 an
rlabel alu1 28 36 28 36 6 b
rlabel alu1 12 36 12 36 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 32 36 32 6 b
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 88 6 88 6 6 vss
rlabel alu1 100 20 100 20 6 z
rlabel ndifct1 84 20 84 20 6 z
rlabel alu1 92 20 92 20 6 z
rlabel alu1 100 44 100 44 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 92 52 92 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 88 74 88 74 6 vdd
rlabel alu1 108 20 108 20 6 z
rlabel alu1 124 28 124 28 6 a1
rlabel alu1 132 28 132 28 6 a1
rlabel alu1 140 28 140 28 6 a1
rlabel alu1 132 40 132 40 6 a2
rlabel alu1 140 44 140 44 6 a2
rlabel alu1 116 36 116 36 6 a1
rlabel alu1 164 32 164 32 6 a2
rlabel alu1 148 36 148 36 6 a1
rlabel alu1 148 44 148 44 6 a2
rlabel alu1 156 44 156 44 6 a2
<< end >>
