magic
tech scmos
timestamp 1199203708
<< ab >>
rect 0 0 128 80
<< nwell >>
rect -5 36 133 88
<< pwell >>
rect -5 -8 133 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 39 53 41 56
rect 49 53 51 56
rect 39 51 51 53
rect 45 49 47 51
rect 49 49 51 51
rect 45 47 51 49
rect 100 63 102 67
rect 110 63 112 67
rect 100 46 102 49
rect 110 46 112 49
rect 100 44 126 46
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 69 39 71 42
rect 79 39 81 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 29 37 65 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 10 24 12 33
rect 19 29 21 33
rect 37 29 39 37
rect 59 35 61 37
rect 63 35 65 37
rect 59 33 65 35
rect 69 37 75 39
rect 69 35 71 37
rect 73 35 75 37
rect 69 33 75 35
rect 79 37 85 39
rect 79 35 81 37
rect 83 35 85 37
rect 89 38 91 42
rect 89 36 103 38
rect 79 33 85 35
rect 97 34 99 36
rect 101 34 103 36
rect 49 31 55 33
rect 49 29 51 31
rect 53 29 55 31
rect 17 27 21 29
rect 17 24 19 27
rect 27 24 29 29
rect 49 27 55 29
rect 49 24 51 27
rect 72 24 74 33
rect 79 24 81 33
rect 97 32 103 34
rect 99 29 101 32
rect 110 30 112 44
rect 120 42 122 44
rect 124 42 126 44
rect 120 40 126 42
rect 89 24 91 29
rect 37 12 39 16
rect 10 6 12 11
rect 17 6 19 11
rect 27 8 29 11
rect 49 8 51 13
rect 27 6 51 8
rect 99 12 101 16
rect 72 6 74 11
rect 79 6 81 11
rect 89 8 91 11
rect 110 8 112 19
rect 89 6 112 8
<< ndif >>
rect 32 24 37 29
rect 2 11 10 24
rect 12 11 17 24
rect 19 21 27 24
rect 19 19 22 21
rect 24 19 27 21
rect 19 11 27 19
rect 29 22 37 24
rect 29 20 32 22
rect 34 20 37 22
rect 29 16 37 20
rect 39 24 47 29
rect 105 29 110 30
rect 94 24 99 29
rect 39 16 49 24
rect 29 11 34 16
rect 41 14 49 16
rect 41 12 43 14
rect 45 13 49 14
rect 51 22 58 24
rect 51 20 54 22
rect 56 20 58 22
rect 51 18 58 20
rect 51 13 56 18
rect 45 12 47 13
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
rect 41 10 47 12
rect 64 11 72 24
rect 74 11 79 24
rect 81 21 89 24
rect 81 19 84 21
rect 86 19 89 21
rect 81 11 89 19
rect 91 22 99 24
rect 91 20 94 22
rect 96 20 99 22
rect 91 16 99 20
rect 101 20 110 29
rect 101 18 104 20
rect 106 19 110 20
rect 112 28 119 30
rect 112 26 115 28
rect 117 26 119 28
rect 112 24 119 26
rect 112 19 117 24
rect 106 18 108 19
rect 101 16 108 18
rect 91 11 96 16
rect 64 9 66 11
rect 68 9 70 11
rect 64 7 70 9
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 57 9 59
rect 4 42 9 57
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 56 39 66
rect 41 61 49 70
rect 41 59 44 61
rect 46 59 49 61
rect 41 56 49 59
rect 51 68 58 70
rect 51 66 54 68
rect 56 66 58 68
rect 51 61 58 66
rect 64 63 69 70
rect 51 59 54 61
rect 56 59 58 61
rect 51 56 58 59
rect 62 61 69 63
rect 62 59 64 61
rect 66 59 69 61
rect 62 57 69 59
rect 31 42 37 56
rect 64 42 69 57
rect 71 53 79 70
rect 71 51 74 53
rect 76 51 79 53
rect 71 42 79 51
rect 81 53 89 70
rect 81 51 84 53
rect 86 51 89 53
rect 81 46 89 51
rect 81 44 84 46
rect 86 44 89 46
rect 81 42 89 44
rect 91 68 98 70
rect 91 66 94 68
rect 96 66 98 68
rect 91 63 98 66
rect 91 49 100 63
rect 102 53 110 63
rect 102 51 105 53
rect 107 51 110 53
rect 102 49 110 51
rect 112 61 120 63
rect 112 59 115 61
rect 117 59 120 61
rect 112 49 120 59
rect 91 42 98 49
<< alu1 >>
rect -2 81 130 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 130 81
rect -2 68 130 79
rect 2 53 18 54
rect 2 51 14 53
rect 16 51 18 53
rect 2 50 18 51
rect 2 22 6 50
rect 41 51 54 54
rect 41 49 47 51
rect 49 49 54 51
rect 41 48 54 49
rect 2 21 26 22
rect 2 19 22 21
rect 24 19 26 21
rect 2 18 26 19
rect 50 31 54 48
rect 50 29 51 31
rect 53 29 54 31
rect 50 27 54 29
rect 113 50 126 55
rect 122 46 126 50
rect 98 36 111 39
rect 98 34 99 36
rect 101 34 111 36
rect 98 33 111 34
rect 105 26 111 33
rect 121 44 126 46
rect 121 42 122 44
rect 124 42 126 44
rect 121 40 126 42
rect 122 33 126 40
rect -2 11 130 12
rect -2 9 4 11
rect 6 9 66 11
rect 68 9 130 11
rect -2 1 130 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 130 1
rect -2 -2 130 -1
<< ptie >>
rect 0 1 128 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 128 1
rect 0 -3 128 -1
<< ntie >>
rect 0 81 128 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 128 81
rect 0 77 128 79
<< nmos >>
rect 10 11 12 24
rect 17 11 19 24
rect 27 11 29 24
rect 37 16 39 29
rect 49 13 51 24
rect 72 11 74 24
rect 79 11 81 24
rect 89 11 91 24
rect 99 16 101 29
rect 110 19 112 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 56 41 70
rect 49 56 51 70
rect 69 42 71 70
rect 79 42 81 70
rect 89 42 91 70
rect 100 49 102 63
rect 110 49 112 63
<< polyct0 >>
rect 11 35 13 37
rect 21 35 23 37
rect 61 35 63 37
rect 71 35 73 37
rect 81 35 83 37
<< polyct1 >>
rect 47 49 49 51
rect 99 34 101 36
rect 51 29 53 31
rect 122 42 124 44
<< ndifct0 >>
rect 32 20 34 22
rect 43 12 45 14
rect 54 20 56 22
rect 84 19 86 21
rect 94 20 96 22
rect 104 18 106 20
rect 115 26 117 28
<< ndifct1 >>
rect 22 19 24 21
rect 4 9 6 11
rect 66 9 68 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
<< pdifct0 >>
rect 4 59 6 61
rect 24 51 26 53
rect 24 44 26 46
rect 34 66 36 68
rect 44 59 46 61
rect 54 66 56 68
rect 54 59 56 61
rect 64 59 66 61
rect 74 51 76 53
rect 84 51 86 53
rect 84 44 86 46
rect 94 66 96 68
rect 105 51 107 53
rect 115 59 117 61
<< pdifct1 >>
rect 14 51 16 53
<< alu0 >>
rect 32 66 34 68
rect 36 66 38 68
rect 32 65 38 66
rect 52 66 54 68
rect 56 66 58 68
rect 2 61 48 62
rect 2 59 4 61
rect 6 59 44 61
rect 46 59 48 61
rect 2 58 48 59
rect 52 61 58 66
rect 92 66 94 68
rect 96 66 98 68
rect 92 65 98 66
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
rect 62 61 94 62
rect 62 59 64 61
rect 66 59 94 61
rect 62 58 94 59
rect 113 61 119 68
rect 113 59 115 61
rect 117 59 119 61
rect 113 58 119 59
rect 22 53 28 54
rect 22 51 24 53
rect 26 51 28 53
rect 22 47 28 51
rect 10 46 28 47
rect 10 44 24 46
rect 26 44 28 46
rect 10 43 28 44
rect 10 37 14 43
rect 32 38 36 58
rect 90 55 94 58
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 19 37 45 38
rect 19 35 21 37
rect 23 35 45 37
rect 19 34 45 35
rect 10 26 35 30
rect 31 22 35 26
rect 31 20 32 22
rect 34 20 35 22
rect 31 18 35 20
rect 41 23 45 34
rect 62 53 78 54
rect 62 51 74 53
rect 76 51 78 53
rect 62 50 78 51
rect 83 53 87 55
rect 83 51 84 53
rect 86 51 87 53
rect 62 38 66 50
rect 83 46 87 51
rect 59 37 66 38
rect 59 35 61 37
rect 63 35 66 37
rect 59 34 66 35
rect 41 22 58 23
rect 41 20 54 22
rect 56 20 58 22
rect 41 19 58 20
rect 62 22 66 34
rect 70 44 84 46
rect 86 44 87 46
rect 70 42 87 44
rect 90 53 108 55
rect 90 51 105 53
rect 107 51 108 53
rect 70 37 74 42
rect 90 38 94 51
rect 104 46 108 51
rect 104 42 118 46
rect 70 35 71 37
rect 73 35 74 37
rect 70 30 74 35
rect 79 37 94 38
rect 79 35 81 37
rect 83 35 94 37
rect 79 34 94 35
rect 70 26 97 30
rect 114 28 118 42
rect 114 26 115 28
rect 117 26 118 28
rect 93 22 97 26
rect 114 24 118 26
rect 62 21 88 22
rect 62 19 84 21
rect 86 19 88 21
rect 62 18 88 19
rect 93 20 94 22
rect 96 20 97 22
rect 93 18 97 20
rect 103 20 107 22
rect 103 18 104 20
rect 106 18 107 20
rect 41 14 47 15
rect 41 12 43 14
rect 45 12 47 14
rect 103 12 107 18
<< labels >>
rlabel alu0 34 48 34 48 6 cn
rlabel alu0 25 60 25 60 6 cn
rlabel alu0 49 21 49 21 6 cn
rlabel polyct0 72 36 72 36 6 an
rlabel alu0 95 24 95 24 6 an
rlabel alu0 86 36 86 36 6 bn
rlabel alu0 85 48 85 48 6 an
rlabel alu0 78 60 78 60 6 bn
rlabel alu0 116 35 116 35 6 bn
rlabel alu0 106 48 106 48 6 bn
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 52 40 52 40 6 c
rlabel alu1 44 52 44 52 6 c
rlabel alu1 64 6 64 6 6 vss
rlabel alu1 64 74 64 74 6 vdd
rlabel alu1 100 36 100 36 6 a
rlabel alu1 108 32 108 32 6 a
rlabel alu1 124 44 124 44 6 b
rlabel alu1 116 52 116 52 6 b
<< end >>
