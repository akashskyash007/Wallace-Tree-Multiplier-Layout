magic
tech scmos
timestamp 1199203295
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 28 66 30 70
rect 35 66 37 70
rect 42 66 44 70
rect 49 66 51 70
rect 9 57 11 61
rect 9 36 11 45
rect 28 36 30 39
rect 9 34 15 36
rect 9 32 11 34
rect 13 32 15 34
rect 9 30 15 32
rect 19 34 30 36
rect 19 32 21 34
rect 23 32 25 34
rect 19 30 25 32
rect 35 30 37 39
rect 9 21 11 30
rect 19 21 21 30
rect 29 28 37 30
rect 29 26 33 28
rect 35 26 37 28
rect 29 24 37 26
rect 42 27 44 39
rect 49 36 51 39
rect 49 34 58 36
rect 52 32 54 34
rect 56 32 58 34
rect 52 30 58 32
rect 42 25 48 27
rect 29 21 31 24
rect 42 23 44 25
rect 46 23 48 25
rect 42 21 48 23
rect 42 18 44 21
rect 52 18 54 30
rect 9 11 11 15
rect 19 11 21 15
rect 29 10 31 15
rect 42 7 44 12
rect 52 7 54 12
<< ndif >>
rect 2 19 9 21
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 15 19 21
rect 21 19 29 21
rect 21 17 24 19
rect 26 17 29 19
rect 21 15 29 17
rect 31 18 40 21
rect 31 15 42 18
rect 13 9 17 15
rect 33 12 42 15
rect 44 16 52 18
rect 44 14 47 16
rect 49 14 52 16
rect 44 12 52 14
rect 54 12 62 18
rect 13 7 19 9
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
rect 33 7 40 12
rect 56 7 62 12
rect 33 5 35 7
rect 37 5 40 7
rect 33 3 40 5
rect 56 5 58 7
rect 60 5 62 7
rect 56 3 62 5
<< pdif >>
rect 13 59 19 61
rect 13 57 15 59
rect 17 57 19 59
rect 4 51 9 57
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 11 55 19 57
rect 11 45 17 55
rect 23 51 28 66
rect 21 49 28 51
rect 21 47 23 49
rect 25 47 28 49
rect 21 45 28 47
rect 23 39 28 45
rect 30 39 35 66
rect 37 39 42 66
rect 44 39 49 66
rect 51 64 59 66
rect 51 62 54 64
rect 56 62 59 64
rect 51 57 59 62
rect 51 55 54 57
rect 56 55 59 57
rect 51 39 59 55
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 66 67
rect -2 64 66 65
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 45 7 47
rect 2 19 6 45
rect 34 42 38 59
rect 20 38 38 42
rect 42 42 46 51
rect 42 38 57 42
rect 20 34 24 38
rect 53 34 57 38
rect 20 32 21 34
rect 23 32 24 34
rect 20 30 24 32
rect 32 30 47 34
rect 53 32 54 34
rect 56 32 57 34
rect 53 30 57 32
rect 32 28 38 30
rect 32 26 33 28
rect 35 26 38 28
rect 2 17 4 19
rect 32 21 38 26
rect 42 25 62 26
rect 42 23 44 25
rect 46 23 62 25
rect 42 22 62 23
rect 6 17 16 18
rect 2 13 16 17
rect 58 13 62 22
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 15 7
rect 17 5 35 7
rect 37 5 58 7
rect 60 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 15 11 21
rect 19 15 21 21
rect 29 15 31 21
rect 42 12 44 18
rect 52 12 54 18
<< pmos >>
rect 9 45 11 57
rect 28 39 30 66
rect 35 39 37 66
rect 42 39 44 66
rect 49 39 51 66
<< polyct0 >>
rect 11 32 13 34
<< polyct1 >>
rect 21 32 23 34
rect 33 26 35 28
rect 54 32 56 34
rect 44 23 46 25
<< ndifct0 >>
rect 24 17 26 19
rect 47 14 49 16
<< ndifct1 >>
rect 4 17 6 19
rect 15 5 17 7
rect 35 5 37 7
rect 58 5 60 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 15 57 17 59
rect 23 47 25 49
rect 54 62 56 64
rect 54 55 56 57
<< pdifct1 >>
rect 4 47 6 49
<< alu0 >>
rect 14 59 18 64
rect 52 62 54 64
rect 56 62 58 64
rect 14 57 15 59
rect 17 57 18 59
rect 14 55 18 57
rect 11 49 27 50
rect 11 47 23 49
rect 25 47 27 49
rect 11 46 27 47
rect 11 36 15 46
rect 52 57 58 62
rect 52 55 54 57
rect 56 55 58 57
rect 52 54 58 55
rect 10 34 15 36
rect 10 32 11 34
rect 13 32 15 34
rect 10 30 15 32
rect 11 26 15 30
rect 11 22 27 26
rect 6 18 7 21
rect 23 19 27 22
rect 23 17 24 19
rect 26 17 27 19
rect 23 16 51 17
rect 23 14 47 16
rect 49 14 51 16
rect 23 13 51 14
<< labels >>
rlabel alu0 13 36 13 36 6 zn
rlabel alu0 19 48 19 48 6 zn
rlabel alu0 37 15 37 15 6 zn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 28 40 28 40 6 d
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 28 36 28 6 c
rlabel alu1 44 32 44 32 6 c
rlabel alu1 36 52 36 52 6 d
rlabel alu1 44 48 44 48 6 a
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 60 16 60 16 6 b
rlabel alu1 52 24 52 24 6 b
rlabel alu1 52 40 52 40 6 a
<< end >>
