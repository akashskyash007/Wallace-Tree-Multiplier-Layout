magic
tech scmos
timestamp 1199202619
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 66 11 71
rect 19 69 21 74
rect 29 69 31 74
rect 39 66 41 71
rect 49 66 51 71
rect 59 60 61 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 33 39
rect 19 35 27 37
rect 29 35 33 37
rect 19 33 33 35
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 37 51 39
rect 38 35 43 37
rect 45 35 51 37
rect 38 33 51 35
rect 55 37 63 39
rect 55 35 59 37
rect 61 35 63 37
rect 55 33 63 35
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 12 6 14 10
rect 19 6 21 10
rect 31 6 33 10
rect 38 6 40 10
rect 48 6 50 10
rect 55 6 57 10
<< ndif >>
rect 5 28 12 30
rect 5 26 7 28
rect 9 26 12 28
rect 5 21 12 26
rect 5 19 7 21
rect 9 19 12 21
rect 5 17 12 19
rect 7 10 12 17
rect 14 10 19 30
rect 21 14 31 30
rect 21 12 25 14
rect 27 12 31 14
rect 21 10 31 12
rect 33 10 38 30
rect 40 21 48 30
rect 40 19 43 21
rect 45 19 48 21
rect 40 10 48 19
rect 50 10 55 30
rect 57 14 65 30
rect 57 12 60 14
rect 62 12 65 14
rect 57 10 65 12
<< pdif >>
rect 14 66 19 69
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 56 9 62
rect 2 54 4 56
rect 6 54 9 56
rect 2 42 9 54
rect 11 53 19 66
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 66 36 69
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 42 49 62
rect 51 60 56 66
rect 51 53 59 60
rect 51 51 54 53
rect 56 51 59 53
rect 51 42 59 51
rect 61 58 68 60
rect 61 56 64 58
rect 66 56 68 58
rect 61 42 68 56
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 12 53 58 54
rect 12 51 14 53
rect 16 51 34 53
rect 36 51 54 53
rect 56 51 58 53
rect 12 50 58 51
rect 12 47 18 50
rect 2 46 18 47
rect 2 44 14 46
rect 16 44 18 46
rect 2 43 18 44
rect 2 29 6 43
rect 25 42 63 46
rect 10 37 21 39
rect 10 35 11 37
rect 13 35 21 37
rect 10 33 21 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 17 30 21 33
rect 41 30 47 35
rect 57 37 63 42
rect 57 35 59 37
rect 61 35 63 37
rect 57 34 63 35
rect 2 28 11 29
rect 2 26 7 28
rect 9 26 11 28
rect 17 26 47 30
rect 2 25 11 26
rect 5 22 11 25
rect 5 21 47 22
rect 5 19 7 21
rect 9 19 43 21
rect 45 19 47 21
rect 5 18 47 19
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 31 10 33 30
rect 38 10 40 30
rect 48 10 50 30
rect 55 10 57 30
<< pmos >>
rect 9 42 11 66
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 66
rect 49 42 51 66
rect 59 42 61 60
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 43 35 45 37
rect 59 35 61 37
<< ndifct0 >>
rect 25 12 27 14
rect 60 12 62 14
<< ndifct1 >>
rect 7 26 9 28
rect 7 19 9 21
rect 43 19 45 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 62 6 64
rect 4 54 6 56
rect 24 65 26 67
rect 24 58 26 60
rect 44 62 46 64
rect 64 56 66 58
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
rect 34 59 36 61
rect 34 51 36 53
rect 54 51 56 53
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 3 56 7 62
rect 22 67 28 68
rect 22 65 24 67
rect 26 65 28 67
rect 22 60 28 65
rect 43 64 47 68
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 43 62 44 64
rect 46 62 47 64
rect 43 60 47 62
rect 3 54 4 56
rect 6 54 7 56
rect 63 58 67 68
rect 63 56 64 58
rect 66 56 67 58
rect 63 54 67 56
rect 3 52 7 54
rect 23 14 29 15
rect 23 12 25 14
rect 27 12 29 14
rect 58 14 64 15
rect 58 12 60 14
rect 62 12 64 14
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 36 4 36 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 28 28 28 6 b
rlabel alu1 28 40 28 40 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel ndifct1 44 20 44 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 b
rlabel alu1 44 32 44 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 52 44 52 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 36 56 36 56 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 40 60 40 6 a
<< end >>
