magic
tech scmos
timestamp 1199203524
<< ab >>
rect 0 0 184 80
<< nwell >>
rect -5 36 189 88
<< pwell >>
rect -5 -8 189 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 72 53 74
rect 29 69 31 72
rect 39 69 41 72
rect 51 55 53 72
rect 63 70 65 74
rect 73 70 75 74
rect 83 70 85 74
rect 93 70 95 74
rect 116 70 118 74
rect 123 70 125 74
rect 133 70 135 74
rect 151 70 153 74
rect 161 70 163 74
rect 48 53 54 55
rect 48 51 50 53
rect 52 51 54 53
rect 48 49 54 51
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 63 41 65 44
rect 73 41 75 44
rect 9 37 22 39
rect 29 37 41 39
rect 61 39 75 41
rect 83 39 85 42
rect 93 39 95 42
rect 116 39 118 42
rect 61 37 67 39
rect 16 35 18 37
rect 20 35 22 37
rect 16 33 22 35
rect 9 28 11 33
rect 16 31 28 33
rect 16 28 18 31
rect 26 28 28 31
rect 33 28 35 37
rect 61 35 63 37
rect 65 35 67 37
rect 80 37 108 39
rect 80 35 82 37
rect 45 30 47 35
rect 55 33 67 35
rect 55 30 57 33
rect 65 30 67 33
rect 75 33 82 35
rect 102 35 104 37
rect 106 35 108 37
rect 102 33 108 35
rect 112 37 118 39
rect 112 35 114 37
rect 116 35 118 37
rect 123 39 125 42
rect 133 39 135 42
rect 151 39 153 42
rect 161 39 163 42
rect 123 36 126 39
rect 133 37 153 39
rect 157 37 163 39
rect 112 33 118 35
rect 75 30 77 33
rect 86 30 92 32
rect 114 30 116 33
rect 124 30 126 36
rect 137 35 139 37
rect 141 35 148 37
rect 137 33 148 35
rect 157 35 159 37
rect 161 35 163 37
rect 157 33 163 35
rect 146 30 148 33
rect 86 28 88 30
rect 90 28 92 30
rect 86 27 92 28
rect 85 25 97 27
rect 85 22 87 25
rect 95 22 97 25
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
rect 45 8 47 16
rect 55 12 57 16
rect 65 12 67 16
rect 75 8 77 16
rect 133 20 139 22
rect 133 18 135 20
rect 137 18 139 20
rect 158 27 160 33
rect 133 16 139 18
rect 114 11 116 16
rect 124 13 126 16
rect 133 13 135 16
rect 146 14 148 19
rect 124 11 135 13
rect 158 11 160 16
rect 45 6 77 8
rect 85 6 87 10
rect 95 6 97 10
<< ndif >>
rect 37 28 45 30
rect 4 22 9 28
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 16 28
rect 18 26 26 28
rect 18 24 21 26
rect 23 24 26 26
rect 18 16 26 24
rect 28 16 33 28
rect 35 16 45 28
rect 47 28 55 30
rect 47 26 50 28
rect 52 26 55 28
rect 47 16 55 26
rect 57 20 65 30
rect 57 18 60 20
rect 62 18 65 20
rect 57 16 65 18
rect 67 28 75 30
rect 67 26 70 28
rect 72 26 75 28
rect 67 21 75 26
rect 67 19 70 21
rect 72 19 75 21
rect 67 16 75 19
rect 77 22 82 30
rect 109 23 114 30
rect 77 20 85 22
rect 77 18 80 20
rect 82 18 85 20
rect 77 16 85 18
rect 37 11 43 16
rect 37 9 39 11
rect 41 9 43 11
rect 37 7 43 9
rect 80 10 85 16
rect 87 20 95 22
rect 87 18 90 20
rect 92 18 95 20
rect 87 10 95 18
rect 97 13 103 22
rect 107 21 114 23
rect 107 19 109 21
rect 111 19 114 21
rect 107 17 114 19
rect 109 16 114 17
rect 116 28 124 30
rect 116 26 119 28
rect 121 26 124 28
rect 116 16 124 26
rect 126 28 133 30
rect 126 26 129 28
rect 131 26 133 28
rect 126 24 133 26
rect 139 28 146 30
rect 139 26 141 28
rect 143 26 146 28
rect 139 24 146 26
rect 126 16 131 24
rect 141 19 146 24
rect 148 27 156 30
rect 148 19 158 27
rect 97 11 105 13
rect 150 16 158 19
rect 160 22 165 27
rect 160 20 167 22
rect 160 18 163 20
rect 165 18 167 20
rect 160 16 167 18
rect 150 11 156 16
rect 97 10 101 11
rect 99 9 101 10
rect 103 9 105 11
rect 99 7 105 9
rect 150 9 152 11
rect 154 9 156 11
rect 150 7 156 9
<< pdif >>
rect 4 63 9 69
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 53 19 69
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 61 29 69
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 46 39 69
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 63 46 69
rect 41 61 48 63
rect 41 59 44 61
rect 46 59 48 61
rect 41 57 48 59
rect 41 42 46 57
rect 56 68 63 70
rect 56 66 58 68
rect 60 66 63 68
rect 56 61 63 66
rect 56 59 58 61
rect 60 59 63 61
rect 56 44 63 59
rect 65 61 73 70
rect 65 59 68 61
rect 70 59 73 61
rect 65 54 73 59
rect 65 52 68 54
rect 70 52 73 54
rect 65 44 73 52
rect 75 68 83 70
rect 75 66 78 68
rect 80 66 83 68
rect 75 44 83 66
rect 78 42 83 44
rect 85 48 93 70
rect 85 46 88 48
rect 90 46 93 48
rect 85 42 93 46
rect 95 68 116 70
rect 95 66 98 68
rect 100 66 106 68
rect 108 66 116 68
rect 95 61 116 66
rect 95 59 106 61
rect 108 59 116 61
rect 95 42 116 59
rect 118 42 123 70
rect 125 62 133 70
rect 125 60 128 62
rect 130 60 133 62
rect 125 42 133 60
rect 135 64 140 70
rect 135 62 142 64
rect 135 60 138 62
rect 140 60 142 62
rect 135 58 142 60
rect 135 42 140 58
rect 146 54 151 70
rect 144 52 151 54
rect 144 50 146 52
rect 148 50 151 52
rect 144 48 151 50
rect 146 42 151 48
rect 153 68 161 70
rect 153 66 156 68
rect 158 66 161 68
rect 153 42 161 66
rect 163 55 168 70
rect 163 53 170 55
rect 163 51 166 53
rect 168 51 170 53
rect 163 46 170 51
rect 163 44 166 46
rect 168 44 170 46
rect 163 42 170 44
<< alu1 >>
rect -2 81 186 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 186 81
rect -2 68 186 79
rect 2 61 48 62
rect 2 59 4 61
rect 6 59 24 61
rect 26 59 44 61
rect 46 59 48 61
rect 2 58 48 59
rect 2 54 6 58
rect 2 52 4 54
rect 2 30 6 52
rect 57 37 87 38
rect 57 35 63 37
rect 65 35 87 37
rect 57 34 87 35
rect 2 26 24 30
rect 20 24 21 26
rect 23 24 24 26
rect 81 32 87 34
rect 81 30 91 32
rect 81 28 88 30
rect 90 28 91 30
rect 81 26 91 28
rect 20 22 24 24
rect 20 20 64 22
rect 20 18 60 20
rect 62 18 64 20
rect 58 17 64 18
rect 129 42 142 46
rect 138 37 142 42
rect 154 39 158 55
rect 138 35 139 37
rect 141 35 142 37
rect 138 33 142 35
rect 146 37 162 39
rect 146 35 159 37
rect 161 35 162 37
rect 146 33 162 35
rect 154 25 158 33
rect -2 11 186 12
rect -2 9 39 11
rect 41 9 101 11
rect 103 9 152 11
rect 154 9 186 11
rect -2 1 186 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 186 1
rect -2 -2 186 -1
<< ptie >>
rect 0 1 184 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 184 1
rect 0 -3 184 -1
<< ntie >>
rect 0 81 184 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 184 81
rect 0 77 184 79
<< nmos >>
rect 9 16 11 28
rect 16 16 18 28
rect 26 16 28 28
rect 33 16 35 28
rect 45 16 47 30
rect 55 16 57 30
rect 65 16 67 30
rect 75 16 77 30
rect 85 10 87 22
rect 95 10 97 22
rect 114 16 116 30
rect 124 16 126 30
rect 146 19 148 30
rect 158 16 160 27
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 63 44 65 70
rect 73 44 75 70
rect 83 42 85 70
rect 93 42 95 70
rect 116 42 118 70
rect 123 42 125 70
rect 133 42 135 70
rect 151 42 153 70
rect 161 42 163 70
<< polyct0 >>
rect 50 51 52 53
rect 18 35 20 37
rect 104 35 106 37
rect 114 35 116 37
rect 135 18 137 20
<< polyct1 >>
rect 63 35 65 37
rect 139 35 141 37
rect 159 35 161 37
rect 88 28 90 30
<< ndifct0 >>
rect 4 18 6 20
rect 50 26 52 28
rect 70 26 72 28
rect 70 19 72 21
rect 80 18 82 20
rect 90 18 92 20
rect 109 19 111 21
rect 119 26 121 28
rect 129 26 131 28
rect 141 26 143 28
rect 163 18 165 20
<< ndifct1 >>
rect 21 24 23 26
rect 60 18 62 20
rect 39 9 41 11
rect 101 9 103 11
rect 152 9 154 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
rect 171 79 173 81
rect 179 79 181 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
rect 171 -1 173 1
rect 179 -1 181 1
<< pdifct0 >>
rect 14 51 16 53
rect 14 44 16 46
rect 34 44 36 46
rect 58 66 60 68
rect 58 59 60 61
rect 68 59 70 61
rect 68 52 70 54
rect 78 66 80 68
rect 88 46 90 48
rect 98 66 100 68
rect 106 66 108 68
rect 106 59 108 61
rect 128 60 130 62
rect 138 60 140 62
rect 146 50 148 52
rect 156 66 158 68
rect 166 51 168 53
rect 166 44 168 46
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
rect 24 59 26 61
rect 44 59 46 61
<< alu0 >>
rect 56 66 58 68
rect 60 66 62 68
rect 56 61 62 66
rect 77 66 78 68
rect 80 66 81 68
rect 77 64 81 66
rect 97 66 98 68
rect 100 66 101 68
rect 97 64 101 66
rect 105 66 106 68
rect 108 66 109 68
rect 56 59 58 61
rect 60 59 62 61
rect 56 58 62 59
rect 67 61 71 63
rect 67 59 68 61
rect 70 59 71 61
rect 67 58 71 59
rect 105 61 109 66
rect 154 66 156 68
rect 158 66 160 68
rect 154 65 160 66
rect 105 59 106 61
rect 108 59 109 61
rect 6 50 7 58
rect 67 54 99 58
rect 105 57 109 59
rect 113 62 132 63
rect 113 60 128 62
rect 130 60 132 62
rect 113 59 132 60
rect 136 62 142 63
rect 136 60 138 62
rect 140 60 169 62
rect 12 53 68 54
rect 12 51 14 53
rect 16 51 50 53
rect 52 52 68 53
rect 70 52 71 54
rect 52 51 71 52
rect 12 50 71 51
rect 12 46 17 50
rect 87 48 91 50
rect 12 44 14 46
rect 16 44 17 46
rect 12 42 17 44
rect 32 46 38 47
rect 87 46 88 48
rect 90 46 91 48
rect 32 44 34 46
rect 36 44 38 46
rect 32 38 38 44
rect 48 42 91 46
rect 48 38 52 42
rect 16 37 52 38
rect 16 35 18 37
rect 20 35 52 37
rect 16 34 52 35
rect 48 29 52 34
rect 48 28 74 29
rect 48 26 50 28
rect 52 26 70 28
rect 72 26 74 28
rect 48 25 74 26
rect 3 20 7 22
rect 3 18 4 20
rect 6 18 7 20
rect 3 12 7 18
rect 69 21 74 25
rect 95 21 99 54
rect 113 53 117 59
rect 136 58 169 60
rect 103 49 117 53
rect 121 52 150 53
rect 121 50 146 52
rect 148 50 150 52
rect 121 49 150 50
rect 103 37 107 49
rect 121 38 125 49
rect 103 35 104 37
rect 106 35 107 37
rect 103 29 107 35
rect 112 37 131 38
rect 112 35 114 37
rect 116 35 131 37
rect 112 34 131 35
rect 127 29 131 34
rect 165 53 169 58
rect 165 51 166 53
rect 168 51 169 53
rect 165 46 169 51
rect 165 44 166 46
rect 168 44 169 46
rect 103 28 123 29
rect 103 26 119 28
rect 121 26 123 28
rect 103 25 123 26
rect 127 28 145 29
rect 127 26 129 28
rect 131 26 141 28
rect 143 26 145 28
rect 127 25 145 26
rect 69 19 70 21
rect 72 19 74 21
rect 69 17 74 19
rect 78 20 84 21
rect 78 18 80 20
rect 82 18 84 20
rect 78 12 84 18
rect 88 20 99 21
rect 88 18 90 20
rect 92 18 99 20
rect 88 17 99 18
rect 107 21 113 22
rect 165 21 169 44
rect 107 19 109 21
rect 111 20 169 21
rect 111 19 135 20
rect 107 18 135 19
rect 137 18 163 20
rect 165 18 169 20
rect 107 17 169 18
<< labels >>
rlabel alu0 14 48 14 48 6 cn
rlabel alu0 35 40 35 40 6 zn
rlabel alu0 41 52 41 52 6 cn
rlabel alu0 61 27 61 27 6 zn
rlabel alu0 71 23 71 23 6 zn
rlabel alu0 93 19 93 19 6 cn
rlabel alu0 69 44 69 44 6 zn
rlabel alu0 105 39 105 39 6 iz
rlabel alu0 83 56 83 56 6 cn
rlabel alu0 113 27 113 27 6 iz
rlabel alu0 136 27 136 27 6 bn
rlabel alu0 123 43 123 43 6 bn
rlabel alu0 122 61 122 61 6 iz
rlabel alu0 138 19 138 19 6 an
rlabel alu0 135 51 135 51 6 bn
rlabel alu0 167 39 167 39 6 an
rlabel alu0 152 60 152 60 6 an
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 20 28 20 28 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 44 20 44 20 6 z
rlabel alu1 76 36 76 36 6 c
rlabel alu1 84 32 84 32 6 c
rlabel alu1 68 36 68 36 6 c
rlabel alu1 60 36 60 36 6 c
rlabel alu1 44 60 44 60 6 z
rlabel alu1 92 6 92 6 6 vss
rlabel alu1 132 44 132 44 6 b
rlabel alu1 92 74 92 74 6 vdd
rlabel polyct1 140 36 140 36 6 b
rlabel alu1 148 36 148 36 6 a
rlabel alu1 156 28 156 28 6 a
rlabel alu1 156 40 156 40 6 a
<< end >>
