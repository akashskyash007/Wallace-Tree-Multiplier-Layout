magic
tech scmos
timestamp 1199202516
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 63 11 68
rect 22 63 24 68
rect 32 63 34 68
rect 44 61 46 65
rect 9 37 11 51
rect 22 47 24 51
rect 16 45 24 47
rect 16 43 18 45
rect 20 43 24 45
rect 16 41 24 43
rect 9 35 15 37
rect 9 33 11 35
rect 13 33 15 35
rect 9 31 15 33
rect 22 31 24 41
rect 32 40 34 51
rect 44 46 46 49
rect 41 44 47 46
rect 41 42 43 44
rect 45 42 47 44
rect 41 40 47 42
rect 32 38 37 40
rect 35 36 37 38
rect 35 34 41 36
rect 35 32 37 34
rect 39 32 41 34
rect 9 26 11 31
rect 22 29 30 31
rect 28 26 30 29
rect 35 30 41 32
rect 35 26 37 30
rect 45 26 47 40
rect 9 15 11 20
rect 28 11 30 16
rect 35 11 37 16
rect 45 15 47 20
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 11 20 17 26
rect 23 24 28 26
rect 13 14 17 20
rect 21 22 28 24
rect 21 20 23 22
rect 25 20 28 22
rect 21 18 28 20
rect 23 16 28 18
rect 30 16 35 26
rect 37 24 45 26
rect 37 22 40 24
rect 42 22 45 24
rect 37 20 45 22
rect 47 24 54 26
rect 47 22 50 24
rect 52 22 54 24
rect 47 20 54 22
rect 37 16 43 20
rect 13 11 19 14
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 4 57 9 63
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 51 9 53
rect 11 61 22 63
rect 11 59 16 61
rect 18 59 22 61
rect 11 51 22 59
rect 24 56 32 63
rect 24 54 27 56
rect 29 54 32 56
rect 24 51 32 54
rect 34 61 42 63
rect 34 59 37 61
rect 39 59 44 61
rect 34 51 44 59
rect 36 49 44 51
rect 46 55 51 61
rect 46 53 53 55
rect 46 51 49 53
rect 51 51 53 53
rect 46 49 53 51
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 26 56 30 63
rect 26 54 27 56
rect 29 54 30 56
rect 10 35 22 39
rect 10 33 11 35
rect 13 33 22 35
rect 10 17 14 33
rect 26 23 30 54
rect 34 47 38 55
rect 34 44 47 47
rect 34 42 43 44
rect 45 42 47 44
rect 34 41 47 42
rect 18 22 30 23
rect 18 20 23 22
rect 25 20 30 22
rect 18 17 30 20
rect -2 11 58 12
rect -2 9 15 11
rect 17 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 20 11 26
rect 28 16 30 26
rect 35 16 37 26
rect 45 20 47 26
<< pmos >>
rect 9 51 11 63
rect 22 51 24 63
rect 32 51 34 63
rect 44 49 46 61
<< polyct0 >>
rect 18 43 20 45
rect 37 32 39 34
<< polyct1 >>
rect 11 33 13 35
rect 43 42 45 44
<< ndifct0 >>
rect 4 22 6 24
rect 40 22 42 24
rect 50 22 52 24
<< ndifct1 >>
rect 23 20 25 22
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 53 6 55
rect 16 59 18 61
rect 37 59 39 61
rect 49 51 51 53
<< pdifct1 >>
rect 27 54 29 56
<< alu0 >>
rect 15 61 19 68
rect 15 59 16 61
rect 18 59 19 61
rect 15 57 19 59
rect 3 55 7 57
rect 3 53 4 55
rect 6 53 7 55
rect 3 46 7 53
rect 35 61 41 68
rect 35 59 37 61
rect 39 59 41 61
rect 35 58 41 59
rect 2 45 22 46
rect 2 43 18 45
rect 20 43 22 45
rect 2 42 22 43
rect 2 26 6 42
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 20 7 22
rect 47 53 54 54
rect 47 51 49 53
rect 51 51 54 53
rect 47 50 54 51
rect 50 35 54 50
rect 35 34 54 35
rect 35 32 37 34
rect 39 32 54 34
rect 35 31 54 32
rect 50 26 54 31
rect 39 24 43 26
rect 39 22 40 24
rect 42 22 43 24
rect 39 12 43 22
rect 49 24 54 26
rect 49 22 50 24
rect 52 22 54 24
rect 49 20 54 22
<< labels >>
rlabel alu0 5 49 5 49 6 bn
rlabel alu0 4 33 4 33 6 bn
rlabel alu0 12 44 12 44 6 bn
rlabel alu0 44 33 44 33 6 an
rlabel alu0 52 37 52 37 6 an
rlabel pdifct0 50 52 50 52 6 an
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 28 12 28 6 b
rlabel alu1 20 36 20 36 6 b
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 48 36 48 6 a
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 44 44 44 6 a
<< end >>
