magic
tech scmos
timestamp 1199203135
<< ab >>
rect 0 0 152 80
<< nwell >>
rect -5 36 157 88
<< pwell >>
rect -5 -8 157 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 46 70 48 74
rect 56 70 58 74
rect 63 70 65 74
rect 73 70 75 74
rect 80 70 82 74
rect 90 70 92 74
rect 97 70 99 74
rect 107 70 109 74
rect 114 70 116 74
rect 124 62 126 67
rect 131 62 133 67
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 46 39 48 42
rect 56 39 58 42
rect 9 37 31 39
rect 9 30 11 37
rect 18 35 20 37
rect 22 35 27 37
rect 29 35 31 37
rect 18 33 31 35
rect 36 37 42 39
rect 46 37 58 39
rect 63 39 65 42
rect 73 39 75 42
rect 63 37 75 39
rect 80 39 82 42
rect 90 39 92 42
rect 80 37 92 39
rect 97 39 99 42
rect 107 39 109 42
rect 114 39 116 42
rect 124 39 126 42
rect 131 39 133 42
rect 97 37 109 39
rect 36 35 38 37
rect 40 35 42 37
rect 36 33 42 35
rect 19 30 21 33
rect 29 30 31 33
rect 40 24 42 29
rect 50 28 52 37
rect 66 35 68 37
rect 70 35 72 37
rect 66 33 72 35
rect 80 35 82 37
rect 84 35 86 37
rect 80 33 86 35
rect 97 35 105 37
rect 107 35 109 37
rect 97 33 109 35
rect 113 37 126 39
rect 130 37 136 39
rect 113 35 115 37
rect 117 35 119 37
rect 113 33 119 35
rect 130 35 132 37
rect 134 35 136 37
rect 130 33 142 35
rect 60 28 62 33
rect 70 30 72 33
rect 83 30 85 33
rect 93 31 105 33
rect 70 12 72 16
rect 93 28 95 31
rect 103 28 105 31
rect 113 30 115 33
rect 130 30 132 33
rect 140 30 142 33
rect 9 6 11 11
rect 19 6 21 11
rect 29 8 31 11
rect 40 8 42 11
rect 29 6 42 8
rect 50 8 52 11
rect 60 8 62 11
rect 83 8 85 14
rect 130 15 132 20
rect 140 15 142 20
rect 50 6 85 8
rect 93 6 95 10
rect 103 6 105 10
rect 113 6 115 10
<< ndif >>
rect 4 22 9 30
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 4 11 9 16
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 11 19 26
rect 21 20 29 30
rect 21 18 24 20
rect 26 18 29 20
rect 21 11 29 18
rect 31 28 38 30
rect 31 26 34 28
rect 36 26 38 28
rect 31 24 38 26
rect 65 28 70 30
rect 45 24 50 28
rect 31 11 40 24
rect 42 22 50 24
rect 42 20 45 22
rect 47 20 50 22
rect 42 11 50 20
rect 52 15 60 28
rect 52 13 55 15
rect 57 13 60 15
rect 52 11 60 13
rect 62 25 70 28
rect 62 23 65 25
rect 67 23 70 25
rect 62 16 70 23
rect 72 20 83 30
rect 72 18 77 20
rect 79 18 83 20
rect 72 16 83 18
rect 62 11 67 16
rect 78 14 83 16
rect 85 28 90 30
rect 108 28 113 30
rect 85 25 93 28
rect 85 23 88 25
rect 90 23 93 25
rect 85 14 93 23
rect 88 10 93 14
rect 95 14 103 28
rect 95 12 98 14
rect 100 12 103 14
rect 95 10 103 12
rect 105 21 113 28
rect 105 19 108 21
rect 110 19 113 21
rect 105 10 113 19
rect 115 20 130 30
rect 132 25 140 30
rect 132 23 135 25
rect 137 23 140 25
rect 132 20 140 23
rect 142 24 149 30
rect 142 22 145 24
rect 147 22 149 24
rect 142 20 149 22
rect 115 14 128 20
rect 115 12 122 14
rect 124 12 128 14
rect 115 10 128 12
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 42 19 59
rect 21 60 29 70
rect 21 58 24 60
rect 26 58 29 60
rect 21 53 29 58
rect 21 51 24 53
rect 26 51 29 53
rect 21 42 29 51
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 42 39 59
rect 41 42 46 70
rect 48 60 56 70
rect 48 58 51 60
rect 53 58 56 60
rect 48 53 56 58
rect 48 51 51 53
rect 53 51 56 53
rect 48 42 56 51
rect 58 42 63 70
rect 65 68 73 70
rect 65 66 68 68
rect 70 66 73 68
rect 65 61 73 66
rect 65 59 68 61
rect 70 59 73 61
rect 65 42 73 59
rect 75 42 80 70
rect 82 60 90 70
rect 82 58 85 60
rect 87 58 90 60
rect 82 53 90 58
rect 82 51 85 53
rect 87 51 90 53
rect 82 42 90 51
rect 92 42 97 70
rect 99 68 107 70
rect 99 66 102 68
rect 104 66 107 68
rect 99 61 107 66
rect 99 59 102 61
rect 104 59 107 61
rect 99 42 107 59
rect 109 42 114 70
rect 116 62 121 70
rect 116 60 124 62
rect 116 58 119 60
rect 121 58 124 60
rect 116 53 124 58
rect 116 51 119 53
rect 121 51 124 53
rect 116 42 124 51
rect 126 42 131 62
rect 133 60 140 62
rect 133 58 136 60
rect 138 58 140 60
rect 133 53 140 58
rect 133 51 136 53
rect 138 51 140 53
rect 133 42 140 51
<< alu1 >>
rect -2 81 154 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 154 81
rect -2 68 154 79
rect 50 60 54 63
rect 50 58 51 60
rect 53 58 54 60
rect 82 60 88 63
rect 82 58 85 60
rect 87 58 88 60
rect 50 54 54 58
rect 82 54 88 58
rect 2 53 127 54
rect 2 51 4 53
rect 6 51 24 53
rect 26 51 51 53
rect 53 51 85 53
rect 87 51 119 53
rect 121 51 127 53
rect 2 50 127 51
rect 2 46 6 50
rect 2 44 4 46
rect 2 30 6 44
rect 25 42 39 46
rect 68 42 135 46
rect 25 38 31 42
rect 68 38 72 42
rect 17 37 31 38
rect 17 35 20 37
rect 22 35 27 37
rect 29 35 31 37
rect 17 34 31 35
rect 36 37 72 38
rect 36 35 38 37
rect 40 35 68 37
rect 70 35 72 37
rect 36 34 72 35
rect 80 37 99 38
rect 80 35 82 37
rect 84 35 99 37
rect 80 34 99 35
rect 113 37 119 38
rect 113 35 115 37
rect 117 35 119 37
rect 95 30 99 34
rect 113 30 119 35
rect 130 37 135 42
rect 130 35 132 37
rect 134 35 135 37
rect 130 33 135 35
rect 2 28 39 30
rect 2 26 14 28
rect 16 26 34 28
rect 36 26 39 28
rect 2 25 39 26
rect 95 26 119 30
rect -2 1 154 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 154 1
rect -2 -2 154 -1
<< ptie >>
rect 0 1 152 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 152 1
rect 0 -3 152 -1
<< ntie >>
rect 0 81 152 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 152 81
rect 0 77 152 79
<< nmos >>
rect 9 11 11 30
rect 19 11 21 30
rect 29 11 31 30
rect 40 11 42 24
rect 50 11 52 28
rect 60 11 62 28
rect 70 16 72 30
rect 83 14 85 30
rect 93 10 95 28
rect 103 10 105 28
rect 113 10 115 30
rect 130 20 132 30
rect 140 20 142 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 46 42 48 70
rect 56 42 58 70
rect 63 42 65 70
rect 73 42 75 70
rect 80 42 82 70
rect 90 42 92 70
rect 97 42 99 70
rect 107 42 109 70
rect 114 42 116 70
rect 124 42 126 62
rect 131 42 133 62
<< polyct0 >>
rect 105 35 107 37
<< polyct1 >>
rect 20 35 22 37
rect 27 35 29 37
rect 38 35 40 37
rect 68 35 70 37
rect 82 35 84 37
rect 115 35 117 37
rect 132 35 134 37
<< ndifct0 >>
rect 4 18 6 20
rect 24 18 26 20
rect 45 20 47 22
rect 55 13 57 15
rect 65 23 67 25
rect 77 18 79 20
rect 88 23 90 25
rect 98 12 100 14
rect 108 19 110 21
rect 135 23 137 25
rect 145 22 147 24
rect 122 12 124 14
<< ndifct1 >>
rect 14 26 16 28
rect 34 26 36 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
<< pdifct0 >>
rect 14 66 16 68
rect 14 59 16 61
rect 24 58 26 60
rect 34 66 36 68
rect 34 59 36 61
rect 68 66 70 68
rect 68 59 70 61
rect 102 66 104 68
rect 102 59 104 61
rect 119 58 121 60
rect 136 58 138 60
rect 136 51 138 53
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 51 26 53
rect 51 58 53 60
rect 51 51 53 53
rect 85 58 87 60
rect 85 51 87 53
rect 119 51 121 53
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 61 18 66
rect 32 66 34 68
rect 36 66 38 68
rect 12 59 14 61
rect 16 59 18 61
rect 12 58 18 59
rect 23 60 27 62
rect 23 58 24 60
rect 26 58 27 60
rect 32 61 38 66
rect 66 66 68 68
rect 70 66 72 68
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 66 61 72 66
rect 100 66 102 68
rect 104 66 106 68
rect 66 59 68 61
rect 70 59 72 61
rect 66 58 72 59
rect 100 61 106 66
rect 100 59 102 61
rect 104 59 106 61
rect 100 58 106 59
rect 118 60 123 62
rect 118 58 119 60
rect 121 58 123 60
rect 23 54 27 58
rect 118 54 123 58
rect 134 60 140 68
rect 134 58 136 60
rect 138 58 140 60
rect 134 53 140 58
rect 134 51 136 53
rect 138 51 140 53
rect 134 50 140 51
rect 6 42 7 50
rect 103 37 109 42
rect 103 35 105 37
rect 107 35 109 37
rect 103 34 109 35
rect 44 25 91 29
rect 44 22 48 25
rect 44 21 45 22
rect 2 20 45 21
rect 47 20 48 22
rect 64 23 65 25
rect 67 23 68 25
rect 64 21 68 23
rect 87 23 88 25
rect 90 23 91 25
rect 87 22 91 23
rect 134 25 138 27
rect 134 23 135 25
rect 137 23 138 25
rect 134 22 138 23
rect 87 21 138 22
rect 2 18 4 20
rect 6 18 24 20
rect 26 18 48 20
rect 2 17 48 18
rect 75 20 81 21
rect 75 18 77 20
rect 79 18 81 20
rect 87 19 108 21
rect 110 19 138 21
rect 87 18 138 19
rect 144 24 148 26
rect 144 22 145 24
rect 147 22 148 24
rect 54 15 58 17
rect 54 13 55 15
rect 57 13 58 15
rect 54 12 58 13
rect 75 12 81 18
rect 96 14 102 15
rect 96 12 98 14
rect 100 12 102 14
rect 120 14 126 15
rect 120 12 122 14
rect 124 12 126 14
rect 144 12 148 22
<< labels >>
rlabel ndifct0 25 19 25 19 6 n1
rlabel alu0 89 23 89 23 6 n1
rlabel alu0 67 27 67 27 6 n1
rlabel alu0 112 20 112 20 6 n1
rlabel alu0 136 22 136 22 6 n1
rlabel alu1 20 28 20 28 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 20 36 20 36 6 b
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 28 28 28 6 z
rlabel alu1 36 28 36 28 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 52 36 52 36 6 a1
rlabel alu1 44 36 44 36 6 a1
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 52 44 52 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 52 56 52 56 6 z
rlabel alu1 76 6 76 6 6 vss
rlabel alu1 60 36 60 36 6 a1
rlabel alu1 84 44 84 44 6 a1
rlabel alu1 84 36 84 36 6 a2
rlabel alu1 76 44 76 44 6 a1
rlabel alu1 68 36 68 36 6 a1
rlabel alu1 76 52 76 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 84 56 84 56 6 z
rlabel alu1 76 74 76 74 6 vdd
rlabel alu1 108 28 108 28 6 a2
rlabel alu1 100 28 100 28 6 a2
rlabel alu1 116 32 116 32 6 a2
rlabel alu1 92 44 92 44 6 a1
rlabel alu1 92 36 92 36 6 a2
rlabel alu1 116 44 116 44 6 a1
rlabel alu1 108 44 108 44 6 a1
rlabel alu1 100 44 100 44 6 a1
rlabel alu1 116 52 116 52 6 z
rlabel alu1 108 52 108 52 6 z
rlabel alu1 100 52 100 52 6 z
rlabel alu1 92 52 92 52 6 z
rlabel alu1 124 44 124 44 6 a1
rlabel alu1 132 40 132 40 6 a1
rlabel alu1 124 52 124 52 6 z
<< end >>
