magic
tech scmos
timestamp 1199203174
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 23 70 25 74
rect 30 70 32 74
rect 37 70 39 74
rect 13 61 15 66
rect 13 39 15 50
rect 23 40 25 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 38 26 40
rect 19 36 22 38
rect 24 36 26 38
rect 19 34 26 36
rect 9 23 11 33
rect 19 23 21 34
rect 30 32 32 43
rect 37 40 39 43
rect 37 38 47 40
rect 41 36 43 38
rect 45 36 47 38
rect 41 34 47 36
rect 30 30 37 32
rect 30 28 33 30
rect 35 28 37 30
rect 30 26 37 28
rect 31 23 33 26
rect 41 23 43 34
rect 9 9 11 14
rect 19 9 21 14
rect 31 9 33 14
rect 41 9 43 14
<< ndif >>
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 14 9 17
rect 11 20 19 23
rect 11 18 14 20
rect 16 18 19 20
rect 11 14 19 18
rect 21 14 31 23
rect 33 20 41 23
rect 33 18 36 20
rect 38 18 41 20
rect 33 14 41 18
rect 43 18 50 23
rect 43 16 46 18
rect 48 16 50 18
rect 43 14 50 16
rect 23 11 29 14
rect 23 9 25 11
rect 27 9 29 11
rect 23 7 29 9
<< pdif >>
rect 5 61 11 63
rect 18 61 23 70
rect 5 59 7 61
rect 9 59 13 61
rect 5 50 13 59
rect 15 54 23 61
rect 15 52 18 54
rect 20 52 23 54
rect 15 50 23 52
rect 18 43 23 50
rect 25 43 30 70
rect 32 43 37 70
rect 39 68 48 70
rect 39 66 43 68
rect 45 66 48 68
rect 39 61 48 66
rect 39 59 43 61
rect 45 59 48 61
rect 39 43 48 59
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 54 22 55
rect 2 52 18 54
rect 20 52 22 54
rect 2 51 22 52
rect 2 49 14 51
rect 2 21 6 49
rect 26 47 30 63
rect 34 49 47 55
rect 18 41 30 47
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 34 30 38 39
rect 42 38 47 49
rect 42 36 43 38
rect 45 36 47 38
rect 42 34 47 36
rect 10 26 23 30
rect 35 28 47 30
rect 34 25 47 28
rect 2 19 4 21
rect 2 17 6 19
rect -2 11 58 12
rect -2 9 25 11
rect 27 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 14 11 23
rect 19 14 21 23
rect 31 14 33 23
rect 41 14 43 23
<< pmos >>
rect 13 50 15 61
rect 23 43 25 70
rect 30 43 32 70
rect 37 43 39 70
<< polyct0 >>
rect 22 36 24 38
rect 33 28 34 30
<< polyct1 >>
rect 11 35 13 37
rect 43 36 45 38
rect 34 28 35 30
<< ndifct0 >>
rect 14 18 16 20
rect 36 18 38 20
rect 46 16 48 18
<< ndifct1 >>
rect 4 19 6 21
rect 25 9 27 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 7 59 9 61
rect 43 66 45 68
rect 43 59 45 61
<< pdifct1 >>
rect 18 52 20 54
<< alu0 >>
rect 5 61 11 68
rect 41 66 43 68
rect 45 66 47 68
rect 5 59 7 61
rect 9 59 11 61
rect 5 58 11 59
rect 41 61 47 66
rect 41 59 43 61
rect 45 59 47 61
rect 41 58 47 59
rect 20 38 26 41
rect 20 36 22 38
rect 24 36 26 38
rect 20 35 26 36
rect 32 30 34 32
rect 32 28 33 30
rect 32 26 34 28
rect 6 17 7 23
rect 12 20 40 21
rect 12 18 14 20
rect 16 18 36 20
rect 38 18 40 20
rect 12 17 40 18
rect 45 18 49 20
rect 45 16 46 18
rect 48 16 49 18
rect 45 12 49 16
<< labels >>
rlabel alu0 26 19 26 19 6 n3
rlabel alu1 4 36 4 36 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 44 20 44 6 a3
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 32 36 32 6 a2
rlabel alu1 28 52 28 52 6 a3
rlabel alu1 36 52 36 52 6 a1
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 44 48 44 48 6 a1
<< end >>
