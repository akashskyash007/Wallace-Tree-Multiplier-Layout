magic
tech scmos
timestamp 1199202922
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 50 66 52 70
rect 60 66 62 70
rect 67 66 69 70
rect 9 29 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 16 33 28 35
rect 33 35 35 38
rect 43 35 45 38
rect 33 33 45 35
rect 50 35 52 38
rect 60 35 62 38
rect 50 33 62 35
rect 22 31 24 33
rect 26 31 28 33
rect 22 29 28 31
rect 35 31 41 33
rect 35 29 37 31
rect 39 29 41 31
rect 50 31 52 33
rect 54 31 56 33
rect 50 29 56 31
rect 9 27 18 29
rect 12 25 14 27
rect 16 25 18 27
rect 12 23 18 25
rect 13 20 15 23
rect 23 20 25 29
rect 35 27 41 29
rect 45 27 56 29
rect 67 27 69 38
rect 35 24 37 27
rect 45 24 47 27
rect 63 25 69 27
rect 63 23 65 25
rect 67 23 69 25
rect 63 21 69 23
rect 13 2 15 7
rect 23 2 25 7
rect 35 2 37 7
rect 45 2 47 7
<< ndif >>
rect 27 20 35 24
rect 4 7 13 20
rect 15 17 23 20
rect 15 15 18 17
rect 20 15 23 17
rect 15 7 23 15
rect 25 7 35 20
rect 37 17 45 24
rect 37 15 40 17
rect 42 15 45 17
rect 37 7 45 15
rect 47 18 55 24
rect 47 16 50 18
rect 52 16 55 18
rect 47 11 55 16
rect 47 9 50 11
rect 52 9 55 11
rect 47 7 55 9
rect 4 5 7 7
rect 9 5 11 7
rect 4 3 11 5
rect 27 5 29 7
rect 31 5 33 7
rect 27 3 33 5
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 38 16 66
rect 18 49 26 66
rect 18 47 21 49
rect 23 47 26 49
rect 18 42 26 47
rect 18 40 21 42
rect 23 40 26 42
rect 18 38 26 40
rect 28 38 33 66
rect 35 64 43 66
rect 35 62 38 64
rect 40 62 43 64
rect 35 57 43 62
rect 35 55 38 57
rect 40 55 43 57
rect 35 38 43 55
rect 45 38 50 66
rect 52 49 60 66
rect 52 47 55 49
rect 57 47 60 49
rect 52 42 60 47
rect 52 40 55 42
rect 57 40 60 42
rect 52 38 60 40
rect 62 38 67 66
rect 69 64 77 66
rect 69 62 72 64
rect 74 62 77 64
rect 69 57 77 62
rect 69 55 72 57
rect 74 55 77 57
rect 69 38 77 55
<< alu1 >>
rect -2 64 82 72
rect 19 49 59 50
rect 19 47 21 49
rect 23 47 55 49
rect 57 47 59 49
rect 19 46 59 47
rect 19 43 24 46
rect 2 42 24 43
rect 54 42 59 46
rect 2 40 21 42
rect 23 40 24 42
rect 2 38 24 40
rect 28 38 50 42
rect 54 40 55 42
rect 57 40 63 42
rect 54 38 63 40
rect 2 18 6 38
rect 28 34 32 38
rect 22 33 32 34
rect 46 34 50 38
rect 46 33 63 34
rect 22 31 24 33
rect 26 31 32 33
rect 22 30 32 31
rect 36 31 40 33
rect 36 29 37 31
rect 39 29 40 31
rect 46 31 52 33
rect 54 31 63 33
rect 46 30 63 31
rect 13 27 17 29
rect 13 25 14 27
rect 16 26 17 27
rect 36 26 40 29
rect 16 25 70 26
rect 13 23 65 25
rect 67 23 70 25
rect 13 22 70 23
rect 2 17 44 18
rect 2 15 18 17
rect 20 15 40 17
rect 42 15 44 17
rect 2 14 44 15
rect 66 13 70 22
rect -2 7 82 8
rect -2 5 7 7
rect 9 5 29 7
rect 31 5 63 7
rect 65 5 71 7
rect 73 5 82 7
rect -2 0 82 5
<< ptie >>
rect 61 7 75 18
rect 61 5 63 7
rect 65 5 71 7
rect 73 5 75 7
rect 61 3 75 5
<< nmos >>
rect 13 7 15 20
rect 23 7 25 20
rect 35 7 37 24
rect 45 7 47 24
<< pmos >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 38 45 66
rect 50 38 52 66
rect 60 38 62 66
rect 67 38 69 66
<< polyct1 >>
rect 24 31 26 33
rect 37 29 39 31
rect 52 31 54 33
rect 14 25 16 27
rect 65 23 67 25
<< ndifct0 >>
rect 50 16 52 18
rect 50 9 52 11
<< ndifct1 >>
rect 18 15 20 17
rect 40 15 42 17
rect 7 5 9 7
rect 29 5 31 7
<< ptiect1 >>
rect 63 5 65 7
rect 71 5 73 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 38 62 40 64
rect 38 55 40 57
rect 72 62 74 64
rect 72 55 74 57
<< pdifct1 >>
rect 21 47 23 49
rect 21 40 23 42
rect 55 47 57 49
rect 55 40 57 42
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 36 62 38 64
rect 40 62 42 64
rect 36 57 42 62
rect 36 55 38 57
rect 40 55 42 57
rect 36 54 42 55
rect 70 62 72 64
rect 74 62 76 64
rect 70 57 76 62
rect 70 55 72 57
rect 74 55 76 57
rect 70 54 76 55
rect 48 18 54 19
rect 48 16 50 18
rect 52 16 54 18
rect 48 11 54 16
rect 48 9 50 11
rect 52 9 54 11
rect 48 8 54 9
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 24 20 24 6 a
rlabel alu1 28 24 28 24 6 a
rlabel alu1 28 32 28 32 6 b
rlabel alu1 12 40 12 40 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 36 16 36 16 6 z
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 52 24 52 24 6 a
rlabel alu1 60 24 60 24 6 a
rlabel alu1 60 32 60 32 6 b
rlabel alu1 52 32 52 32 6 b
rlabel alu1 60 40 60 40 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 68 16 68 16 6 a
<< end >>
