magic
tech scmos
timestamp 1199202429
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 13 60 15 65
rect 13 39 15 45
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 29 11 33
rect 9 17 11 22
<< ndif >>
rect 2 27 9 29
rect 2 25 4 27
rect 6 25 9 27
rect 2 22 9 25
rect 11 22 19 29
rect 13 21 19 22
rect 13 19 15 21
rect 17 19 19 21
rect 13 17 19 19
<< pdif >>
rect 5 61 11 63
rect 5 59 7 61
rect 9 60 11 61
rect 9 59 13 60
rect 5 45 13 59
rect 15 55 20 60
rect 15 53 22 55
rect 15 51 18 53
rect 20 51 22 53
rect 15 49 22 51
rect 15 45 20 49
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 68 26 79
rect 2 53 22 54
rect 2 51 18 53
rect 20 51 22 53
rect 2 50 22 51
rect 2 29 6 50
rect 10 37 22 39
rect 10 35 11 37
rect 13 35 22 37
rect 10 33 22 35
rect 2 27 7 29
rect 2 25 4 27
rect 6 25 7 27
rect 18 25 22 33
rect 2 23 7 25
rect -2 1 26 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 22 11 29
<< pmos >>
rect 13 45 15 60
<< polyct1 >>
rect 11 35 13 37
<< ndifct0 >>
rect 15 19 17 21
<< ndifct1 >>
rect 4 25 6 27
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct0 >>
rect 7 59 9 61
<< pdifct1 >>
rect 18 51 20 53
<< alu0 >>
rect 5 61 11 68
rect 5 59 7 61
rect 9 59 11 61
rect 5 58 11 59
rect 13 21 19 22
rect 13 19 15 21
rect 17 19 19 21
rect 13 12 19 19
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 32 20 32 6 a
<< end >>
