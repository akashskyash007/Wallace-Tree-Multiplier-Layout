magic
tech scmos
timestamp 1199202113
<< ab >>
rect 0 0 152 72
<< nwell >>
rect -5 32 157 77
<< pwell >>
rect -5 -5 157 32
<< poly >>
rect 19 65 21 70
rect 29 65 31 70
rect 39 65 41 70
rect 49 65 51 70
rect 59 65 61 70
rect 71 65 73 70
rect 78 65 80 70
rect 88 65 90 70
rect 95 65 97 70
rect 107 65 109 70
rect 117 65 119 70
rect 127 65 129 70
rect 9 55 11 60
rect 137 55 139 60
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 71 35 73 38
rect 78 35 80 38
rect 88 35 90 38
rect 95 35 97 38
rect 9 33 21 35
rect 9 31 11 33
rect 13 31 21 33
rect 9 29 21 31
rect 25 33 32 35
rect 25 31 27 33
rect 29 31 32 33
rect 25 29 32 31
rect 39 33 52 35
rect 39 31 48 33
rect 50 31 52 33
rect 39 29 52 31
rect 59 33 73 35
rect 59 31 67 33
rect 69 31 73 33
rect 59 29 73 31
rect 77 33 90 35
rect 77 31 86 33
rect 88 31 90 33
rect 77 29 90 31
rect 94 33 102 35
rect 94 31 98 33
rect 100 31 102 33
rect 94 29 102 31
rect 107 29 109 38
rect 117 29 119 38
rect 127 34 129 38
rect 137 34 139 38
rect 9 26 11 29
rect 19 26 21 29
rect 30 26 32 29
rect 40 26 42 29
rect 50 26 52 29
rect 60 26 62 29
rect 70 26 72 29
rect 77 26 79 29
rect 87 26 89 29
rect 94 26 96 29
rect 106 27 119 29
rect 9 11 11 15
rect 19 11 21 15
rect 30 7 32 12
rect 40 7 42 12
rect 50 7 52 12
rect 60 7 62 12
rect 70 11 72 15
rect 77 10 79 15
rect 106 25 115 27
rect 117 25 119 27
rect 106 23 119 25
rect 126 32 139 34
rect 126 30 135 32
rect 137 30 139 32
rect 126 28 139 30
rect 106 20 108 23
rect 116 20 118 23
rect 126 20 128 28
rect 136 20 138 28
rect 87 8 89 13
rect 94 8 96 13
rect 106 2 108 6
rect 116 2 118 6
rect 126 4 128 9
rect 136 4 138 9
<< ndif >>
rect 2 15 9 26
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 15 19 22
rect 21 16 30 26
rect 21 15 25 16
rect 2 9 7 15
rect 23 14 25 15
rect 27 14 30 16
rect 23 12 30 14
rect 32 17 40 26
rect 32 15 35 17
rect 37 15 40 17
rect 32 12 40 15
rect 42 24 50 26
rect 42 22 45 24
rect 47 22 50 24
rect 42 12 50 22
rect 52 17 60 26
rect 52 15 55 17
rect 57 15 60 17
rect 52 12 60 15
rect 62 15 70 26
rect 72 15 77 26
rect 79 24 87 26
rect 79 22 82 24
rect 84 22 87 24
rect 79 15 87 22
rect 62 12 68 15
rect 2 7 8 9
rect 2 5 4 7
rect 6 5 8 7
rect 2 3 8 5
rect 64 9 68 12
rect 82 13 87 15
rect 89 13 94 26
rect 96 20 104 26
rect 96 13 106 20
rect 64 7 70 9
rect 98 10 106 13
rect 98 8 100 10
rect 102 8 106 10
rect 64 5 66 7
rect 68 5 70 7
rect 98 6 106 8
rect 108 17 116 20
rect 108 15 111 17
rect 113 15 116 17
rect 108 6 116 15
rect 118 13 126 20
rect 118 11 121 13
rect 123 11 126 13
rect 118 9 126 11
rect 128 18 136 20
rect 128 16 131 18
rect 133 16 136 18
rect 128 9 136 16
rect 138 13 146 20
rect 138 11 141 13
rect 143 11 146 13
rect 138 9 146 11
rect 118 6 124 9
rect 64 3 70 5
<< pdif >>
rect 99 67 105 69
rect 99 65 101 67
rect 103 65 105 67
rect 14 55 19 65
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 45 9 51
rect 2 43 4 45
rect 6 43 9 45
rect 2 38 9 43
rect 11 49 19 55
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 63 29 65
rect 21 61 24 63
rect 26 61 29 63
rect 21 56 29 61
rect 21 54 24 56
rect 26 54 29 56
rect 21 38 29 54
rect 31 56 39 65
rect 31 54 34 56
rect 36 54 39 56
rect 31 38 39 54
rect 41 42 49 65
rect 41 40 44 42
rect 46 40 49 42
rect 41 38 49 40
rect 51 56 59 65
rect 51 54 54 56
rect 56 54 59 56
rect 51 38 59 54
rect 61 63 71 65
rect 61 61 65 63
rect 67 61 71 63
rect 61 38 71 61
rect 73 38 78 65
rect 80 42 88 65
rect 80 40 83 42
rect 85 40 88 42
rect 80 38 88 40
rect 90 38 95 65
rect 97 38 107 65
rect 109 56 117 65
rect 109 54 112 56
rect 114 54 117 56
rect 109 49 117 54
rect 109 47 112 49
rect 114 47 117 49
rect 109 38 117 47
rect 119 63 127 65
rect 119 61 122 63
rect 124 61 127 63
rect 119 55 127 61
rect 119 53 122 55
rect 124 53 127 55
rect 119 38 127 53
rect 129 55 134 65
rect 129 50 137 55
rect 129 48 132 50
rect 134 48 137 50
rect 129 43 137 48
rect 129 41 132 43
rect 134 41 137 43
rect 129 38 137 41
rect 139 53 146 55
rect 139 51 142 53
rect 144 51 146 53
rect 139 45 146 51
rect 139 43 142 45
rect 144 43 146 45
rect 139 38 146 43
<< alu1 >>
rect -2 67 154 72
rect -2 65 5 67
rect 7 65 101 67
rect 103 65 141 67
rect 143 65 154 67
rect -2 64 154 65
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 2 13 6 29
rect 34 42 48 43
rect 34 40 44 42
rect 46 40 48 42
rect 34 38 48 40
rect 34 26 38 38
rect 57 34 63 42
rect 46 33 63 34
rect 46 31 48 33
rect 50 31 63 33
rect 46 30 63 31
rect 74 42 87 43
rect 74 40 83 42
rect 85 40 87 42
rect 74 38 87 40
rect 74 26 78 38
rect 34 24 87 26
rect 34 22 45 24
rect 47 22 82 24
rect 84 22 87 24
rect 74 21 87 22
rect 130 32 142 35
rect 130 30 135 32
rect 137 30 142 32
rect 130 29 142 30
rect 138 21 142 29
rect -2 7 154 8
rect -2 5 4 7
rect 6 5 14 7
rect 16 5 66 7
rect 68 5 154 7
rect -2 0 154 5
<< ptie >>
rect 12 7 18 9
rect 12 5 14 7
rect 16 5 18 7
rect 12 3 18 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 139 67 145 69
rect 139 65 141 67
rect 143 65 145 67
rect 3 63 9 65
rect 139 63 145 65
<< nmos >>
rect 9 15 11 26
rect 19 15 21 26
rect 30 12 32 26
rect 40 12 42 26
rect 50 12 52 26
rect 60 12 62 26
rect 70 15 72 26
rect 77 15 79 26
rect 87 13 89 26
rect 94 13 96 26
rect 106 6 108 20
rect 116 6 118 20
rect 126 9 128 20
rect 136 9 138 20
<< pmos >>
rect 9 38 11 55
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 65
rect 49 38 51 65
rect 59 38 61 65
rect 71 38 73 65
rect 78 38 80 65
rect 88 38 90 65
rect 95 38 97 65
rect 107 38 109 65
rect 117 38 119 65
rect 127 38 129 65
rect 137 38 139 55
<< polyct0 >>
rect 27 31 29 33
rect 67 31 69 33
rect 86 31 88 33
rect 98 31 100 33
rect 115 25 117 27
<< polyct1 >>
rect 11 31 13 33
rect 48 31 50 33
rect 135 30 137 32
<< ndifct0 >>
rect 14 22 16 24
rect 25 14 27 16
rect 35 15 37 17
rect 55 15 57 17
rect 100 8 102 10
rect 111 15 113 17
rect 121 11 123 13
rect 131 16 133 18
rect 141 11 143 13
<< ndifct1 >>
rect 45 22 47 24
rect 82 22 84 24
rect 4 5 6 7
rect 66 5 68 7
<< ntiect1 >>
rect 5 65 7 67
rect 141 65 143 67
<< ptiect1 >>
rect 14 5 16 7
<< pdifct0 >>
rect 4 51 6 53
rect 4 43 6 45
rect 14 47 16 49
rect 14 40 16 42
rect 24 61 26 63
rect 24 54 26 56
rect 34 54 36 56
rect 54 54 56 56
rect 65 61 67 63
rect 112 54 114 56
rect 112 47 114 49
rect 122 61 124 63
rect 122 53 124 55
rect 132 48 134 50
rect 132 41 134 43
rect 142 51 144 53
rect 142 43 144 45
<< pdifct1 >>
rect 101 65 103 67
rect 44 40 46 42
rect 83 40 85 42
<< alu0 >>
rect 3 53 7 64
rect 22 63 28 64
rect 22 61 24 63
rect 26 61 28 63
rect 22 56 28 61
rect 63 63 69 64
rect 63 61 65 63
rect 67 61 69 63
rect 63 60 69 61
rect 121 63 125 64
rect 121 61 122 63
rect 124 61 125 63
rect 22 54 24 56
rect 26 54 28 56
rect 22 53 28 54
rect 32 56 116 57
rect 32 54 34 56
rect 36 54 54 56
rect 56 54 112 56
rect 114 54 116 56
rect 32 53 116 54
rect 3 51 4 53
rect 6 51 7 53
rect 3 45 7 51
rect 3 43 4 45
rect 6 43 7 45
rect 3 41 7 43
rect 12 49 101 50
rect 12 47 14 49
rect 16 47 101 49
rect 12 46 101 47
rect 110 49 116 53
rect 121 55 125 61
rect 121 53 122 55
rect 124 53 125 55
rect 121 51 125 53
rect 141 53 145 64
rect 110 47 112 49
rect 114 47 116 49
rect 110 46 116 47
rect 131 50 135 52
rect 131 48 132 50
rect 134 48 135 50
rect 12 42 18 46
rect 12 40 14 42
rect 16 40 18 42
rect 12 39 18 40
rect 26 33 30 46
rect 26 31 27 33
rect 29 31 30 33
rect 26 25 30 31
rect 12 24 30 25
rect 12 22 14 24
rect 16 22 30 24
rect 66 33 70 46
rect 66 31 67 33
rect 69 31 70 33
rect 66 29 70 31
rect 84 33 94 34
rect 84 31 86 33
rect 88 31 94 33
rect 84 30 94 31
rect 12 21 30 22
rect 43 21 49 22
rect 90 25 94 30
rect 97 33 101 46
rect 131 43 135 48
rect 97 31 98 33
rect 100 31 101 33
rect 97 29 101 31
rect 114 41 132 43
rect 134 41 135 43
rect 141 51 142 53
rect 144 51 145 53
rect 141 45 145 51
rect 141 43 142 45
rect 144 43 145 45
rect 141 41 145 43
rect 114 39 135 41
rect 114 27 118 39
rect 114 25 115 27
rect 117 25 118 27
rect 90 21 134 25
rect 130 18 134 21
rect 33 17 115 18
rect 23 16 29 17
rect 23 14 25 16
rect 27 14 29 16
rect 33 15 35 17
rect 37 15 55 17
rect 57 15 111 17
rect 113 15 115 17
rect 130 16 131 18
rect 133 16 134 18
rect 33 14 115 15
rect 23 8 29 14
rect 120 13 124 15
rect 130 14 134 16
rect 120 11 121 13
rect 123 11 124 13
rect 98 10 104 11
rect 98 8 100 10
rect 102 8 104 10
rect 120 8 124 11
rect 140 13 144 15
rect 140 11 141 13
rect 143 11 144 13
rect 140 8 144 11
<< labels >>
rlabel alu0 21 23 21 23 6 an
rlabel alu0 28 35 28 35 6 an
rlabel alu0 15 44 15 44 6 an
rlabel alu0 68 39 68 39 6 an
rlabel alu0 89 32 89 32 6 bn
rlabel alu0 99 39 99 39 6 an
rlabel alu0 74 16 74 16 6 n3
rlabel alu0 132 19 132 19 6 bn
rlabel alu0 116 32 116 32 6 bn
rlabel alu0 133 45 133 45 6 bn
rlabel alu0 113 51 113 51 6 n1
rlabel alu0 74 55 74 55 6 n1
rlabel alu1 4 24 4 24 6 a
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 68 24 68 24 6 z
rlabel alu1 60 24 60 24 6 z
rlabel alu1 52 32 52 32 6 c
rlabel alu1 52 24 52 24 6 z
rlabel alu1 44 24 44 24 6 z
rlabel alu1 44 40 44 40 6 z
rlabel alu1 60 36 60 36 6 c
rlabel alu1 36 36 36 36 6 z
rlabel alu1 76 4 76 4 6 vss
rlabel alu1 76 32 76 32 6 z
rlabel alu1 84 24 84 24 6 z
rlabel alu1 84 40 84 40 6 z
rlabel alu1 76 68 76 68 6 vdd
rlabel alu1 132 32 132 32 6 b
rlabel alu1 140 28 140 28 6 b
<< end >>
