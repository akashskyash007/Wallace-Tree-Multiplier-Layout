magic
tech scmos
timestamp 1199203139
<< ab >>
rect 0 0 192 72
<< nwell >>
rect -5 32 197 77
<< pwell >>
rect -5 -5 197 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 56 66 58 70
rect 66 66 68 70
rect 73 66 75 70
rect 83 66 85 70
rect 90 66 92 70
rect 100 66 102 70
rect 107 66 109 70
rect 117 66 119 70
rect 124 66 126 70
rect 134 66 136 70
rect 141 66 143 70
rect 151 66 153 70
rect 158 66 160 70
rect 168 59 170 64
rect 175 59 177 64
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 9 33 41 35
rect 9 31 27 33
rect 29 31 31 33
rect 9 29 31 31
rect 9 26 11 29
rect 19 26 21 29
rect 29 26 31 29
rect 39 26 41 33
rect 45 33 51 35
rect 56 35 58 38
rect 66 35 68 38
rect 56 33 68 35
rect 73 35 75 38
rect 83 35 85 38
rect 73 33 85 35
rect 90 35 92 38
rect 100 35 102 38
rect 90 33 102 35
rect 107 35 109 38
rect 117 35 119 38
rect 124 35 126 38
rect 134 35 136 38
rect 107 33 119 35
rect 123 33 136 35
rect 141 35 143 38
rect 151 35 153 38
rect 141 33 153 35
rect 158 35 160 38
rect 168 35 170 38
rect 158 33 170 35
rect 175 35 177 38
rect 175 33 183 35
rect 45 31 47 33
rect 49 31 51 33
rect 45 29 51 31
rect 59 25 61 33
rect 76 31 78 33
rect 80 31 82 33
rect 76 29 82 31
rect 70 25 72 29
rect 80 25 82 29
rect 90 31 92 33
rect 94 31 96 33
rect 90 29 96 31
rect 107 31 112 33
rect 114 31 116 33
rect 107 29 116 31
rect 123 31 129 33
rect 123 29 125 31
rect 127 29 129 31
rect 141 31 143 33
rect 145 31 147 33
rect 141 29 147 31
rect 158 31 162 33
rect 164 31 168 33
rect 158 29 168 31
rect 175 31 179 33
rect 181 31 183 33
rect 175 29 183 31
rect 49 21 51 25
rect 90 24 92 29
rect 100 27 116 29
rect 122 27 129 29
rect 134 27 147 29
rect 156 27 168 29
rect 100 24 102 27
rect 112 24 114 27
rect 122 24 124 27
rect 134 24 136 27
rect 144 24 146 27
rect 156 24 158 27
rect 166 24 168 27
rect 177 26 179 29
rect 80 8 82 12
rect 9 2 11 6
rect 19 2 21 6
rect 29 2 31 6
rect 39 4 41 7
rect 49 4 51 7
rect 39 2 51 4
rect 59 4 61 7
rect 70 4 72 7
rect 90 4 92 12
rect 59 2 92 4
rect 100 2 102 6
rect 112 2 114 6
rect 122 2 124 6
rect 177 11 179 15
rect 134 2 136 6
rect 144 2 146 6
rect 156 4 158 9
rect 166 4 168 9
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 6 9 13
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 6 19 22
rect 21 16 29 26
rect 21 14 24 16
rect 26 14 29 16
rect 21 6 29 14
rect 31 24 39 26
rect 31 22 34 24
rect 36 22 39 24
rect 31 7 39 22
rect 41 21 46 26
rect 54 21 59 25
rect 41 16 49 21
rect 41 14 44 16
rect 46 14 49 16
rect 41 7 49 14
rect 51 19 59 21
rect 51 17 54 19
rect 56 17 59 19
rect 51 7 59 17
rect 61 11 70 25
rect 61 9 65 11
rect 67 9 70 11
rect 61 7 70 9
rect 72 21 80 25
rect 72 19 75 21
rect 77 19 80 21
rect 72 12 80 19
rect 82 24 87 25
rect 170 24 177 26
rect 82 16 90 24
rect 82 14 85 16
rect 87 14 90 16
rect 82 12 90 14
rect 92 21 100 24
rect 92 19 95 21
rect 97 19 100 21
rect 92 12 100 19
rect 72 7 77 12
rect 31 6 36 7
rect 95 6 100 12
rect 102 7 112 24
rect 102 6 106 7
rect 104 5 106 6
rect 108 6 112 7
rect 114 16 122 24
rect 114 14 117 16
rect 119 14 122 16
rect 114 6 122 14
rect 124 7 134 24
rect 124 6 128 7
rect 108 5 110 6
rect 104 3 110 5
rect 126 5 128 6
rect 130 6 134 7
rect 136 16 144 24
rect 136 14 139 16
rect 141 14 144 16
rect 136 6 144 14
rect 146 9 156 24
rect 158 16 166 24
rect 158 14 161 16
rect 163 14 166 16
rect 158 9 166 14
rect 168 15 177 24
rect 179 24 186 26
rect 179 22 182 24
rect 184 22 186 24
rect 179 20 186 22
rect 179 15 184 20
rect 168 13 175 15
rect 168 11 171 13
rect 173 11 175 13
rect 168 9 175 11
rect 146 7 154 9
rect 146 6 150 7
rect 130 5 132 6
rect 126 3 132 5
rect 148 5 150 6
rect 152 5 154 7
rect 148 3 154 5
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 49 39 55
rect 31 47 34 49
rect 36 47 39 49
rect 31 38 39 47
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 38 49 55
rect 51 38 56 66
rect 58 57 66 66
rect 58 55 61 57
rect 63 55 66 57
rect 58 49 66 55
rect 58 47 61 49
rect 63 47 66 49
rect 58 38 66 47
rect 68 38 73 66
rect 75 64 83 66
rect 75 62 78 64
rect 80 62 83 64
rect 75 57 83 62
rect 75 55 78 57
rect 80 55 83 57
rect 75 38 83 55
rect 85 38 90 66
rect 92 56 100 66
rect 92 54 95 56
rect 97 54 100 56
rect 92 49 100 54
rect 92 47 95 49
rect 97 47 100 49
rect 92 38 100 47
rect 102 38 107 66
rect 109 64 117 66
rect 109 62 112 64
rect 114 62 117 64
rect 109 57 117 62
rect 109 55 112 57
rect 114 55 117 57
rect 109 38 117 55
rect 119 38 124 66
rect 126 57 134 66
rect 126 55 129 57
rect 131 55 134 57
rect 126 49 134 55
rect 126 47 129 49
rect 131 47 134 49
rect 126 38 134 47
rect 136 38 141 66
rect 143 64 151 66
rect 143 62 146 64
rect 148 62 151 64
rect 143 57 151 62
rect 143 55 146 57
rect 148 55 151 57
rect 143 38 151 55
rect 153 38 158 66
rect 160 59 165 66
rect 160 57 168 59
rect 160 55 163 57
rect 165 55 168 57
rect 160 50 168 55
rect 160 48 163 50
rect 165 48 168 50
rect 160 38 168 48
rect 170 38 175 59
rect 177 57 185 59
rect 177 55 180 57
rect 182 55 185 57
rect 177 50 185 55
rect 177 48 180 50
rect 182 48 185 50
rect 177 38 185 48
<< alu1 >>
rect -2 67 194 72
rect -2 65 185 67
rect 187 65 194 67
rect -2 64 194 65
rect 33 57 38 59
rect 33 55 34 57
rect 36 55 38 57
rect 33 50 38 55
rect 58 57 64 59
rect 58 55 61 57
rect 63 55 64 57
rect 58 50 64 55
rect 128 57 134 59
rect 128 55 129 57
rect 131 55 134 57
rect 128 50 134 55
rect 162 57 166 59
rect 162 55 163 57
rect 165 55 166 57
rect 162 50 166 55
rect 12 49 163 50
rect 12 47 14 49
rect 16 47 34 49
rect 36 47 61 49
rect 63 47 95 49
rect 97 47 129 49
rect 131 48 163 49
rect 165 48 166 50
rect 131 47 166 48
rect 12 46 166 47
rect 12 43 17 46
rect 2 42 17 43
rect 170 42 174 51
rect 2 40 14 42
rect 16 40 17 42
rect 2 38 17 40
rect 25 38 39 42
rect 78 38 183 42
rect 2 24 6 38
rect 2 22 4 24
rect 2 17 6 22
rect 25 34 31 38
rect 78 34 82 38
rect 17 33 31 34
rect 17 31 27 33
rect 29 31 31 33
rect 17 30 31 31
rect 41 33 82 34
rect 41 31 47 33
rect 49 31 78 33
rect 80 31 82 33
rect 41 30 82 31
rect 89 33 106 34
rect 89 31 92 33
rect 94 31 106 33
rect 89 30 106 31
rect 102 26 106 30
rect 153 33 167 34
rect 153 31 162 33
rect 164 31 167 33
rect 153 30 167 31
rect 177 33 183 38
rect 177 31 179 33
rect 181 31 183 33
rect 177 30 183 31
rect 153 26 159 30
rect 102 22 159 26
rect 2 15 4 17
rect 6 16 48 17
rect 6 15 24 16
rect 2 14 24 15
rect 26 14 44 16
rect 46 14 48 16
rect 2 13 48 14
rect -2 7 194 8
rect -2 5 106 7
rect 108 5 128 7
rect 130 5 150 7
rect 152 5 183 7
rect 185 5 194 7
rect -2 0 194 5
<< ptie >>
rect 179 7 189 9
rect 179 5 183 7
rect 185 5 189 7
rect 179 3 189 5
<< ntie >>
rect 183 67 189 69
rect 183 65 185 67
rect 187 65 189 67
rect 183 63 189 65
<< nmos >>
rect 9 6 11 26
rect 19 6 21 26
rect 29 6 31 26
rect 39 7 41 26
rect 49 7 51 21
rect 59 7 61 25
rect 70 7 72 25
rect 80 12 82 25
rect 90 12 92 24
rect 100 6 102 24
rect 112 6 114 24
rect 122 6 124 24
rect 134 6 136 24
rect 144 6 146 24
rect 156 9 158 24
rect 166 9 168 24
rect 177 15 179 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 56 38 58 66
rect 66 38 68 66
rect 73 38 75 66
rect 83 38 85 66
rect 90 38 92 66
rect 100 38 102 66
rect 107 38 109 66
rect 117 38 119 66
rect 124 38 126 66
rect 134 38 136 66
rect 141 38 143 66
rect 151 38 153 66
rect 158 38 160 66
rect 168 38 170 59
rect 175 38 177 59
<< polyct0 >>
rect 112 31 114 33
rect 125 29 127 31
rect 143 31 145 33
<< polyct1 >>
rect 27 31 29 33
rect 47 31 49 33
rect 78 31 80 33
rect 92 31 94 33
rect 162 31 164 33
rect 179 31 181 33
<< ndifct0 >>
rect 14 22 16 24
rect 34 22 36 24
rect 54 17 56 19
rect 65 9 67 11
rect 75 19 77 21
rect 85 14 87 16
rect 95 19 97 21
rect 117 14 119 16
rect 139 14 141 16
rect 161 14 163 16
rect 182 22 184 24
rect 171 11 173 13
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
rect 24 14 26 16
rect 44 14 46 16
rect 106 5 108 7
rect 128 5 130 7
rect 150 5 152 7
<< ntiect1 >>
rect 185 65 187 67
<< ptiect1 >>
rect 183 5 185 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 24 62 26 64
rect 24 55 26 57
rect 44 62 46 64
rect 44 55 46 57
rect 78 62 80 64
rect 78 55 80 57
rect 95 54 97 56
rect 112 62 114 64
rect 112 55 114 57
rect 146 62 148 64
rect 146 55 148 57
rect 180 55 182 57
rect 180 48 182 50
<< pdifct1 >>
rect 14 47 16 49
rect 14 40 16 42
rect 34 55 36 57
rect 34 47 36 49
rect 61 55 63 57
rect 61 47 63 49
rect 95 47 97 49
rect 129 55 131 57
rect 129 47 131 49
rect 163 55 165 57
rect 163 48 165 50
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 22 62 24 64
rect 26 62 28 64
rect 22 57 28 62
rect 42 62 44 64
rect 46 62 48 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 42 57 48 62
rect 76 62 78 64
rect 80 62 82 64
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 76 57 82 62
rect 110 62 112 64
rect 114 62 116 64
rect 76 55 78 57
rect 80 55 82 57
rect 76 54 82 55
rect 94 56 98 58
rect 94 54 95 56
rect 97 54 98 56
rect 110 57 116 62
rect 144 62 146 64
rect 148 62 150 64
rect 110 55 112 57
rect 114 55 116 57
rect 110 54 116 55
rect 94 50 98 54
rect 144 57 150 62
rect 144 55 146 57
rect 148 55 150 57
rect 144 54 150 55
rect 179 57 183 64
rect 179 55 180 57
rect 182 55 183 57
rect 179 50 183 55
rect 179 48 180 50
rect 182 48 183 50
rect 179 46 183 48
rect 6 17 7 38
rect 110 33 116 38
rect 141 33 147 38
rect 110 31 112 33
rect 114 31 116 33
rect 110 30 116 31
rect 124 31 128 33
rect 124 29 125 31
rect 127 29 128 31
rect 141 31 143 33
rect 145 31 147 33
rect 141 30 147 31
rect 124 26 128 29
rect 12 24 98 25
rect 12 22 14 24
rect 16 22 34 24
rect 36 22 98 24
rect 162 24 186 25
rect 162 22 182 24
rect 184 22 186 24
rect 12 21 98 22
rect 53 19 57 21
rect 53 17 54 19
rect 56 17 57 19
rect 74 19 75 21
rect 77 19 78 21
rect 74 17 78 19
rect 94 19 95 21
rect 97 19 98 21
rect 94 17 98 19
rect 162 21 186 22
rect 162 17 166 21
rect 53 15 57 17
rect 83 16 89 17
rect 83 14 85 16
rect 87 14 89 16
rect 64 11 68 13
rect 64 9 65 11
rect 67 9 68 11
rect 64 8 68 9
rect 83 8 89 14
rect 94 16 166 17
rect 94 14 117 16
rect 119 14 139 16
rect 141 14 161 16
rect 163 14 166 16
rect 94 13 166 14
rect 170 13 174 15
rect 170 11 171 13
rect 173 11 174 13
rect 170 8 174 11
<< labels >>
rlabel alu0 55 20 55 20 6 n1
rlabel alu0 96 19 96 19 6 n1
rlabel alu0 55 23 55 23 6 n1
rlabel alu0 130 15 130 15 6 n1
rlabel alu0 174 23 174 23 6 n1
rlabel alu1 20 32 20 32 6 b
rlabel alu1 4 28 4 28 6 z
rlabel alu1 28 36 28 36 6 b
rlabel alu1 12 40 12 40 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 52 32 52 32 6 a1
rlabel alu1 60 32 60 32 6 a1
rlabel alu1 68 32 68 32 6 a1
rlabel alu1 36 40 36 40 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 96 4 96 4 6 vss
rlabel alu1 108 24 108 24 6 a2
rlabel alu1 92 32 92 32 6 a2
rlabel alu1 100 32 100 32 6 a2
rlabel alu1 76 32 76 32 6 a1
rlabel alu1 100 40 100 40 6 a1
rlabel alu1 108 40 108 40 6 a1
rlabel alu1 84 40 84 40 6 a1
rlabel alu1 92 40 92 40 6 a1
rlabel alu1 76 48 76 48 6 z
rlabel alu1 100 48 100 48 6 z
rlabel alu1 108 48 108 48 6 z
rlabel alu1 84 48 84 48 6 z
rlabel alu1 92 48 92 48 6 z
rlabel alu1 96 68 96 68 6 vdd
rlabel alu1 116 24 116 24 6 a2
rlabel alu1 132 24 132 24 6 a2
rlabel alu1 140 24 140 24 6 a2
rlabel alu1 148 24 148 24 6 a2
rlabel alu1 124 24 124 24 6 a2
rlabel alu1 116 40 116 40 6 a1
rlabel alu1 132 40 132 40 6 a1
rlabel alu1 140 40 140 40 6 a1
rlabel alu1 148 40 148 40 6 a1
rlabel alu1 124 40 124 40 6 a1
rlabel alu1 116 48 116 48 6 z
rlabel alu1 132 52 132 52 6 z
rlabel alu1 140 48 140 48 6 z
rlabel alu1 148 48 148 48 6 z
rlabel alu1 124 48 124 48 6 z
rlabel alu1 164 32 164 32 6 a2
rlabel alu1 156 28 156 28 6 a2
rlabel alu1 156 40 156 40 6 a1
rlabel alu1 164 40 164 40 6 a1
rlabel alu1 180 36 180 36 6 a1
rlabel alu1 172 44 172 44 6 a1
rlabel alu1 156 48 156 48 6 z
rlabel pdifct1 164 56 164 56 6 z
<< end >>
