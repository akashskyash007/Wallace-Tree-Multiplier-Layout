magic
tech scmos
timestamp 1199202564
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 60 11 64
rect 19 62 21 67
rect 29 62 31 67
rect 39 64 41 68
rect 49 64 51 69
rect 9 38 11 44
rect 19 39 21 44
rect 29 39 31 44
rect 9 36 15 38
rect 9 34 11 36
rect 13 34 15 36
rect 9 32 15 34
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 19 33 31 35
rect 12 29 14 32
rect 19 29 21 33
rect 29 22 31 33
rect 39 31 41 44
rect 49 39 51 42
rect 45 37 51 39
rect 45 35 47 37
rect 49 35 51 37
rect 45 33 51 35
rect 35 29 41 31
rect 49 30 51 33
rect 35 27 37 29
rect 39 27 41 29
rect 35 25 41 27
rect 36 22 38 25
rect 49 15 51 19
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 11
rect 36 6 38 11
<< ndif >>
rect 4 14 12 29
rect 4 12 7 14
rect 9 12 12 14
rect 4 10 12 12
rect 14 10 19 29
rect 21 22 26 29
rect 43 22 49 30
rect 21 20 29 22
rect 21 18 24 20
rect 26 18 29 20
rect 21 11 29 18
rect 31 11 36 22
rect 38 19 49 22
rect 51 28 58 30
rect 51 26 54 28
rect 56 26 58 28
rect 51 24 58 26
rect 51 19 56 24
rect 38 17 43 19
rect 45 17 47 19
rect 38 11 47 17
rect 21 10 26 11
<< pdif >>
rect 34 62 39 64
rect 14 60 19 62
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 44 9 56
rect 11 53 19 60
rect 11 51 14 53
rect 16 51 19 53
rect 11 44 19 51
rect 21 60 29 62
rect 21 58 24 60
rect 26 58 29 60
rect 21 44 29 58
rect 31 60 39 62
rect 31 58 34 60
rect 36 58 39 60
rect 31 53 39 58
rect 31 51 34 53
rect 36 51 39 53
rect 31 44 39 51
rect 41 60 49 64
rect 41 58 44 60
rect 46 58 49 60
rect 41 53 49 58
rect 41 51 44 53
rect 46 51 49 53
rect 41 44 49 51
rect 43 42 49 44
rect 51 55 56 64
rect 51 53 58 55
rect 51 51 54 53
rect 56 51 58 53
rect 51 46 58 51
rect 51 44 54 46
rect 56 44 58 46
rect 51 42 58 44
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 33 60 38 63
rect 33 58 34 60
rect 36 58 38 60
rect 33 54 38 58
rect 12 53 38 54
rect 12 51 14 53
rect 16 51 34 53
rect 36 51 38 53
rect 12 50 38 51
rect 2 22 6 47
rect 17 42 30 46
rect 26 37 30 42
rect 41 39 47 46
rect 26 35 27 37
rect 29 35 30 37
rect 26 33 30 35
rect 34 37 50 39
rect 34 35 47 37
rect 49 35 50 37
rect 34 33 50 35
rect 2 20 28 22
rect 2 18 24 20
rect 26 18 28 20
rect 22 17 28 18
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 12 10 14 29
rect 19 10 21 29
rect 29 11 31 22
rect 36 11 38 22
rect 49 19 51 30
<< pmos >>
rect 9 44 11 60
rect 19 44 21 62
rect 29 44 31 62
rect 39 44 41 64
rect 49 42 51 64
<< polyct0 >>
rect 11 34 13 36
rect 37 27 39 29
<< polyct1 >>
rect 27 35 29 37
rect 47 35 49 37
<< ndifct0 >>
rect 7 12 9 14
rect 54 26 56 28
rect 43 17 45 19
<< ndifct1 >>
rect 24 18 26 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 56 6 58
rect 24 58 26 60
rect 44 58 46 60
rect 44 51 46 53
rect 54 51 56 53
rect 54 44 56 46
<< pdifct1 >>
rect 14 51 16 53
rect 34 58 36 60
rect 34 51 36 53
<< alu0 >>
rect 3 58 7 68
rect 3 56 4 58
rect 6 56 7 58
rect 22 60 28 68
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 3 54 7 56
rect 10 50 12 54
rect 42 60 48 68
rect 42 58 44 60
rect 46 58 48 60
rect 42 53 48 58
rect 42 51 44 53
rect 46 51 48 53
rect 42 50 48 51
rect 53 53 57 55
rect 53 51 54 53
rect 56 51 57 53
rect 10 47 14 50
rect 6 43 14 47
rect 53 46 57 51
rect 10 36 14 38
rect 10 34 11 36
rect 13 34 14 36
rect 10 30 14 34
rect 53 44 54 46
rect 56 44 57 46
rect 53 30 57 44
rect 10 29 57 30
rect 10 27 37 29
rect 39 28 57 29
rect 39 27 54 28
rect 10 26 54 27
rect 56 26 57 28
rect 53 24 57 26
rect 42 19 46 21
rect 42 17 43 19
rect 45 17 46 19
rect 5 14 11 15
rect 5 12 7 14
rect 9 12 11 14
rect 42 12 46 17
<< labels >>
rlabel alu0 12 32 12 32 6 an
rlabel alu0 33 28 33 28 6 an
rlabel alu0 55 39 55 39 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel polyct1 28 36 28 36 6 b
rlabel alu1 20 44 20 44 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 36 36 36 6 a
rlabel alu1 44 40 44 40 6 a
rlabel alu1 36 60 36 60 6 z
rlabel alu1 32 74 32 74 6 vdd
<< end >>
