magic
tech scmos
timestamp 1199203242
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 63 11 68
rect 19 62 25 64
rect 19 60 21 62
rect 23 60 25 62
rect 19 58 25 60
rect 22 55 24 58
rect 29 55 31 60
rect 9 41 11 45
rect 9 39 15 41
rect 9 37 11 39
rect 13 37 15 39
rect 22 37 24 45
rect 9 35 15 37
rect 19 35 24 37
rect 29 39 31 45
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 9 30 11 35
rect 19 30 21 35
rect 29 33 35 35
rect 29 30 31 33
rect 9 16 11 21
rect 19 19 21 24
rect 29 19 31 24
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 21 9 24
rect 11 24 19 30
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 24 29 26
rect 31 28 38 30
rect 31 26 34 28
rect 36 26 38 28
rect 31 24 38 26
rect 11 21 17 24
rect 13 17 17 21
rect 13 15 19 17
rect 13 13 15 15
rect 17 13 19 15
rect 13 11 19 13
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 66 19 69
rect 13 63 17 66
rect 4 58 9 63
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 11 55 17 63
rect 11 45 22 55
rect 24 45 29 55
rect 31 53 38 55
rect 31 51 34 53
rect 36 51 38 53
rect 31 49 38 51
rect 31 45 36 49
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 71 42 79
rect -2 69 15 71
rect 17 69 42 71
rect -2 68 42 69
rect 2 56 6 63
rect 10 62 25 63
rect 10 60 21 62
rect 23 60 25 62
rect 2 54 4 56
rect 2 49 6 54
rect 2 47 4 49
rect 2 31 6 47
rect 10 57 25 60
rect 10 49 14 57
rect 34 39 38 47
rect 2 28 14 31
rect 2 26 4 28
rect 6 26 14 28
rect 2 25 14 26
rect 26 37 38 39
rect 26 35 31 37
rect 33 35 38 37
rect 26 33 38 35
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 21 11 30
rect 19 24 21 30
rect 29 24 31 30
<< pmos >>
rect 9 45 11 63
rect 22 45 24 55
rect 29 45 31 55
<< polyct0 >>
rect 11 37 13 39
<< polyct1 >>
rect 21 60 23 62
rect 31 35 33 37
<< ndifct0 >>
rect 24 26 26 28
rect 34 26 36 28
rect 15 13 17 15
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 34 51 36 53
<< pdifct1 >>
rect 15 69 17 71
rect 4 54 6 56
rect 4 47 6 49
<< alu0 >>
rect 6 45 7 58
rect 18 53 38 54
rect 18 51 34 53
rect 36 51 38 53
rect 18 50 38 51
rect 18 41 22 50
rect 10 39 22 41
rect 10 37 11 39
rect 13 37 22 39
rect 10 35 22 37
rect 18 29 22 35
rect 18 28 28 29
rect 18 26 24 28
rect 26 26 28 28
rect 18 25 28 26
rect 32 28 38 29
rect 32 26 34 28
rect 36 26 38 28
rect 14 15 18 17
rect 14 13 15 15
rect 17 13 18 15
rect 14 12 18 13
rect 32 12 38 26
<< labels >>
rlabel alu0 23 27 23 27 6 zn
rlabel alu0 16 38 16 38 6 zn
rlabel alu0 28 52 28 52 6 zn
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 56 12 56 6 a
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 60 20 60 6 a
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 40 36 40 6 b
<< end >>
