magic
tech scmos
timestamp 1199203542
<< ab >>
rect 0 0 160 80
<< nwell >>
rect -5 36 165 88
<< pwell >>
rect -5 -8 165 36
<< poly >>
rect 22 70 24 74
rect 29 70 31 74
rect 39 70 41 74
rect 46 70 48 74
rect 56 70 58 74
rect 66 70 68 74
rect 76 70 78 74
rect 86 70 88 74
rect 93 70 95 74
rect 104 72 130 74
rect 104 64 106 72
rect 111 64 113 68
rect 121 64 123 68
rect 128 64 130 72
rect 139 70 141 74
rect 149 70 151 74
rect 22 39 24 42
rect 20 36 24 39
rect 29 39 31 42
rect 39 39 41 42
rect 29 37 42 39
rect 20 30 22 36
rect 29 35 31 37
rect 33 35 38 37
rect 40 35 42 37
rect 29 33 42 35
rect 46 35 48 42
rect 56 39 58 42
rect 66 39 68 42
rect 76 39 78 42
rect 86 39 88 42
rect 56 37 78 39
rect 82 37 88 39
rect 93 39 95 42
rect 104 39 106 42
rect 93 37 106 39
rect 46 33 52 35
rect 30 30 32 33
rect 40 30 42 33
rect 50 30 52 33
rect 72 31 74 37
rect 82 35 84 37
rect 86 35 88 37
rect 82 33 88 35
rect 72 29 78 31
rect 72 27 74 29
rect 76 27 78 29
rect 72 25 78 27
rect 82 23 84 33
rect 104 28 106 37
rect 111 39 113 42
rect 121 39 123 42
rect 128 39 130 42
rect 139 39 141 42
rect 149 39 151 42
rect 111 37 123 39
rect 127 37 133 39
rect 111 35 113 37
rect 115 35 117 37
rect 111 33 117 35
rect 127 35 129 37
rect 131 35 133 37
rect 127 33 133 35
rect 137 37 151 39
rect 137 35 139 37
rect 141 35 143 37
rect 137 33 143 35
rect 92 26 106 28
rect 92 23 94 26
rect 104 23 106 26
rect 114 23 116 33
rect 137 28 139 33
rect 127 26 139 28
rect 127 23 129 26
rect 137 23 139 26
rect 59 20 65 22
rect 59 18 61 20
rect 63 18 65 20
rect 59 16 65 18
rect 20 8 22 16
rect 30 12 32 16
rect 40 12 42 16
rect 50 13 52 16
rect 59 13 61 16
rect 50 11 61 13
rect 50 8 52 11
rect 20 6 52 8
rect 82 6 84 11
rect 92 6 94 11
rect 104 6 106 11
rect 114 6 116 11
rect 127 6 129 10
rect 137 6 139 10
<< ndif >>
rect 13 28 20 30
rect 13 26 15 28
rect 17 26 20 28
rect 13 24 20 26
rect 15 16 20 24
rect 22 28 30 30
rect 22 26 25 28
rect 27 26 30 28
rect 22 21 30 26
rect 22 19 25 21
rect 27 19 30 21
rect 22 16 30 19
rect 32 20 40 30
rect 32 18 35 20
rect 37 18 40 20
rect 32 16 40 18
rect 42 28 50 30
rect 42 26 45 28
rect 47 26 50 28
rect 42 16 50 26
rect 52 28 59 30
rect 52 26 55 28
rect 57 26 59 28
rect 52 24 59 26
rect 52 16 57 24
rect 74 11 82 23
rect 84 20 92 23
rect 84 18 87 20
rect 89 18 92 20
rect 84 11 92 18
rect 94 11 104 23
rect 106 20 114 23
rect 106 18 109 20
rect 111 18 114 20
rect 106 11 114 18
rect 116 11 127 23
rect 74 9 76 11
rect 78 9 80 11
rect 74 7 80 9
rect 96 9 98 11
rect 100 9 102 11
rect 96 7 102 9
rect 118 9 120 11
rect 122 10 127 11
rect 129 20 137 23
rect 129 18 132 20
rect 134 18 137 20
rect 129 10 137 18
rect 139 11 147 23
rect 139 10 143 11
rect 122 9 124 10
rect 118 7 124 9
rect 141 9 143 10
rect 145 9 147 11
rect 141 7 147 9
<< pdif >>
rect 17 55 22 70
rect 15 53 22 55
rect 15 51 17 53
rect 19 51 22 53
rect 15 46 22 51
rect 15 44 17 46
rect 19 44 22 46
rect 15 42 22 44
rect 24 42 29 70
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 60 39 66
rect 31 58 34 60
rect 36 58 39 60
rect 31 42 39 58
rect 41 42 46 70
rect 48 61 56 70
rect 48 59 51 61
rect 53 59 56 61
rect 48 42 56 59
rect 58 46 66 70
rect 58 44 61 46
rect 63 44 66 46
rect 58 42 66 44
rect 68 61 76 70
rect 68 59 71 61
rect 73 59 76 61
rect 68 42 76 59
rect 78 46 86 70
rect 78 44 81 46
rect 83 44 86 46
rect 78 42 86 44
rect 88 42 93 70
rect 95 68 102 70
rect 95 66 98 68
rect 100 66 102 68
rect 95 64 102 66
rect 132 68 139 70
rect 132 66 134 68
rect 136 66 139 68
rect 132 64 139 66
rect 95 42 104 64
rect 106 42 111 64
rect 113 53 121 64
rect 113 51 116 53
rect 118 51 121 53
rect 113 46 121 51
rect 113 44 116 46
rect 118 44 121 46
rect 113 42 121 44
rect 123 42 128 64
rect 130 61 139 64
rect 130 59 134 61
rect 136 59 139 61
rect 130 42 139 59
rect 141 61 149 70
rect 141 59 144 61
rect 146 59 149 61
rect 141 54 149 59
rect 141 52 144 54
rect 146 52 149 54
rect 141 42 149 52
rect 151 63 158 70
rect 151 61 154 63
rect 156 61 158 63
rect 151 42 158 61
<< alu1 >>
rect -2 81 162 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 162 81
rect -2 68 162 79
rect 42 61 79 62
rect 42 59 51 61
rect 53 59 71 61
rect 73 59 79 61
rect 42 58 79 59
rect 2 46 20 47
rect 42 46 46 58
rect 2 44 17 46
rect 19 44 46 46
rect 2 42 46 44
rect 2 21 6 42
rect 24 28 49 30
rect 24 26 25 28
rect 27 26 45 28
rect 47 26 49 28
rect 24 25 49 26
rect 24 21 28 25
rect 105 38 111 46
rect 130 38 134 47
rect 81 37 117 38
rect 81 35 84 37
rect 86 35 113 37
rect 115 35 117 37
rect 81 34 117 35
rect 121 37 134 38
rect 121 35 129 37
rect 131 35 134 37
rect 121 34 134 35
rect 138 37 142 47
rect 138 35 139 37
rect 141 35 142 37
rect 138 30 142 35
rect 72 29 142 30
rect 72 27 74 29
rect 76 27 142 29
rect 72 26 142 27
rect 2 19 25 21
rect 27 19 28 21
rect 2 17 28 19
rect 122 17 126 26
rect -2 11 162 12
rect -2 9 76 11
rect 78 9 98 11
rect 100 9 120 11
rect 122 9 143 11
rect 145 9 162 11
rect -2 1 162 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 162 1
rect -2 -2 162 -1
<< ptie >>
rect 0 1 160 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 160 1
rect 0 -3 160 -1
<< ntie >>
rect 0 81 160 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 160 81
rect 0 77 160 79
<< nmos >>
rect 20 16 22 30
rect 30 16 32 30
rect 40 16 42 30
rect 50 16 52 30
rect 82 11 84 23
rect 92 11 94 23
rect 104 11 106 23
rect 114 11 116 23
rect 127 10 129 23
rect 137 10 139 23
<< pmos >>
rect 22 42 24 70
rect 29 42 31 70
rect 39 42 41 70
rect 46 42 48 70
rect 56 42 58 70
rect 66 42 68 70
rect 76 42 78 70
rect 86 42 88 70
rect 93 42 95 70
rect 104 42 106 64
rect 111 42 113 64
rect 121 42 123 64
rect 128 42 130 64
rect 139 42 141 70
rect 149 42 151 70
<< polyct0 >>
rect 31 35 33 37
rect 38 35 40 37
rect 61 18 63 20
<< polyct1 >>
rect 84 35 86 37
rect 74 27 76 29
rect 113 35 115 37
rect 129 35 131 37
rect 139 35 141 37
<< ndifct0 >>
rect 15 26 17 28
rect 35 18 37 20
rect 55 26 57 28
rect 87 18 89 20
rect 109 18 111 20
rect 132 18 134 20
<< ndifct1 >>
rect 25 26 27 28
rect 25 19 27 21
rect 45 26 47 28
rect 76 9 78 11
rect 98 9 100 11
rect 120 9 122 11
rect 143 9 145 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
<< pdifct0 >>
rect 17 51 19 53
rect 34 66 36 68
rect 34 58 36 60
rect 61 44 63 46
rect 81 44 83 46
rect 98 66 100 68
rect 134 66 136 68
rect 116 51 118 53
rect 116 44 118 46
rect 134 59 136 61
rect 144 59 146 61
rect 144 52 146 54
rect 154 61 156 63
<< pdifct1 >>
rect 17 44 19 46
rect 51 59 53 61
rect 71 59 73 61
<< alu0 >>
rect 33 66 34 68
rect 36 66 37 68
rect 33 60 37 66
rect 96 66 98 68
rect 100 66 102 68
rect 96 65 102 66
rect 132 66 134 68
rect 136 66 138 68
rect 33 58 34 60
rect 36 58 37 60
rect 33 56 37 58
rect 86 58 128 62
rect 132 61 138 66
rect 153 63 157 68
rect 132 59 134 61
rect 136 59 138 61
rect 132 58 138 59
rect 143 61 148 62
rect 143 59 144 61
rect 146 59 148 61
rect 153 61 154 63
rect 156 61 157 63
rect 153 59 157 61
rect 16 53 20 55
rect 16 51 17 53
rect 19 51 20 53
rect 16 47 20 51
rect 86 55 90 58
rect 50 51 90 55
rect 124 55 128 58
rect 143 55 148 59
rect 124 54 150 55
rect 94 53 120 54
rect 94 51 116 53
rect 118 51 120 53
rect 124 52 144 54
rect 146 52 150 54
rect 124 51 150 52
rect 50 38 54 51
rect 94 50 120 51
rect 94 47 98 50
rect 59 46 98 47
rect 115 46 120 50
rect 59 44 61 46
rect 63 44 81 46
rect 83 44 98 46
rect 59 43 98 44
rect 13 37 59 38
rect 13 35 31 37
rect 33 35 38 37
rect 40 35 59 37
rect 13 34 59 35
rect 13 28 19 34
rect 13 26 15 28
rect 17 26 19 28
rect 13 25 19 26
rect 53 28 59 34
rect 53 26 55 28
rect 57 26 59 28
rect 53 25 59 26
rect 64 21 68 43
rect 115 44 116 46
rect 118 44 120 46
rect 115 42 120 44
rect 33 20 113 21
rect 33 18 35 20
rect 37 18 61 20
rect 63 18 87 20
rect 89 18 109 20
rect 111 18 113 20
rect 33 17 113 18
rect 146 21 150 51
rect 130 20 150 21
rect 130 18 132 20
rect 134 18 150 20
rect 130 17 150 18
<< labels >>
rlabel alu0 16 31 16 31 6 bn
rlabel alu0 56 31 56 31 6 bn
rlabel alu0 73 19 73 19 6 an
rlabel alu0 78 45 78 45 6 an
rlabel alu0 117 48 117 48 6 an
rlabel alu0 107 52 107 52 6 an
rlabel alu0 140 19 140 19 6 bn
rlabel alu0 137 53 137 53 6 bn
rlabel alu0 145 56 145 56 6 bn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 28 28 28 28 6 z
rlabel alu1 36 28 36 28 6 z
rlabel alu1 44 28 44 28 6 z
rlabel alu1 28 44 28 44 6 z
rlabel alu1 36 44 36 44 6 z
rlabel alu1 44 52 44 52 6 z
rlabel pdifct1 52 60 52 60 6 z
rlabel alu1 60 60 60 60 6 z
rlabel alu1 80 6 80 6 6 vss
rlabel alu1 76 28 76 28 6 b
rlabel alu1 84 28 84 28 6 b
rlabel alu1 92 28 92 28 6 b
rlabel alu1 84 36 84 36 6 a2
rlabel alu1 92 36 92 36 6 a2
rlabel alu1 68 60 68 60 6 z
rlabel alu1 76 60 76 60 6 z
rlabel alu1 80 74 80 74 6 vdd
rlabel alu1 100 28 100 28 6 b
rlabel alu1 108 28 108 28 6 b
rlabel alu1 116 28 116 28 6 b
rlabel alu1 124 24 124 24 6 b
rlabel alu1 100 36 100 36 6 a2
rlabel alu1 108 40 108 40 6 a2
rlabel alu1 124 36 124 36 6 a1
rlabel alu1 132 28 132 28 6 b
rlabel alu1 132 44 132 44 6 a1
rlabel alu1 140 40 140 40 6 b
<< end >>
