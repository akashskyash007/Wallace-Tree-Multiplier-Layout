magic
tech scmos
timestamp 1199469652
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 83 49 88
rect 11 52 13 55
rect 23 52 25 55
rect 11 50 25 52
rect 11 48 21 50
rect 23 48 25 50
rect 11 46 25 48
rect 11 35 13 46
rect 23 35 25 46
rect 35 52 37 55
rect 47 52 49 55
rect 35 50 49 52
rect 35 48 37 50
rect 39 48 49 50
rect 35 46 49 48
rect 35 35 37 46
rect 47 35 49 46
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 47 12 49 17
<< ndif >>
rect 3 31 11 35
rect 3 29 5 31
rect 7 29 11 31
rect 3 21 11 29
rect 3 19 5 21
rect 7 19 11 21
rect 3 17 11 19
rect 13 31 23 35
rect 13 29 17 31
rect 19 29 23 31
rect 13 21 23 29
rect 13 19 17 21
rect 19 19 23 21
rect 13 17 23 19
rect 25 31 35 35
rect 25 29 29 31
rect 31 29 35 31
rect 25 21 35 29
rect 25 19 29 21
rect 31 19 35 21
rect 25 17 35 19
rect 37 31 47 35
rect 37 29 41 31
rect 43 29 47 31
rect 37 21 47 29
rect 37 19 41 21
rect 43 19 47 21
rect 37 17 47 19
rect 49 31 57 35
rect 49 29 53 31
rect 55 29 57 31
rect 49 21 57 29
rect 49 19 53 21
rect 55 19 57 21
rect 49 17 57 19
<< pdif >>
rect 3 91 11 94
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 55 11 69
rect 13 71 23 94
rect 13 69 17 71
rect 19 69 23 71
rect 13 61 23 69
rect 13 59 17 61
rect 19 59 23 61
rect 13 55 23 59
rect 25 91 35 94
rect 25 89 29 91
rect 31 89 35 91
rect 25 81 35 89
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 55 35 69
rect 37 83 42 94
rect 37 71 47 83
rect 37 69 41 71
rect 43 69 47 71
rect 37 61 47 69
rect 37 59 41 61
rect 43 59 47 61
rect 37 55 47 59
rect 49 81 57 83
rect 49 79 53 81
rect 55 79 57 81
rect 49 71 57 79
rect 49 69 53 71
rect 55 69 57 71
rect 49 55 57 69
<< alu1 >>
rect -2 95 62 100
rect -2 93 51 95
rect 53 93 62 95
rect -2 91 62 93
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 62 91
rect -2 88 62 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 28 81 32 88
rect 28 79 29 81
rect 31 79 32 81
rect 4 69 5 71
rect 7 69 8 71
rect 4 67 8 69
rect 16 71 22 73
rect 16 69 17 71
rect 19 69 22 71
rect 16 63 22 69
rect 28 71 32 79
rect 52 81 56 88
rect 52 79 53 81
rect 55 79 56 81
rect 28 69 29 71
rect 31 69 32 71
rect 28 67 32 69
rect 38 71 44 73
rect 38 69 41 71
rect 43 69 44 71
rect 38 63 44 69
rect 52 71 56 79
rect 52 69 53 71
rect 55 69 56 71
rect 52 67 56 69
rect 8 61 44 63
rect 8 59 17 61
rect 19 59 41 61
rect 43 59 44 61
rect 8 58 44 59
rect 8 42 12 58
rect 48 52 52 63
rect 17 50 52 52
rect 17 48 21 50
rect 23 48 37 50
rect 39 48 52 50
rect 17 47 52 48
rect 8 37 44 42
rect 48 37 52 47
rect 4 31 8 33
rect 4 29 5 31
rect 7 29 8 31
rect 4 21 8 29
rect 4 19 5 21
rect 7 19 8 21
rect 4 12 8 19
rect 16 31 22 37
rect 16 29 17 31
rect 19 29 22 31
rect 16 21 22 29
rect 16 19 17 21
rect 19 19 22 21
rect 16 17 22 19
rect 28 31 32 33
rect 28 29 29 31
rect 31 29 32 31
rect 28 21 32 29
rect 28 19 29 21
rect 31 19 32 21
rect 28 12 32 19
rect 38 31 44 37
rect 38 29 41 31
rect 43 29 44 31
rect 38 21 44 29
rect 38 19 41 21
rect 43 19 44 21
rect 38 17 44 19
rect 52 31 56 33
rect 52 29 53 31
rect 55 29 56 31
rect 52 21 56 29
rect 52 19 53 21
rect 55 19 56 21
rect 52 12 56 19
rect -2 7 62 12
rect -2 5 22 7
rect 24 5 32 7
rect 34 5 62 7
rect -2 0 62 5
<< ptie >>
rect 20 7 36 9
rect 20 5 22 7
rect 24 5 32 7
rect 34 5 36 7
rect 20 3 36 5
<< ntie >>
rect 49 95 55 97
rect 49 93 51 95
rect 53 93 55 95
rect 49 91 55 93
<< nmos >>
rect 11 17 13 35
rect 23 17 25 35
rect 35 17 37 35
rect 47 17 49 35
<< pmos >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 55 37 94
rect 47 55 49 83
<< polyct1 >>
rect 21 48 23 50
rect 37 48 39 50
<< ndifct1 >>
rect 5 29 7 31
rect 5 19 7 21
rect 17 29 19 31
rect 17 19 19 21
rect 29 29 31 31
rect 29 19 31 21
rect 41 29 43 31
rect 41 19 43 21
rect 53 29 55 31
rect 53 19 55 21
<< ntiect1 >>
rect 51 93 53 95
<< ptiect1 >>
rect 22 5 24 7
rect 32 5 34 7
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 5 69 7 71
rect 17 69 19 71
rect 17 59 19 61
rect 29 89 31 91
rect 29 79 31 81
rect 29 69 31 71
rect 41 69 43 71
rect 41 59 43 61
rect 53 79 55 81
rect 53 69 55 71
<< labels >>
rlabel alu1 10 50 10 50 6 z
rlabel alu1 20 30 20 30 6 z
rlabel alu1 20 50 20 50 6 a
rlabel alu1 20 65 20 65 6 z
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 30 40 30 40 6 z
rlabel alu1 40 30 40 30 6 z
rlabel alu1 40 50 40 50 6 a
rlabel alu1 30 50 30 50 6 a
rlabel alu1 30 60 30 60 6 z
rlabel alu1 40 65 40 65 6 z
rlabel alu1 30 94 30 94 6 vdd
rlabel alu1 50 50 50 50 6 a
<< end >>
