magic
tech scmos
timestamp 1199202340
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 11 58 13 63
rect 21 58 23 63
rect 11 39 13 42
rect 21 39 23 42
rect 11 37 23 39
rect 11 35 19 37
rect 21 35 23 37
rect 11 33 23 35
rect 15 30 17 33
rect 15 17 17 22
<< ndif >>
rect 8 28 15 30
rect 8 26 10 28
rect 12 26 15 28
rect 8 24 15 26
rect 10 22 15 24
rect 17 26 25 30
rect 17 24 20 26
rect 22 24 25 26
rect 17 22 25 24
<< pdif >>
rect 2 56 11 58
rect 2 54 4 56
rect 6 54 11 56
rect 2 49 11 54
rect 2 47 4 49
rect 6 47 11 49
rect 2 42 11 47
rect 13 54 21 58
rect 13 52 16 54
rect 18 52 21 54
rect 13 47 21 52
rect 13 45 16 47
rect 18 45 21 47
rect 13 42 21 45
rect 23 56 30 58
rect 23 54 26 56
rect 28 54 30 56
rect 23 49 30 54
rect 23 47 26 49
rect 28 47 30 49
rect 23 42 30 47
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 15 54 22 56
rect 15 52 16 54
rect 18 52 22 54
rect 15 49 22 52
rect 15 47 19 49
rect 10 45 16 47
rect 18 45 19 47
rect 10 43 19 45
rect 10 30 14 43
rect 18 37 30 39
rect 18 35 19 37
rect 21 35 30 37
rect 18 33 30 35
rect 9 28 14 30
rect 9 26 10 28
rect 12 26 14 28
rect 9 24 14 26
rect 26 25 30 33
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 15 22 17 30
<< pmos >>
rect 11 42 13 58
rect 21 42 23 58
<< polyct1 >>
rect 19 35 21 37
<< ndifct0 >>
rect 20 24 22 26
<< ndifct1 >>
rect 10 26 12 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 54 6 56
rect 4 47 6 49
rect 26 54 28 56
rect 26 47 28 49
<< pdifct1 >>
rect 16 52 18 54
rect 16 45 18 47
<< alu0 >>
rect 3 56 7 68
rect 25 56 29 68
rect 3 54 4 56
rect 6 54 7 56
rect 3 49 7 54
rect 3 47 4 49
rect 6 47 7 49
rect 25 54 26 56
rect 28 54 29 56
rect 25 49 29 54
rect 3 45 7 47
rect 25 47 26 49
rect 28 47 29 49
rect 25 45 29 47
rect 19 26 23 28
rect 19 24 20 26
rect 22 24 23 26
rect 19 12 23 24
<< labels >>
rlabel alu1 12 36 12 36 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel polyct1 20 36 20 36 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 32 28 32 6 a
<< end >>
