magic
tech scmos
timestamp 1199542023
<< ab >>
rect 0 0 180 100
<< nwell >>
rect -2 48 182 104
<< pwell >>
rect -2 -4 182 48
<< poly >>
rect 11 95 13 98
rect 23 95 25 98
rect 155 95 157 98
rect 167 95 169 98
rect 35 83 37 86
rect 47 83 49 86
rect 83 77 85 80
rect 95 77 97 80
rect 107 77 109 80
rect 119 77 121 80
rect 131 77 133 80
rect 71 71 73 74
rect 11 43 13 55
rect 23 43 25 55
rect 35 53 37 65
rect 47 63 49 65
rect 47 61 53 63
rect 47 59 49 61
rect 51 59 53 61
rect 47 57 53 59
rect 29 51 37 53
rect 71 53 73 55
rect 83 53 85 55
rect 71 51 85 53
rect 95 53 97 55
rect 95 51 103 53
rect 29 49 31 51
rect 33 49 37 51
rect 29 47 37 49
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 97 49 99 51
rect 101 49 103 51
rect 97 47 103 49
rect 11 41 25 43
rect 37 41 43 43
rect 11 39 39 41
rect 41 39 43 41
rect 11 37 25 39
rect 37 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 63 41 69 43
rect 107 41 109 55
rect 119 43 121 55
rect 131 53 133 55
rect 127 51 133 53
rect 127 49 129 51
rect 131 49 133 51
rect 127 47 133 49
rect 155 43 157 55
rect 167 43 169 55
rect 63 39 65 41
rect 67 39 109 41
rect 63 37 69 39
rect 11 25 13 37
rect 23 25 25 37
rect 29 31 37 33
rect 29 29 31 31
rect 33 29 37 31
rect 47 29 49 37
rect 97 33 103 35
rect 77 31 83 33
rect 97 31 99 33
rect 101 31 103 33
rect 77 29 79 31
rect 81 29 83 31
rect 95 29 103 31
rect 29 27 37 29
rect 35 25 37 27
rect 71 27 85 29
rect 95 27 97 29
rect 107 27 109 39
rect 117 41 123 43
rect 137 41 143 43
rect 117 39 119 41
rect 121 39 139 41
rect 141 39 143 41
rect 117 37 123 39
rect 137 37 143 39
rect 147 41 169 43
rect 147 39 149 41
rect 151 39 169 41
rect 147 37 169 39
rect 127 31 133 33
rect 127 29 129 31
rect 131 29 133 31
rect 119 27 133 29
rect 71 25 73 27
rect 83 25 85 27
rect 35 12 37 15
rect 47 12 49 15
rect 71 14 73 17
rect 119 25 121 27
rect 131 25 133 27
rect 155 25 157 37
rect 167 25 169 37
rect 83 12 85 15
rect 95 12 97 15
rect 107 12 109 15
rect 119 12 121 15
rect 131 14 133 17
rect 11 2 13 5
rect 23 2 25 5
rect 155 2 157 5
rect 167 2 169 5
<< ndif >>
rect 39 25 47 29
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 11 11 19
rect 3 9 5 11
rect 7 9 11 11
rect 3 5 11 9
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 5 23 19
rect 25 15 35 25
rect 37 15 47 25
rect 49 21 57 29
rect 87 25 95 27
rect 49 19 53 21
rect 55 19 57 21
rect 49 15 57 19
rect 63 21 71 25
rect 63 19 65 21
rect 67 19 71 21
rect 63 17 71 19
rect 73 17 83 25
rect 25 11 33 15
rect 75 15 83 17
rect 85 15 95 25
rect 97 23 107 27
rect 97 21 101 23
rect 103 21 107 23
rect 97 15 107 21
rect 109 25 117 27
rect 135 31 143 33
rect 135 29 139 31
rect 141 29 143 31
rect 135 27 143 29
rect 135 25 141 27
rect 109 15 119 25
rect 121 17 131 25
rect 133 17 141 25
rect 151 21 155 25
rect 121 15 129 17
rect 25 9 29 11
rect 31 9 33 11
rect 75 11 81 15
rect 75 9 77 11
rect 79 9 81 11
rect 123 11 129 15
rect 123 9 125 11
rect 127 9 129 11
rect 25 5 33 9
rect 75 7 81 9
rect 123 7 129 9
rect 147 11 155 21
rect 147 9 149 11
rect 151 9 155 11
rect 147 5 155 9
rect 157 21 167 25
rect 157 19 161 21
rect 163 19 167 21
rect 157 5 167 19
rect 169 21 177 25
rect 169 19 173 21
rect 175 19 177 21
rect 169 11 177 19
rect 169 9 173 11
rect 175 9 177 11
rect 169 5 177 9
<< pdif >>
rect 3 91 11 95
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 81 23 95
rect 13 79 17 81
rect 19 79 23 81
rect 13 71 23 79
rect 13 69 17 71
rect 19 69 23 71
rect 13 61 23 69
rect 13 59 17 61
rect 19 59 23 61
rect 13 55 23 59
rect 25 91 33 95
rect 25 89 29 91
rect 31 89 33 91
rect 25 83 33 89
rect 51 91 57 93
rect 51 89 53 91
rect 55 89 57 91
rect 51 83 57 89
rect 75 91 81 93
rect 123 91 129 93
rect 75 89 77 91
rect 79 89 81 91
rect 25 65 35 83
rect 37 71 47 83
rect 37 69 41 71
rect 43 69 47 71
rect 37 65 47 69
rect 49 65 57 83
rect 75 77 81 89
rect 123 89 125 91
rect 127 89 129 91
rect 123 77 129 89
rect 147 91 155 95
rect 147 89 149 91
rect 151 89 155 91
rect 147 81 155 89
rect 147 79 149 81
rect 151 79 155 81
rect 75 71 83 77
rect 25 55 33 65
rect 63 61 71 71
rect 63 59 65 61
rect 67 59 71 61
rect 63 55 71 59
rect 73 55 83 71
rect 85 71 95 77
rect 85 69 89 71
rect 91 69 95 71
rect 85 55 95 69
rect 97 61 107 77
rect 97 59 101 61
rect 103 59 107 61
rect 97 55 107 59
rect 109 71 119 77
rect 109 69 113 71
rect 115 69 119 71
rect 109 61 119 69
rect 109 59 113 61
rect 115 59 119 61
rect 109 55 119 59
rect 121 55 131 77
rect 133 61 141 77
rect 147 71 155 79
rect 147 69 149 71
rect 151 69 155 71
rect 147 67 155 69
rect 133 59 143 61
rect 133 57 139 59
rect 141 57 143 59
rect 133 55 143 57
rect 151 55 155 67
rect 157 81 167 95
rect 157 79 161 81
rect 163 79 167 81
rect 157 71 167 79
rect 157 69 161 71
rect 163 69 167 71
rect 157 61 167 69
rect 157 59 161 61
rect 163 59 167 61
rect 157 55 167 59
rect 169 91 177 95
rect 169 89 173 91
rect 175 89 177 91
rect 169 81 177 89
rect 169 79 173 81
rect 175 79 177 81
rect 169 71 177 79
rect 169 69 173 71
rect 175 69 177 71
rect 169 61 177 69
rect 169 59 173 61
rect 175 59 177 61
rect 169 55 177 59
<< alu1 >>
rect -2 95 182 100
rect -2 93 65 95
rect 67 93 89 95
rect 91 93 101 95
rect 103 93 113 95
rect 115 93 137 95
rect 139 93 182 95
rect -2 91 182 93
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 53 91
rect 55 89 77 91
rect 79 89 125 91
rect 127 89 149 91
rect 151 89 173 91
rect 175 89 182 91
rect -2 88 182 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 16 81 22 82
rect 16 79 17 81
rect 19 79 22 81
rect 16 78 22 79
rect 18 72 22 78
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 16 71 22 72
rect 16 69 17 71
rect 19 69 22 71
rect 16 68 22 69
rect 18 62 22 68
rect 4 59 5 61
rect 7 59 8 61
rect 4 58 8 59
rect 16 61 22 62
rect 16 59 17 61
rect 19 59 22 61
rect 16 58 22 59
rect 18 22 22 58
rect 4 21 8 22
rect 4 19 5 21
rect 7 19 8 21
rect 4 12 8 19
rect 16 21 22 22
rect 16 19 17 21
rect 19 19 22 21
rect 16 18 22 19
rect 28 81 32 82
rect 148 81 152 88
rect 28 79 131 81
rect 28 52 32 79
rect 40 71 44 72
rect 78 71 82 72
rect 40 69 41 71
rect 43 69 44 71
rect 40 68 44 69
rect 51 69 82 71
rect 28 51 34 52
rect 28 49 31 51
rect 33 49 34 51
rect 28 48 34 49
rect 28 32 32 48
rect 40 42 42 68
rect 51 62 53 69
rect 48 61 53 62
rect 48 59 49 61
rect 51 59 53 61
rect 64 61 68 62
rect 64 59 65 61
rect 67 59 68 61
rect 48 58 52 59
rect 64 58 68 59
rect 49 42 51 58
rect 65 42 67 58
rect 78 51 82 69
rect 88 71 92 72
rect 112 71 116 72
rect 88 69 89 71
rect 91 69 113 71
rect 115 69 116 71
rect 88 68 92 69
rect 112 68 116 69
rect 113 62 115 68
rect 100 61 104 62
rect 78 49 79 51
rect 81 49 82 51
rect 38 41 42 42
rect 38 39 39 41
rect 41 39 42 41
rect 38 38 42 39
rect 48 41 52 42
rect 48 39 49 41
rect 51 39 52 41
rect 48 38 52 39
rect 64 41 68 42
rect 64 39 65 41
rect 67 39 68 41
rect 64 38 68 39
rect 28 31 34 32
rect 28 29 31 31
rect 33 29 34 31
rect 28 28 34 29
rect 28 18 32 28
rect 40 21 42 38
rect 65 22 67 38
rect 78 31 82 49
rect 78 29 79 31
rect 81 29 82 31
rect 52 21 56 22
rect 40 19 53 21
rect 55 19 56 21
rect 52 18 56 19
rect 64 21 68 22
rect 64 19 65 21
rect 67 19 68 21
rect 64 18 68 19
rect 78 18 82 29
rect 89 59 101 61
rect 103 59 104 61
rect 89 21 91 59
rect 100 58 104 59
rect 112 61 116 62
rect 112 59 113 61
rect 115 59 116 61
rect 112 58 116 59
rect 129 52 131 79
rect 148 79 149 81
rect 151 79 152 81
rect 148 71 152 79
rect 148 69 149 71
rect 151 69 152 71
rect 148 68 152 69
rect 158 81 164 82
rect 158 79 161 81
rect 163 79 164 81
rect 158 78 164 79
rect 172 81 176 88
rect 172 79 173 81
rect 175 79 176 81
rect 158 72 162 78
rect 158 71 164 72
rect 158 69 161 71
rect 163 69 164 71
rect 158 68 164 69
rect 172 71 176 79
rect 172 69 173 71
rect 175 69 176 71
rect 158 62 162 68
rect 158 61 164 62
rect 138 59 142 60
rect 138 57 139 59
rect 141 57 142 59
rect 138 56 142 57
rect 158 59 161 61
rect 163 59 164 61
rect 158 58 164 59
rect 172 61 176 69
rect 172 59 173 61
rect 175 59 176 61
rect 172 58 176 59
rect 98 51 102 52
rect 128 51 132 52
rect 98 49 99 51
rect 101 49 129 51
rect 131 49 132 51
rect 98 48 102 49
rect 128 48 132 49
rect 118 41 122 42
rect 109 39 119 41
rect 121 39 122 41
rect 98 33 102 34
rect 109 33 111 39
rect 118 38 122 39
rect 98 31 99 33
rect 101 31 111 33
rect 129 32 131 48
rect 139 42 141 56
rect 138 41 142 42
rect 138 39 139 41
rect 141 39 142 41
rect 138 38 142 39
rect 148 41 152 42
rect 148 39 149 41
rect 151 39 152 41
rect 148 38 152 39
rect 139 32 141 38
rect 128 31 132 32
rect 98 30 102 31
rect 128 29 129 31
rect 131 29 132 31
rect 128 28 132 29
rect 138 31 142 32
rect 138 29 139 31
rect 141 29 142 31
rect 138 28 142 29
rect 100 23 104 24
rect 100 21 101 23
rect 103 21 104 23
rect 149 21 151 38
rect 89 19 151 21
rect 158 22 162 58
rect 158 21 164 22
rect 158 19 161 21
rect 163 19 164 21
rect 158 18 164 19
rect 172 21 176 22
rect 172 19 173 21
rect 175 19 176 21
rect 172 12 176 19
rect -2 11 182 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 77 11
rect 79 9 125 11
rect 127 9 149 11
rect 151 9 173 11
rect 175 9 182 11
rect -2 7 182 9
rect -2 5 41 7
rect 43 5 53 7
rect 55 5 65 7
rect 67 5 89 7
rect 91 5 101 7
rect 103 5 113 7
rect 115 5 182 7
rect -2 0 182 5
<< ptie >>
rect 39 7 69 9
rect 87 7 117 9
rect 39 5 41 7
rect 43 5 53 7
rect 55 5 65 7
rect 67 5 69 7
rect 39 3 69 5
rect 87 5 89 7
rect 91 5 101 7
rect 103 5 113 7
rect 115 5 117 7
rect 87 3 117 5
<< ntie >>
rect 63 95 69 97
rect 63 93 65 95
rect 67 93 69 95
rect 87 95 117 97
rect 87 93 89 95
rect 91 93 101 95
rect 103 93 113 95
rect 115 93 117 95
rect 135 95 141 97
rect 135 93 137 95
rect 139 93 141 95
rect 63 85 69 93
rect 87 91 117 93
rect 135 85 141 93
<< nmos >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 15 37 25
rect 47 15 49 29
rect 71 17 73 25
rect 83 15 85 25
rect 95 15 97 27
rect 107 15 109 27
rect 119 15 121 25
rect 131 17 133 25
rect 155 5 157 25
rect 167 5 169 25
<< pmos >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 65 37 83
rect 47 65 49 83
rect 71 55 73 71
rect 83 55 85 77
rect 95 55 97 77
rect 107 55 109 77
rect 119 55 121 77
rect 131 55 133 77
rect 155 55 157 95
rect 167 55 169 95
<< polyct1 >>
rect 49 59 51 61
rect 31 49 33 51
rect 79 49 81 51
rect 99 49 101 51
rect 39 39 41 41
rect 49 39 51 41
rect 129 49 131 51
rect 65 39 67 41
rect 31 29 33 31
rect 99 31 101 33
rect 79 29 81 31
rect 119 39 121 41
rect 139 39 141 41
rect 149 39 151 41
rect 129 29 131 31
<< ndifct1 >>
rect 5 19 7 21
rect 5 9 7 11
rect 17 19 19 21
rect 53 19 55 21
rect 65 19 67 21
rect 101 21 103 23
rect 139 29 141 31
rect 29 9 31 11
rect 77 9 79 11
rect 125 9 127 11
rect 149 9 151 11
rect 161 19 163 21
rect 173 19 175 21
rect 173 9 175 11
<< ntiect1 >>
rect 65 93 67 95
rect 89 93 91 95
rect 101 93 103 95
rect 113 93 115 95
rect 137 93 139 95
<< ptiect1 >>
rect 41 5 43 7
rect 53 5 55 7
rect 65 5 67 7
rect 89 5 91 7
rect 101 5 103 7
rect 113 5 115 7
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 5 69 7 71
rect 5 59 7 61
rect 17 79 19 81
rect 17 69 19 71
rect 17 59 19 61
rect 29 89 31 91
rect 53 89 55 91
rect 77 89 79 91
rect 41 69 43 71
rect 125 89 127 91
rect 149 89 151 91
rect 149 79 151 81
rect 65 59 67 61
rect 89 69 91 71
rect 101 59 103 61
rect 113 69 115 71
rect 113 59 115 61
rect 149 69 151 71
rect 139 57 141 59
rect 161 79 163 81
rect 161 69 163 71
rect 161 59 163 61
rect 173 89 175 91
rect 173 79 175 81
rect 173 69 175 71
rect 173 59 175 61
<< labels >>
rlabel alu1 30 50 30 50 6 a
rlabel alu1 20 50 20 50 6 cout
rlabel ptiect1 90 6 90 6 6 vss
rlabel alu1 80 45 80 45 6 b
rlabel ntiect1 90 94 90 94 6 vdd
rlabel alu1 160 50 160 50 6 sout
<< end >>
