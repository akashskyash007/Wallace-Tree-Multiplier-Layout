magic
tech scmos
timestamp 1199203346
<< ab >>
rect 0 0 24 72
<< nwell >>
rect -5 32 29 77
<< pwell >>
rect -5 -5 29 32
<< poly >>
rect 12 57 14 61
rect 12 34 14 38
rect 4 32 14 34
rect 4 30 6 32
rect 8 30 14 32
rect 4 28 14 30
rect 12 25 14 28
rect 12 11 14 15
<< ndif >>
rect 3 23 12 25
rect 3 21 6 23
rect 8 21 12 23
rect 3 15 12 21
rect 14 23 22 25
rect 14 21 18 23
rect 20 21 22 23
rect 14 15 22 21
rect 3 13 6 15
rect 8 13 10 15
rect 3 7 10 13
rect 3 5 6 7
rect 8 5 10 7
rect 3 3 10 5
<< pdif >>
rect 3 65 10 68
rect 3 63 6 65
rect 8 63 10 65
rect 3 58 10 63
rect 3 56 6 58
rect 8 57 10 58
rect 8 56 12 57
rect 3 51 12 56
rect 3 49 6 51
rect 8 49 12 51
rect 3 38 12 49
rect 14 49 22 57
rect 14 47 18 49
rect 20 47 22 49
rect 14 42 22 47
rect 14 40 18 42
rect 20 40 22 42
rect 14 38 22 40
<< alu1 >>
rect -2 67 26 72
rect -2 65 17 67
rect 19 65 26 67
rect -2 64 6 65
rect 8 64 26 65
rect 17 49 22 59
rect 17 47 18 49
rect 20 47 22 49
rect 17 43 22 47
rect 2 42 22 43
rect 2 40 18 42
rect 20 40 22 42
rect 2 37 22 40
rect 17 23 22 37
rect 17 21 18 23
rect 20 21 22 23
rect 17 13 22 21
rect -2 7 26 8
rect -2 5 6 7
rect 8 5 17 7
rect 19 5 26 7
rect -2 0 26 5
<< ptie >>
rect 15 7 21 9
rect 15 5 17 7
rect 19 5 21 7
rect 15 3 21 5
<< ntie >>
rect 15 67 21 69
rect 15 65 17 67
rect 19 65 21 67
rect 15 63 21 65
<< nmos >>
rect 12 15 14 25
<< pmos >>
rect 12 38 14 57
<< polyct0 >>
rect 6 30 8 32
<< ndifct0 >>
rect 6 21 8 23
rect 6 13 8 15
<< ndifct1 >>
rect 18 21 20 23
rect 6 5 8 7
<< ntiect1 >>
rect 17 65 19 67
<< ptiect1 >>
rect 17 5 19 7
<< pdifct0 >>
rect 6 63 8 64
rect 6 56 8 58
rect 6 49 8 51
<< pdifct1 >>
rect 6 64 8 65
rect 18 47 20 49
rect 18 40 20 42
<< alu0 >>
rect 5 63 6 64
rect 8 63 9 64
rect 5 58 9 63
rect 5 56 6 58
rect 8 56 9 58
rect 5 51 9 56
rect 5 49 6 51
rect 8 49 9 51
rect 5 47 9 49
rect 4 32 10 33
rect 4 30 6 32
rect 8 30 10 32
rect 4 23 10 30
rect 4 21 6 23
rect 8 21 10 23
rect 4 15 10 21
rect 4 13 6 15
rect 8 13 10 15
rect 4 8 10 13
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 4 12 4 6 vss
rlabel alu1 12 40 12 40 6 z
rlabel alu1 12 68 12 68 6 vdd
rlabel alu1 20 36 20 36 6 z
<< end >>
