magic
tech scmos
timestamp 1199541846
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 59 94 61 98
rect 11 53 13 56
rect 11 51 19 53
rect 11 49 15 51
rect 17 49 19 51
rect 11 47 19 49
rect 23 43 25 55
rect 35 43 37 55
rect 47 43 49 55
rect 59 43 61 55
rect 3 41 61 43
rect 3 39 5 41
rect 7 39 61 41
rect 3 37 61 39
rect 11 31 19 33
rect 11 29 15 31
rect 17 29 19 31
rect 11 27 19 29
rect 11 24 13 27
rect 23 25 25 37
rect 35 25 37 37
rect 47 25 49 37
rect 59 25 61 37
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
rect 59 2 61 6
<< ndif >>
rect 18 24 23 25
rect 3 21 11 24
rect 3 19 5 21
rect 7 19 11 21
rect 3 6 11 19
rect 13 11 23 24
rect 13 9 17 11
rect 19 9 23 11
rect 13 6 23 9
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 6 35 19
rect 37 21 47 25
rect 37 19 41 21
rect 43 19 47 21
rect 37 11 47 19
rect 37 9 41 11
rect 43 9 47 11
rect 37 6 47 9
rect 49 21 59 25
rect 49 19 53 21
rect 55 19 59 21
rect 49 6 59 19
rect 61 21 69 25
rect 61 19 65 21
rect 67 19 69 21
rect 61 11 69 19
rect 61 9 65 11
rect 67 9 69 11
rect 61 6 69 9
<< pdif >>
rect 3 81 11 94
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 56 11 59
rect 13 91 23 94
rect 13 89 17 91
rect 19 89 23 91
rect 13 56 23 89
rect 18 55 23 56
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 91 47 94
rect 37 89 41 91
rect 43 89 47 91
rect 37 81 47 89
rect 37 79 41 81
rect 43 79 47 81
rect 37 71 47 79
rect 37 69 41 71
rect 43 69 47 71
rect 37 61 47 69
rect 37 59 41 61
rect 43 59 47 61
rect 37 55 47 59
rect 49 81 59 94
rect 49 79 53 81
rect 55 79 59 81
rect 49 71 59 79
rect 49 69 53 71
rect 55 69 59 71
rect 49 61 59 69
rect 49 59 53 61
rect 55 59 59 61
rect 49 55 59 59
rect 61 91 69 94
rect 61 89 65 91
rect 67 89 69 91
rect 61 81 69 89
rect 61 79 65 81
rect 67 79 69 81
rect 61 77 69 79
rect 61 55 66 77
<< alu1 >>
rect -2 91 82 100
rect -2 89 17 91
rect 19 89 41 91
rect 43 89 65 91
rect 67 89 82 91
rect -2 88 82 89
rect 4 81 8 83
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 4 59 5 61
rect 7 59 8 61
rect 4 41 8 59
rect 18 52 22 83
rect 13 51 22 52
rect 13 49 15 51
rect 17 49 22 51
rect 13 48 22 49
rect 4 39 5 41
rect 7 39 8 41
rect 4 21 8 39
rect 18 32 22 48
rect 13 31 22 32
rect 13 29 15 31
rect 17 29 22 31
rect 13 28 22 29
rect 4 19 5 21
rect 7 19 8 21
rect 4 17 8 19
rect 18 17 22 28
rect 28 81 32 83
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 28 42 32 59
rect 40 81 44 88
rect 40 79 41 81
rect 43 79 44 81
rect 40 71 44 79
rect 40 69 41 71
rect 43 69 44 71
rect 40 61 44 69
rect 40 59 41 61
rect 43 59 44 61
rect 40 57 44 59
rect 52 81 56 83
rect 52 79 53 81
rect 55 79 56 81
rect 52 71 56 79
rect 52 69 53 71
rect 55 69 56 71
rect 52 61 56 69
rect 64 81 68 88
rect 64 79 65 81
rect 67 79 68 81
rect 64 70 68 79
rect 72 70 76 71
rect 64 69 76 70
rect 64 67 73 69
rect 75 67 76 69
rect 64 66 76 67
rect 52 59 53 61
rect 55 59 56 61
rect 52 42 56 59
rect 72 59 76 66
rect 72 57 73 59
rect 75 57 76 59
rect 72 55 76 57
rect 28 38 56 42
rect 28 21 32 38
rect 28 19 29 21
rect 31 19 32 21
rect 28 17 32 19
rect 40 21 44 23
rect 40 19 41 21
rect 43 19 44 21
rect 40 12 44 19
rect 52 21 56 38
rect 52 19 53 21
rect 55 19 56 21
rect 52 17 56 19
rect 64 36 68 37
rect 64 35 77 36
rect 64 33 65 35
rect 67 33 73 35
rect 75 33 77 35
rect 64 32 77 33
rect 64 21 68 32
rect 64 19 65 21
rect 67 19 68 21
rect 64 12 68 19
rect -2 11 82 12
rect -2 9 17 11
rect 19 9 41 11
rect 43 9 65 11
rect 67 9 82 11
rect -2 0 82 9
<< ptie >>
rect 63 35 77 37
rect 63 33 65 35
rect 67 33 73 35
rect 75 33 77 35
rect 63 31 77 33
<< ntie >>
rect 71 69 77 71
rect 71 67 73 69
rect 75 67 77 69
rect 71 59 77 67
rect 71 57 73 59
rect 75 57 77 59
rect 71 55 77 57
<< nmos >>
rect 11 6 13 24
rect 23 6 25 25
rect 35 6 37 25
rect 47 6 49 25
rect 59 6 61 25
<< pmos >>
rect 11 56 13 94
rect 23 55 25 94
rect 35 55 37 94
rect 47 55 49 94
rect 59 55 61 94
<< polyct1 >>
rect 15 49 17 51
rect 5 39 7 41
rect 15 29 17 31
<< ndifct1 >>
rect 5 19 7 21
rect 17 9 19 11
rect 29 19 31 21
rect 41 19 43 21
rect 41 9 43 11
rect 53 19 55 21
rect 65 19 67 21
rect 65 9 67 11
<< ntiect1 >>
rect 73 67 75 69
rect 73 57 75 59
<< ptiect1 >>
rect 65 33 67 35
rect 73 33 75 35
<< pdifct1 >>
rect 5 79 7 81
rect 5 69 7 71
rect 5 59 7 61
rect 17 89 19 91
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
rect 41 89 43 91
rect 41 79 43 81
rect 41 69 43 71
rect 41 59 43 61
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
rect 65 89 67 91
rect 65 79 67 81
<< labels >>
rlabel alu1 30 50 30 50 6 q
rlabel alu1 20 50 20 50 6 i
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 40 40 40 40 6 q
rlabel alu1 50 40 50 40 6 q
rlabel alu1 40 94 40 94 6 vdd
<< end >>
