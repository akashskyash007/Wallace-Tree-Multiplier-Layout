magic
tech scmos
timestamp 1199201925
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 58 11 63
rect 19 58 21 63
rect 30 59 32 64
rect 40 59 42 64
rect 9 33 11 50
rect 19 47 21 50
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 19 41 25 43
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 9 27 15 29
rect 12 24 14 27
rect 19 24 21 41
rect 30 33 32 50
rect 40 47 42 50
rect 39 45 47 47
rect 39 43 43 45
rect 45 43 47 45
rect 39 41 47 43
rect 25 31 34 33
rect 25 29 27 31
rect 29 29 34 31
rect 25 27 34 29
rect 32 24 34 27
rect 39 24 41 41
rect 12 12 14 17
rect 19 12 21 17
rect 32 12 34 17
rect 39 12 41 17
<< ndif >>
rect 5 22 12 24
rect 5 20 7 22
rect 9 20 12 22
rect 5 17 12 20
rect 14 17 19 24
rect 21 21 32 24
rect 21 19 27 21
rect 29 19 32 21
rect 21 17 32 19
rect 34 17 39 24
rect 41 22 48 24
rect 41 20 44 22
rect 46 20 48 22
rect 41 17 48 20
<< pdif >>
rect 23 58 30 59
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 50 9 54
rect 11 54 19 58
rect 11 52 14 54
rect 16 52 19 54
rect 11 50 19 52
rect 21 56 30 58
rect 21 54 25 56
rect 27 54 30 56
rect 21 50 30 54
rect 32 54 40 59
rect 32 52 35 54
rect 37 52 40 54
rect 32 50 40 52
rect 42 56 50 59
rect 42 54 46 56
rect 48 54 50 56
rect 42 50 50 54
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 10 54 17 56
rect 10 52 14 54
rect 16 52 17 54
rect 10 50 17 52
rect 10 47 14 50
rect 2 43 14 47
rect 2 23 6 43
rect 41 45 54 47
rect 41 43 43 45
rect 45 43 54 45
rect 41 42 54 43
rect 10 31 14 39
rect 26 31 30 39
rect 10 29 11 31
rect 13 29 22 31
rect 10 27 22 29
rect 2 22 14 23
rect 2 20 7 22
rect 9 20 14 22
rect 2 17 14 20
rect 18 17 22 27
rect 26 29 27 31
rect 29 29 38 31
rect 26 25 38 29
rect 50 25 54 42
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 12 17 14 24
rect 19 17 21 24
rect 32 17 34 24
rect 39 17 41 24
<< pmos >>
rect 9 50 11 58
rect 19 50 21 58
rect 30 50 32 59
rect 40 50 42 59
<< polyct0 >>
rect 21 43 23 45
<< polyct1 >>
rect 11 29 13 31
rect 43 43 45 45
rect 27 29 29 31
<< ndifct0 >>
rect 27 19 29 21
rect 44 20 46 22
<< ndifct1 >>
rect 7 20 9 22
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 54 6 56
rect 25 54 27 56
rect 35 52 37 54
rect 46 54 48 56
<< pdifct1 >>
rect 14 52 16 54
<< alu0 >>
rect 3 56 7 68
rect 24 56 28 68
rect 45 56 49 68
rect 3 54 4 56
rect 6 54 7 56
rect 3 52 7 54
rect 24 54 25 56
rect 27 54 28 56
rect 24 52 28 54
rect 34 54 38 56
rect 34 52 35 54
rect 37 52 38 54
rect 45 54 46 56
rect 48 54 49 56
rect 45 52 49 54
rect 34 46 38 52
rect 19 45 38 46
rect 19 43 21 45
rect 23 43 38 45
rect 19 42 38 43
rect 34 38 38 42
rect 34 34 47 38
rect 43 22 47 34
rect 25 21 31 22
rect 25 19 27 21
rect 29 19 31 21
rect 25 12 31 19
rect 43 20 44 22
rect 46 20 47 22
rect 43 18 47 20
<< labels >>
rlabel alu0 28 44 28 44 6 an
rlabel alu0 45 28 45 28 6 an
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 36 12 36 6 b
rlabel alu1 20 24 20 24 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 32 28 32 6 a1
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 52 36 52 36 6 a2
rlabel polyct1 44 44 44 44 6 a2
<< end >>
