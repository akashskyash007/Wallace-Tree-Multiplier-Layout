magic
tech scmos
timestamp 1199542146
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -5 48 95 105
<< pwell >>
rect -5 -5 95 48
<< poly >>
rect 75 94 77 98
rect 11 85 13 89
rect 23 85 25 89
rect 31 85 33 89
rect 47 85 49 89
rect 55 85 57 89
rect 11 41 13 65
rect 23 63 25 66
rect 17 61 25 63
rect 17 59 19 61
rect 21 59 23 61
rect 17 57 23 59
rect 31 43 33 66
rect 47 57 49 66
rect 55 63 57 66
rect 55 61 63 63
rect 57 59 59 61
rect 61 59 63 61
rect 57 57 63 59
rect 47 55 53 57
rect 47 53 49 55
rect 51 53 53 55
rect 47 51 53 53
rect 37 49 43 51
rect 37 47 39 49
rect 41 47 43 49
rect 75 47 77 55
rect 37 45 77 47
rect 27 41 33 43
rect 11 39 29 41
rect 31 39 49 41
rect 11 15 13 39
rect 27 37 33 39
rect 17 31 23 33
rect 17 29 19 31
rect 21 29 23 31
rect 17 27 25 29
rect 23 14 25 27
rect 29 21 35 23
rect 29 19 31 21
rect 33 19 35 21
rect 29 17 35 19
rect 31 14 33 17
rect 47 15 49 39
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 55 27 63 29
rect 55 15 57 27
rect 75 25 77 45
rect 11 2 13 6
rect 23 2 25 6
rect 31 2 33 6
rect 47 2 49 6
rect 55 2 57 6
rect 75 2 77 6
<< ndif >>
rect 3 21 9 25
rect 3 19 5 21
rect 7 19 9 21
rect 3 15 9 19
rect 37 31 45 33
rect 37 29 39 31
rect 41 29 45 31
rect 3 6 11 15
rect 13 14 18 15
rect 37 15 45 29
rect 59 21 75 25
rect 59 19 69 21
rect 71 19 75 21
rect 59 15 75 19
rect 37 14 47 15
rect 13 11 23 14
rect 13 9 17 11
rect 19 9 23 11
rect 13 6 23 9
rect 25 6 31 14
rect 33 6 47 14
rect 49 6 55 15
rect 57 11 75 15
rect 57 9 69 11
rect 71 9 75 11
rect 57 6 75 9
rect 77 21 85 25
rect 77 19 81 21
rect 83 19 85 21
rect 77 6 85 19
<< pdif >>
rect 15 91 21 93
rect 59 91 75 94
rect 15 89 17 91
rect 19 89 21 91
rect 59 89 69 91
rect 71 89 75 91
rect 15 85 21 89
rect 59 85 75 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 66 23 85
rect 25 66 31 85
rect 33 81 47 85
rect 33 79 39 81
rect 41 79 47 81
rect 33 71 47 79
rect 33 69 39 71
rect 41 69 47 71
rect 33 66 47 69
rect 49 66 55 85
rect 57 81 75 85
rect 57 79 69 81
rect 71 79 75 81
rect 57 71 75 79
rect 57 69 69 71
rect 71 69 75 71
rect 57 66 75 69
rect 13 65 18 66
rect 59 65 75 66
rect 67 61 75 65
rect 67 59 69 61
rect 71 59 75 61
rect 67 55 75 59
rect 77 81 85 94
rect 77 79 81 81
rect 83 79 85 81
rect 77 71 85 79
rect 77 69 81 71
rect 83 69 85 71
rect 77 61 85 69
rect 77 59 81 61
rect 83 59 85 61
rect 77 55 85 59
<< alu1 >>
rect -2 95 92 100
rect -2 93 29 95
rect 31 93 39 95
rect 41 93 49 95
rect 51 93 92 95
rect -2 91 92 93
rect -2 89 17 91
rect 19 89 69 91
rect 71 89 92 91
rect -2 88 92 89
rect 4 81 8 83
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 4 69 5 71
rect 7 69 8 71
rect 4 22 8 69
rect 18 61 22 83
rect 18 59 19 61
rect 21 59 22 61
rect 18 31 22 59
rect 18 29 19 31
rect 21 29 22 31
rect 18 27 22 29
rect 28 41 32 83
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 81 42 83
rect 38 79 39 81
rect 41 79 42 81
rect 38 71 42 79
rect 38 69 39 71
rect 41 69 42 71
rect 38 49 42 69
rect 58 61 62 83
rect 58 59 59 61
rect 61 59 62 61
rect 38 47 39 49
rect 41 47 42 49
rect 38 31 42 47
rect 38 29 39 31
rect 41 29 42 31
rect 38 27 42 29
rect 48 55 52 57
rect 48 53 49 55
rect 51 53 52 55
rect 48 22 52 53
rect 4 21 52 22
rect 4 19 5 21
rect 7 19 31 21
rect 33 19 52 21
rect 4 18 52 19
rect 58 31 62 59
rect 68 81 72 88
rect 68 79 69 81
rect 71 79 72 81
rect 68 71 72 79
rect 68 69 69 71
rect 71 69 72 71
rect 68 61 72 69
rect 68 59 69 61
rect 71 59 72 61
rect 68 57 72 59
rect 78 82 82 83
rect 78 81 85 82
rect 78 79 81 81
rect 83 79 85 81
rect 78 78 85 79
rect 78 72 82 78
rect 78 71 85 72
rect 78 69 81 71
rect 83 69 85 71
rect 78 68 85 69
rect 78 62 82 68
rect 78 61 85 62
rect 78 59 81 61
rect 83 59 85 61
rect 78 58 85 59
rect 58 29 59 31
rect 61 29 62 31
rect 4 17 8 18
rect 58 17 62 29
rect 68 21 72 23
rect 68 19 69 21
rect 71 19 72 21
rect 68 12 72 19
rect 78 22 82 58
rect 78 21 85 22
rect 78 19 81 21
rect 83 19 85 21
rect 78 18 85 19
rect 78 17 82 18
rect -2 11 92 12
rect -2 9 17 11
rect 19 9 69 11
rect 71 9 92 11
rect -2 0 92 9
<< ntie >>
rect 27 95 53 97
rect 27 93 29 95
rect 31 93 39 95
rect 41 93 49 95
rect 51 93 53 95
rect 27 91 53 93
<< nmos >>
rect 11 6 13 15
rect 23 6 25 14
rect 31 6 33 14
rect 47 6 49 15
rect 55 6 57 15
rect 75 6 77 25
<< pmos >>
rect 11 65 13 85
rect 23 66 25 85
rect 31 66 33 85
rect 47 66 49 85
rect 55 66 57 85
rect 75 55 77 94
<< polyct1 >>
rect 19 59 21 61
rect 59 59 61 61
rect 49 53 51 55
rect 39 47 41 49
rect 29 39 31 41
rect 19 29 21 31
rect 31 19 33 21
rect 59 29 61 31
<< ndifct1 >>
rect 5 19 7 21
rect 39 29 41 31
rect 69 19 71 21
rect 17 9 19 11
rect 69 9 71 11
rect 81 19 83 21
<< ntiect1 >>
rect 29 93 31 95
rect 39 93 41 95
rect 49 93 51 95
<< pdifct1 >>
rect 17 89 19 91
rect 69 89 71 91
rect 5 79 7 81
rect 5 69 7 71
rect 39 79 41 81
rect 39 69 41 71
rect 69 79 71 81
rect 69 69 71 71
rect 69 59 71 61
rect 81 79 83 81
rect 81 69 83 71
rect 81 59 83 61
<< labels >>
rlabel alu1 20 55 20 55 6 i0
rlabel alu1 30 55 30 55 6 cmd
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 60 50 60 50 6 i1
rlabel alu1 45 94 45 94 6 vdd
rlabel alu1 80 50 80 50 6 q
<< end >>
