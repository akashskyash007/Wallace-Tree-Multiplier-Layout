magic
tech scmos
timestamp 1199202125
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 12 65 14 70
rect 22 65 24 70
rect 29 65 31 70
rect 39 65 41 70
rect 49 65 51 70
rect 59 65 61 70
rect 12 35 14 38
rect 22 35 24 38
rect 9 33 24 35
rect 9 31 11 33
rect 13 31 24 33
rect 29 32 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 9 29 24 31
rect 28 29 31 32
rect 35 33 41 35
rect 35 31 37 33
rect 39 31 41 33
rect 35 29 41 31
rect 48 33 55 35
rect 48 31 51 33
rect 53 31 55 33
rect 48 29 55 31
rect 59 33 65 35
rect 59 31 61 33
rect 63 31 65 33
rect 59 29 65 31
rect 9 24 11 29
rect 21 26 23 29
rect 28 26 30 29
rect 38 26 40 29
rect 48 26 50 29
rect 59 26 61 29
rect 9 7 11 12
rect 21 9 23 14
rect 28 5 30 14
rect 38 9 40 14
rect 48 5 50 14
rect 59 9 61 14
rect 28 3 50 5
<< ndif >>
rect 13 24 21 26
rect 4 18 9 24
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 14 21 24
rect 23 14 28 26
rect 30 24 38 26
rect 30 22 33 24
rect 35 22 38 24
rect 30 14 38 22
rect 40 18 48 26
rect 40 16 43 18
rect 45 16 48 18
rect 40 14 48 16
rect 50 18 59 26
rect 50 16 53 18
rect 55 16 59 18
rect 50 14 59 16
rect 61 24 68 26
rect 61 22 64 24
rect 66 22 68 24
rect 61 20 68 22
rect 61 14 66 20
rect 11 12 19 14
rect 13 7 19 12
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
<< pdif >>
rect 7 59 12 65
rect 5 57 12 59
rect 5 55 7 57
rect 9 55 12 57
rect 5 50 12 55
rect 5 48 7 50
rect 9 48 12 50
rect 5 46 12 48
rect 7 38 12 46
rect 14 63 22 65
rect 14 61 17 63
rect 19 61 22 63
rect 14 56 22 61
rect 14 54 17 56
rect 19 54 22 56
rect 14 38 22 54
rect 24 38 29 65
rect 31 49 39 65
rect 31 47 34 49
rect 36 47 39 49
rect 31 42 39 47
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 58 49 65
rect 41 56 44 58
rect 46 56 49 58
rect 41 38 49 56
rect 51 63 59 65
rect 51 61 54 63
rect 56 61 59 63
rect 51 56 59 61
rect 51 54 54 56
rect 56 54 59 56
rect 51 38 59 54
rect 61 57 66 65
rect 61 55 68 57
rect 61 53 64 55
rect 66 53 68 55
rect 61 48 68 53
rect 61 46 64 48
rect 66 46 68 48
rect 61 44 68 46
rect 61 38 66 44
<< alu1 >>
rect -2 64 74 72
rect 33 49 38 51
rect 33 47 34 49
rect 36 47 38 49
rect 2 35 6 43
rect 33 42 38 47
rect 18 40 34 42
rect 36 40 38 42
rect 18 38 38 40
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 18 26 22 38
rect 33 33 47 34
rect 33 31 37 33
rect 39 31 47 33
rect 33 30 47 31
rect 18 24 37 26
rect 18 22 33 24
rect 35 22 37 24
rect 41 22 47 30
rect 57 35 63 42
rect 57 33 70 35
rect 57 31 61 33
rect 63 31 70 33
rect 57 29 70 31
rect 18 21 37 22
rect -2 7 74 8
rect -2 5 15 7
rect 17 5 74 7
rect -2 0 74 5
<< nmos >>
rect 9 12 11 24
rect 21 14 23 26
rect 28 14 30 26
rect 38 14 40 26
rect 48 14 50 26
rect 59 14 61 26
<< pmos >>
rect 12 38 14 65
rect 22 38 24 65
rect 29 38 31 65
rect 39 38 41 65
rect 49 38 51 65
rect 59 38 61 65
<< polyct0 >>
rect 51 31 53 33
<< polyct1 >>
rect 11 31 13 33
rect 37 31 39 33
rect 61 31 63 33
<< ndifct0 >>
rect 4 14 6 16
rect 43 16 45 18
rect 53 16 55 18
rect 64 22 66 24
<< ndifct1 >>
rect 33 22 35 24
rect 15 5 17 7
<< pdifct0 >>
rect 7 55 9 57
rect 7 48 9 50
rect 17 61 19 63
rect 17 54 19 56
rect 44 56 46 58
rect 54 61 56 63
rect 54 54 56 56
rect 64 53 66 55
rect 64 46 66 48
<< pdifct1 >>
rect 34 47 36 49
rect 34 40 36 42
<< alu0 >>
rect 15 63 21 64
rect 15 61 17 63
rect 19 61 21 63
rect 6 57 10 59
rect 6 55 7 57
rect 9 55 10 57
rect 6 50 10 55
rect 15 56 21 61
rect 53 63 57 64
rect 53 61 54 63
rect 56 61 57 63
rect 15 54 17 56
rect 19 54 21 56
rect 15 53 21 54
rect 24 58 48 59
rect 24 56 44 58
rect 46 56 48 58
rect 24 55 48 56
rect 53 56 57 61
rect 24 50 28 55
rect 53 54 54 56
rect 56 54 57 56
rect 53 52 57 54
rect 62 55 68 56
rect 62 53 64 55
rect 66 53 68 55
rect 6 48 7 50
rect 9 48 28 50
rect 6 46 28 48
rect 62 49 68 53
rect 50 48 68 49
rect 50 46 64 48
rect 66 46 68 48
rect 50 45 68 46
rect 50 33 54 45
rect 50 31 51 33
rect 53 31 54 33
rect 50 26 54 31
rect 50 24 68 26
rect 50 22 64 24
rect 66 22 68 24
rect 62 21 68 22
rect 41 18 47 19
rect 41 17 43 18
rect 2 16 43 17
rect 45 16 47 18
rect 2 14 4 16
rect 6 14 47 16
rect 2 13 47 14
rect 51 18 57 19
rect 51 16 53 18
rect 55 16 57 18
rect 51 8 57 16
<< labels >>
rlabel alu0 8 52 8 52 6 n1
rlabel alu0 24 15 24 15 6 n3
rlabel alu0 44 16 44 16 6 n3
rlabel alu0 36 57 36 57 6 n1
rlabel ndifct0 65 23 65 23 6 bn
rlabel alu0 52 35 52 35 6 bn
rlabel alu0 59 47 59 47 6 bn
rlabel alu0 65 50 65 50 6 bn
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 4 36 4 36 6 a
rlabel alu1 20 28 20 28 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 36 32 36 32 6 c
rlabel alu1 44 28 44 28 6 c
rlabel alu1 36 48 36 48 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 68 32 68 32 6 b
rlabel alu1 60 36 60 36 6 b
<< end >>
