magic
tech scmos
timestamp 1199202734
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 69 41 74
rect 49 69 51 74
rect 59 69 61 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 33 39
rect 19 35 27 37
rect 29 35 33 37
rect 19 33 33 35
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 37 51 39
rect 38 35 43 37
rect 45 35 51 37
rect 38 33 51 35
rect 55 37 61 39
rect 55 35 57 37
rect 59 35 61 37
rect 55 33 61 35
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 12 15 14 19
rect 19 14 21 19
rect 31 6 33 10
rect 38 6 40 10
rect 48 6 50 10
rect 55 6 57 10
<< ndif >>
rect 5 28 12 30
rect 5 26 7 28
rect 9 26 12 28
rect 5 24 12 26
rect 7 19 12 24
rect 14 19 19 30
rect 21 19 31 30
rect 23 14 31 19
rect 23 12 25 14
rect 27 12 31 14
rect 23 10 31 12
rect 33 10 38 30
rect 40 21 48 30
rect 40 19 43 21
rect 45 19 48 21
rect 40 10 48 19
rect 50 10 55 30
rect 57 11 66 30
rect 57 10 61 11
rect 59 9 61 10
rect 63 9 66 11
rect 59 7 66 9
<< pdif >>
rect 2 67 9 69
rect 2 65 4 67
rect 6 65 9 67
rect 2 60 9 65
rect 2 58 4 60
rect 6 58 9 60
rect 2 42 9 58
rect 11 61 19 69
rect 11 59 14 61
rect 16 59 19 61
rect 11 53 19 59
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 61 39 69
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 67 49 69
rect 41 65 44 67
rect 46 65 49 67
rect 41 60 49 65
rect 41 58 44 60
rect 46 58 49 60
rect 41 42 49 58
rect 51 61 59 69
rect 51 59 54 61
rect 56 59 59 61
rect 51 54 59 59
rect 51 52 54 54
rect 56 52 59 54
rect 51 42 59 52
rect 61 67 68 69
rect 61 65 64 67
rect 66 65 68 67
rect 61 60 68 65
rect 61 58 64 60
rect 66 58 68 60
rect 61 42 68 58
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 2 53 54 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 52 54 53
rect 56 52 63 54
rect 36 51 63 52
rect 2 50 63 51
rect 2 29 6 50
rect 25 42 63 46
rect 10 37 21 39
rect 10 35 11 37
rect 13 35 21 37
rect 10 33 21 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 17 30 21 33
rect 41 30 47 35
rect 2 28 11 29
rect 2 26 7 28
rect 9 26 11 28
rect 17 26 55 30
rect 2 25 11 26
rect 7 22 11 25
rect 7 21 47 22
rect 7 19 43 21
rect 45 19 47 21
rect 7 18 47 19
rect -2 11 74 12
rect -2 9 61 11
rect 63 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 12 19 14 30
rect 19 19 21 30
rect 31 10 33 30
rect 38 10 40 30
rect 48 10 50 30
rect 55 10 57 30
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 49 42 51 69
rect 59 42 61 69
<< polyct0 >>
rect 57 35 59 37
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 43 35 45 37
<< ndifct0 >>
rect 25 12 27 14
<< ndifct1 >>
rect 7 26 9 28
rect 43 19 45 21
rect 61 9 63 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 65 6 67
rect 4 58 6 60
rect 14 59 16 61
rect 24 65 26 67
rect 24 58 26 60
rect 44 65 46 67
rect 44 58 46 60
rect 54 59 56 61
rect 64 65 66 67
rect 64 58 66 60
<< pdifct1 >>
rect 14 51 16 53
rect 34 59 36 61
rect 34 51 36 53
rect 54 52 56 54
<< alu0 >>
rect 2 67 8 68
rect 2 65 4 67
rect 6 65 8 67
rect 2 60 8 65
rect 22 67 28 68
rect 22 65 24 67
rect 26 65 28 67
rect 2 58 4 60
rect 6 58 8 60
rect 2 57 8 58
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 60 28 65
rect 42 67 48 68
rect 42 65 44 67
rect 46 65 48 67
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 42 60 48 65
rect 62 67 68 68
rect 62 65 64 67
rect 66 65 68 67
rect 42 58 44 60
rect 46 58 48 60
rect 42 57 48 58
rect 53 61 57 63
rect 53 59 54 61
rect 56 59 57 61
rect 53 54 57 59
rect 62 60 68 65
rect 62 58 64 60
rect 66 58 68 60
rect 62 57 68 58
rect 55 37 61 42
rect 55 35 57 37
rect 59 35 61 37
rect 55 34 61 35
rect 23 14 29 15
rect 23 12 25 14
rect 27 12 29 14
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 b
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 b
rlabel alu1 28 40 28 40 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel ndifct1 44 20 44 20 6 z
rlabel alu1 52 28 52 28 6 b
rlabel alu1 44 32 44 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 52 44 52 44 6 a
rlabel alu1 52 52 52 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 60 44 60 44 6 a
rlabel alu1 60 52 60 52 6 z
<< end >>
