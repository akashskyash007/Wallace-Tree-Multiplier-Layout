magic
tech scmos
timestamp 1199202798
<< ab >>
rect 0 0 136 80
<< nwell >>
rect -5 36 141 88
<< pwell >>
rect -5 -8 141 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 99 70 101 74
rect 109 70 111 74
rect 119 61 121 65
rect 9 39 11 48
rect 19 47 21 50
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 19 41 25 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 36 15 37
rect 13 35 17 36
rect 9 33 17 35
rect 15 30 17 33
rect 22 30 24 41
rect 29 39 31 50
rect 39 39 41 50
rect 49 47 51 50
rect 45 45 51 47
rect 45 43 47 45
rect 49 43 51 45
rect 45 41 51 43
rect 29 37 41 39
rect 29 35 37 37
rect 39 35 41 37
rect 29 33 41 35
rect 29 30 31 33
rect 39 30 41 33
rect 46 30 48 41
rect 59 35 61 50
rect 69 35 71 50
rect 79 47 81 50
rect 79 45 85 47
rect 79 43 81 45
rect 83 43 85 45
rect 79 41 85 43
rect 53 33 77 35
rect 53 30 55 33
rect 62 29 68 33
rect 75 30 77 33
rect 82 30 84 41
rect 89 39 91 50
rect 99 39 101 50
rect 109 46 111 50
rect 105 44 111 46
rect 105 42 107 44
rect 109 42 111 44
rect 105 40 111 42
rect 89 37 101 39
rect 89 35 92 37
rect 94 35 101 37
rect 89 33 101 35
rect 89 30 91 33
rect 99 30 101 33
rect 106 30 108 40
rect 119 39 121 43
rect 119 37 127 39
rect 119 35 123 37
rect 125 35 127 37
rect 113 33 127 35
rect 113 30 115 33
rect 62 27 64 29
rect 66 27 68 29
rect 62 25 68 27
rect 15 6 17 10
rect 22 6 24 10
rect 29 6 31 10
rect 39 6 41 10
rect 46 6 48 10
rect 53 6 55 10
rect 75 6 77 10
rect 82 6 84 10
rect 89 6 91 10
rect 99 6 101 10
rect 106 6 108 10
rect 113 6 115 10
<< ndif >>
rect 7 14 15 30
rect 7 12 10 14
rect 12 12 15 14
rect 7 10 15 12
rect 17 10 22 30
rect 24 10 29 30
rect 31 21 39 30
rect 31 19 34 21
rect 36 19 39 21
rect 31 10 39 19
rect 41 10 46 30
rect 48 10 53 30
rect 55 22 60 30
rect 70 22 75 30
rect 55 14 75 22
rect 55 12 58 14
rect 60 12 70 14
rect 72 12 75 14
rect 55 10 75 12
rect 77 10 82 30
rect 84 10 89 30
rect 91 21 99 30
rect 91 19 94 21
rect 96 19 99 21
rect 91 10 99 19
rect 101 10 106 30
rect 108 10 113 30
rect 115 21 123 30
rect 115 19 118 21
rect 120 19 123 21
rect 115 14 123 19
rect 115 12 118 14
rect 120 12 123 14
rect 115 10 123 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 48 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 50 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 50 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 50 39 52
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 61 49 66
rect 41 59 44 61
rect 46 59 49 61
rect 41 50 49 59
rect 51 61 59 70
rect 51 59 54 61
rect 56 59 59 61
rect 51 54 59 59
rect 51 52 54 54
rect 56 52 59 54
rect 51 50 59 52
rect 61 68 69 70
rect 61 66 64 68
rect 66 66 69 68
rect 61 61 69 66
rect 61 59 64 61
rect 66 59 69 61
rect 61 50 69 59
rect 71 61 79 70
rect 71 59 74 61
rect 76 59 79 61
rect 71 54 79 59
rect 71 52 74 54
rect 76 52 79 54
rect 71 50 79 52
rect 81 68 89 70
rect 81 66 84 68
rect 86 66 89 68
rect 81 61 89 66
rect 81 59 84 61
rect 86 59 89 61
rect 81 50 89 59
rect 91 61 99 70
rect 91 59 94 61
rect 96 59 99 61
rect 91 54 99 59
rect 91 52 94 54
rect 96 52 99 54
rect 91 50 99 52
rect 101 68 109 70
rect 101 66 104 68
rect 106 66 109 68
rect 101 61 109 66
rect 101 59 104 61
rect 106 59 109 61
rect 101 50 109 59
rect 111 61 116 70
rect 111 57 119 61
rect 111 55 114 57
rect 116 55 119 57
rect 111 50 119 55
rect 11 48 16 50
rect 114 43 119 50
rect 121 59 129 61
rect 121 57 125 59
rect 127 57 129 59
rect 121 52 129 57
rect 121 50 125 52
rect 127 50 129 52
rect 121 43 129 50
<< alu1 >>
rect -2 81 138 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 138 81
rect -2 68 138 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 73 61 78 63
rect 73 59 74 61
rect 76 59 78 61
rect 73 54 78 59
rect 113 57 119 63
rect 113 55 114 57
rect 116 55 119 57
rect 113 54 119 55
rect 2 52 14 54
rect 16 52 34 54
rect 36 52 54 54
rect 56 52 74 54
rect 76 52 94 54
rect 96 52 119 54
rect 2 50 119 52
rect 2 22 6 50
rect 19 45 119 46
rect 19 43 21 45
rect 23 43 47 45
rect 49 43 81 45
rect 83 44 119 45
rect 83 43 107 44
rect 19 42 107 43
rect 109 42 119 44
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 33 37 96 38
rect 33 35 37 37
rect 39 35 92 37
rect 94 35 96 37
rect 33 34 96 35
rect 105 34 111 42
rect 121 37 127 38
rect 121 35 123 37
rect 125 35 127 37
rect 121 30 127 35
rect 10 29 127 30
rect 10 27 64 29
rect 66 27 127 29
rect 10 26 127 27
rect 2 21 103 22
rect 2 19 34 21
rect 36 19 94 21
rect 96 19 103 21
rect 2 18 103 19
rect -2 1 138 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 138 1
rect -2 -2 138 -1
<< ptie >>
rect 0 1 136 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 136 1
rect 0 -3 136 -1
<< ntie >>
rect 0 81 136 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 136 81
rect 0 77 136 79
<< nmos >>
rect 15 10 17 30
rect 22 10 24 30
rect 29 10 31 30
rect 39 10 41 30
rect 46 10 48 30
rect 53 10 55 30
rect 75 10 77 30
rect 82 10 84 30
rect 89 10 91 30
rect 99 10 101 30
rect 106 10 108 30
rect 113 10 115 30
<< pmos >>
rect 9 48 11 70
rect 19 50 21 70
rect 29 50 31 70
rect 39 50 41 70
rect 49 50 51 70
rect 59 50 61 70
rect 69 50 71 70
rect 79 50 81 70
rect 89 50 91 70
rect 99 50 101 70
rect 109 50 111 70
rect 119 43 121 61
<< polyct1 >>
rect 21 43 23 45
rect 11 35 13 37
rect 47 43 49 45
rect 37 35 39 37
rect 81 43 83 45
rect 107 42 109 44
rect 92 35 94 37
rect 123 35 125 37
rect 64 27 66 29
<< ndifct0 >>
rect 10 12 12 14
rect 58 12 60 14
rect 70 12 72 14
rect 118 19 120 21
rect 118 12 120 14
<< ndifct1 >>
rect 34 19 36 21
rect 94 19 96 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 59 16 61
rect 24 66 26 68
rect 24 59 26 61
rect 44 66 46 68
rect 44 59 46 61
rect 54 59 56 61
rect 64 66 66 68
rect 64 59 66 61
rect 84 66 86 68
rect 84 59 86 61
rect 94 59 96 61
rect 104 66 106 68
rect 104 59 106 61
rect 125 57 127 59
rect 125 50 127 52
<< pdifct1 >>
rect 14 52 16 54
rect 34 59 36 61
rect 34 52 36 54
rect 54 52 56 54
rect 74 59 76 61
rect 74 52 76 54
rect 94 52 96 54
rect 114 55 116 57
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 61 28 66
rect 42 66 44 68
rect 46 66 48 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 42 61 48 66
rect 62 66 64 68
rect 66 66 68 68
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 53 61 57 63
rect 53 59 54 61
rect 56 59 57 61
rect 53 54 57 59
rect 62 61 68 66
rect 82 66 84 68
rect 86 66 88 68
rect 62 59 64 61
rect 66 59 68 61
rect 62 58 68 59
rect 82 61 88 66
rect 102 66 104 68
rect 106 66 108 68
rect 82 59 84 61
rect 86 59 88 61
rect 82 58 88 59
rect 93 61 97 63
rect 93 59 94 61
rect 96 59 97 61
rect 93 54 97 59
rect 102 61 108 66
rect 102 59 104 61
rect 106 59 108 61
rect 102 58 108 59
rect 123 59 129 68
rect 123 57 125 59
rect 127 57 129 59
rect 123 52 129 57
rect 123 50 125 52
rect 127 50 129 52
rect 123 49 129 50
rect 116 21 122 22
rect 116 19 118 21
rect 120 19 122 21
rect 8 14 14 15
rect 8 12 10 14
rect 12 12 14 14
rect 56 14 62 15
rect 56 12 58 14
rect 60 12 62 14
rect 68 14 74 15
rect 68 12 70 14
rect 72 12 74 14
rect 116 14 122 19
rect 116 12 118 14
rect 120 12 122 14
<< labels >>
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 44 28 44 6 b
rlabel alu1 44 44 44 44 6 b
rlabel alu1 44 36 44 36 6 c
rlabel alu1 36 44 36 44 6 b
rlabel alu1 36 36 36 36 6 c
rlabel alu1 44 52 44 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 68 6 68 6 6 vss
rlabel alu1 52 20 52 20 6 z
rlabel alu1 52 28 52 28 6 a
rlabel alu1 68 28 68 28 6 a
rlabel alu1 76 28 76 28 6 a
rlabel alu1 76 20 76 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 60 28 60 28 6 a
rlabel alu1 60 20 60 20 6 z
rlabel alu1 52 36 52 36 6 c
rlabel alu1 52 44 52 44 6 b
rlabel alu1 68 44 68 44 6 b
rlabel alu1 76 44 76 44 6 b
rlabel alu1 76 36 76 36 6 c
rlabel alu1 68 36 68 36 6 c
rlabel alu1 60 44 60 44 6 b
rlabel alu1 60 36 60 36 6 c
rlabel alu1 60 52 60 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 76 56 76 56 6 z
rlabel alu1 68 74 68 74 6 vdd
rlabel alu1 84 20 84 20 6 z
rlabel alu1 84 28 84 28 6 a
rlabel alu1 92 28 92 28 6 a
rlabel alu1 108 28 108 28 6 a
rlabel alu1 100 28 100 28 6 a
rlabel alu1 100 20 100 20 6 z
rlabel alu1 92 20 92 20 6 z
rlabel alu1 84 36 84 36 6 c
rlabel alu1 84 44 84 44 6 b
rlabel alu1 92 44 92 44 6 b
rlabel alu1 108 40 108 40 6 b
rlabel alu1 100 44 100 44 6 b
rlabel alu1 92 36 92 36 6 c
rlabel alu1 92 52 92 52 6 z
rlabel alu1 108 52 108 52 6 z
rlabel alu1 100 52 100 52 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 116 28 116 28 6 a
rlabel alu1 124 32 124 32 6 a
rlabel alu1 116 44 116 44 6 b
rlabel alu1 116 56 116 56 6 z
<< end >>
