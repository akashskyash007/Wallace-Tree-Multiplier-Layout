magic
tech scmos
timestamp 1199202091
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 61 31 65
rect 9 38 11 42
rect 19 38 21 42
rect 29 40 31 45
rect 26 38 32 40
rect 9 36 22 38
rect 9 34 18 36
rect 20 34 22 36
rect 26 36 28 38
rect 30 36 32 38
rect 26 34 32 36
rect 9 32 22 34
rect 9 27 11 32
rect 19 27 21 32
rect 29 27 31 34
rect 29 15 31 19
rect 9 8 11 13
rect 19 8 21 13
<< ndif >>
rect 4 19 9 27
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 11 21 19 27
rect 11 19 14 21
rect 16 19 19 21
rect 11 13 19 19
rect 21 23 29 27
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 31 25 38 27
rect 31 23 34 25
rect 36 23 38 25
rect 31 21 38 23
rect 31 19 36 21
rect 21 13 27 19
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 61 27 70
rect 21 56 29 61
rect 21 54 24 56
rect 26 54 29 56
rect 21 45 29 54
rect 31 59 38 61
rect 31 57 34 59
rect 36 57 38 59
rect 31 52 38 57
rect 31 50 34 52
rect 36 50 38 52
rect 31 48 38 50
rect 31 45 36 48
rect 21 42 26 45
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 31 6 50
rect 17 42 31 46
rect 25 38 31 42
rect 25 36 28 38
rect 30 36 31 38
rect 25 34 31 36
rect 2 25 14 31
rect 10 23 14 25
rect 10 21 17 23
rect 10 19 14 21
rect 16 19 17 21
rect 10 17 17 19
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 13 11 27
rect 19 13 21 27
rect 29 19 31 27
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 45 31 61
<< polyct0 >>
rect 18 34 20 36
<< polyct1 >>
rect 28 36 30 38
<< ndifct0 >>
rect 4 15 6 17
rect 24 21 26 23
rect 34 23 36 25
<< ndifct1 >>
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 54 26 56
rect 34 57 36 59
rect 34 50 36 52
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 23 56 27 68
rect 23 54 24 56
rect 26 54 27 56
rect 23 52 27 54
rect 32 59 38 60
rect 32 57 34 59
rect 36 57 38 59
rect 32 52 38 57
rect 32 50 34 52
rect 36 50 38 52
rect 32 49 38 50
rect 17 36 21 38
rect 17 34 18 36
rect 20 34 21 36
rect 17 31 21 34
rect 34 31 38 49
rect 17 27 38 31
rect 33 25 38 27
rect 22 23 28 24
rect 3 17 7 19
rect 22 21 24 23
rect 26 21 28 23
rect 33 23 34 25
rect 36 23 38 25
rect 33 21 38 23
rect 3 15 4 17
rect 6 15 7 17
rect 3 12 7 15
rect 22 12 28 21
<< labels >>
rlabel alu0 19 32 19 32 6 an
rlabel alu0 36 40 36 40 6 an
rlabel alu0 35 54 35 54 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 40 28 40 6 a
rlabel alu1 20 44 20 44 6 a
rlabel alu1 20 74 20 74 6 vdd
<< end >>
