magic
tech scmos
timestamp 1199202106
<< ab >>
rect 0 0 88 72
<< nwell >>
rect -5 32 93 77
<< pwell >>
rect -5 -5 93 32
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 39 65 41 70
rect 46 65 48 70
rect 56 65 58 70
rect 66 65 68 70
rect 76 65 78 70
rect 9 35 11 38
rect 19 35 21 38
rect 39 35 41 38
rect 46 35 48 38
rect 56 35 58 38
rect 66 35 68 38
rect 76 35 78 38
rect 5 33 11 35
rect 5 31 7 33
rect 9 31 11 33
rect 5 29 11 31
rect 17 33 23 35
rect 17 31 19 33
rect 21 31 23 33
rect 17 29 23 31
rect 32 33 42 35
rect 32 31 34 33
rect 36 31 42 33
rect 46 32 49 35
rect 32 29 42 31
rect 9 26 11 29
rect 19 26 21 29
rect 40 26 42 29
rect 47 26 49 32
rect 55 33 61 35
rect 55 31 57 33
rect 59 31 61 33
rect 55 29 61 31
rect 65 33 71 35
rect 65 31 67 33
rect 69 31 71 33
rect 65 29 71 31
rect 76 33 86 35
rect 76 31 82 33
rect 84 31 86 33
rect 76 29 86 31
rect 57 26 59 29
rect 67 26 69 29
rect 77 26 79 29
rect 9 7 11 12
rect 19 7 21 12
rect 40 9 42 14
rect 47 4 49 14
rect 57 8 59 12
rect 67 4 69 12
rect 77 7 79 12
rect 47 2 69 4
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 12 9 15
rect 11 16 19 26
rect 11 14 14 16
rect 16 14 19 16
rect 11 12 19 14
rect 21 18 26 26
rect 21 16 28 18
rect 21 14 24 16
rect 26 14 28 16
rect 21 12 28 14
rect 32 14 40 26
rect 42 14 47 26
rect 49 24 57 26
rect 49 22 52 24
rect 54 22 57 24
rect 49 14 57 22
rect 32 7 38 14
rect 32 5 34 7
rect 36 5 38 7
rect 32 3 38 5
rect 52 12 57 14
rect 59 16 67 26
rect 59 14 62 16
rect 64 14 67 16
rect 59 12 67 14
rect 69 16 77 26
rect 69 14 72 16
rect 74 14 77 16
rect 69 12 77 14
rect 79 24 86 26
rect 79 22 82 24
rect 84 22 86 24
rect 79 17 86 22
rect 79 15 82 17
rect 84 15 86 17
rect 79 12 86 15
<< pdif >>
rect 4 59 9 65
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 4 38 9 46
rect 11 63 19 65
rect 11 61 14 63
rect 16 61 19 63
rect 11 56 19 61
rect 11 54 14 56
rect 16 54 19 56
rect 11 38 19 54
rect 21 59 26 65
rect 32 63 39 65
rect 32 61 34 63
rect 36 61 39 63
rect 21 57 28 59
rect 21 55 24 57
rect 26 55 28 57
rect 21 50 28 55
rect 21 48 24 50
rect 26 48 28 50
rect 21 46 28 48
rect 32 56 39 61
rect 32 54 34 56
rect 36 54 39 56
rect 21 38 26 46
rect 32 38 39 54
rect 41 38 46 65
rect 48 44 56 65
rect 48 42 51 44
rect 53 42 56 44
rect 48 38 56 42
rect 58 58 66 65
rect 58 56 61 58
rect 63 56 66 58
rect 58 38 66 56
rect 68 63 76 65
rect 68 61 71 63
rect 73 61 76 63
rect 68 56 76 61
rect 68 54 71 56
rect 73 54 76 56
rect 68 38 76 54
rect 78 59 83 65
rect 78 57 85 59
rect 78 55 81 57
rect 83 55 85 57
rect 78 50 85 55
rect 78 48 81 50
rect 83 48 85 50
rect 78 46 85 48
rect 78 38 83 46
<< alu1 >>
rect -2 64 90 72
rect 50 44 54 51
rect 50 43 51 44
rect 2 35 6 43
rect 2 33 14 35
rect 2 31 7 33
rect 9 31 14 33
rect 2 29 14 31
rect 42 42 51 43
rect 53 42 54 44
rect 42 39 54 42
rect 42 25 46 39
rect 58 35 62 51
rect 50 33 62 35
rect 50 31 57 33
rect 59 31 62 33
rect 50 29 62 31
rect 82 35 86 43
rect 74 33 86 35
rect 74 31 82 33
rect 84 31 86 33
rect 74 29 86 31
rect 42 24 56 25
rect 42 22 52 24
rect 54 22 56 24
rect 42 21 56 22
rect -2 7 90 8
rect -2 5 34 7
rect 36 5 90 7
rect -2 0 90 5
<< nmos >>
rect 9 12 11 26
rect 19 12 21 26
rect 40 14 42 26
rect 47 14 49 26
rect 57 12 59 26
rect 67 12 69 26
rect 77 12 79 26
<< pmos >>
rect 9 38 11 65
rect 19 38 21 65
rect 39 38 41 65
rect 46 38 48 65
rect 56 38 58 65
rect 66 38 68 65
rect 76 38 78 65
<< polyct0 >>
rect 19 31 21 33
rect 34 31 36 33
rect 67 31 69 33
<< polyct1 >>
rect 7 31 9 33
rect 57 31 59 33
rect 82 31 84 33
<< ndifct0 >>
rect 4 22 6 24
rect 4 15 6 17
rect 14 14 16 16
rect 24 14 26 16
rect 62 14 64 16
rect 72 14 74 16
rect 82 22 84 24
rect 82 15 84 17
<< ndifct1 >>
rect 52 22 54 24
rect 34 5 36 7
<< pdifct0 >>
rect 4 55 6 57
rect 4 48 6 50
rect 14 61 16 63
rect 14 54 16 56
rect 34 61 36 63
rect 24 55 26 57
rect 24 48 26 50
rect 34 54 36 56
rect 61 56 63 58
rect 71 61 73 63
rect 71 54 73 56
rect 81 55 83 57
rect 81 48 83 50
<< pdifct1 >>
rect 51 42 53 44
<< alu0 >>
rect 12 63 18 64
rect 12 61 14 63
rect 16 61 18 63
rect 3 57 7 59
rect 3 55 4 57
rect 6 55 7 57
rect 3 50 7 55
rect 12 56 18 61
rect 32 63 38 64
rect 32 61 34 63
rect 36 61 38 63
rect 12 54 14 56
rect 16 54 18 56
rect 12 53 18 54
rect 23 57 27 59
rect 23 55 24 57
rect 26 55 27 57
rect 23 50 27 55
rect 32 56 38 61
rect 69 63 75 64
rect 69 61 71 63
rect 73 61 75 63
rect 32 54 34 56
rect 36 54 38 56
rect 32 53 38 54
rect 42 58 65 59
rect 42 56 61 58
rect 63 56 65 58
rect 42 55 65 56
rect 69 56 75 61
rect 42 50 46 55
rect 69 54 71 56
rect 73 54 75 56
rect 69 53 75 54
rect 80 57 84 59
rect 80 55 81 57
rect 83 55 84 57
rect 3 48 4 50
rect 6 48 17 50
rect 3 46 17 48
rect 23 48 24 50
rect 26 48 46 50
rect 23 46 46 48
rect 13 43 17 46
rect 13 39 22 43
rect 18 34 22 39
rect 18 33 38 34
rect 18 31 19 33
rect 21 31 34 33
rect 36 31 38 33
rect 18 30 38 31
rect 18 26 22 30
rect 3 24 22 26
rect 3 22 4 24
rect 6 22 22 24
rect 80 50 84 55
rect 66 48 81 50
rect 83 48 84 50
rect 66 46 84 48
rect 66 33 70 46
rect 66 31 67 33
rect 69 31 70 33
rect 66 26 70 31
rect 66 24 85 26
rect 66 22 82 24
rect 84 22 85 24
rect 3 17 7 22
rect 81 17 85 22
rect 3 15 4 17
rect 6 15 7 17
rect 3 13 7 15
rect 12 16 18 17
rect 12 14 14 16
rect 16 14 18 16
rect 12 8 18 14
rect 22 16 66 17
rect 22 14 24 16
rect 26 14 62 16
rect 64 14 66 16
rect 22 13 66 14
rect 70 16 76 17
rect 70 14 72 16
rect 74 14 76 16
rect 70 8 76 14
rect 81 15 82 17
rect 84 15 85 17
rect 81 13 85 15
<< labels >>
rlabel alu0 5 19 5 19 6 an
rlabel alu0 5 52 5 52 6 an
rlabel alu0 28 32 28 32 6 an
rlabel alu0 25 52 25 52 6 n1
rlabel alu0 44 15 44 15 6 n3
rlabel alu0 68 36 68 36 6 bn
rlabel alu0 53 57 53 57 6 n1
rlabel alu1 12 32 12 32 6 a
rlabel alu1 4 36 4 36 6 a
rlabel alu1 44 4 44 4 6 vss
rlabel alu1 44 32 44 32 6 z
rlabel alu1 52 32 52 32 6 c
rlabel alu1 60 40 60 40 6 c
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 68 44 68 6 vdd
rlabel alu1 76 32 76 32 6 b
rlabel alu1 84 36 84 36 6 b
<< end >>
