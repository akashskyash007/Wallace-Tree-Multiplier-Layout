magic
tech scmos
timestamp 1199203050
<< ab >>
rect 0 0 112 72
<< nwell >>
rect -5 32 117 77
<< pwell >>
rect -5 -5 117 32
<< poly >>
rect 14 65 16 70
rect 21 65 23 70
rect 28 65 30 70
rect 35 65 37 70
rect 47 65 49 70
rect 54 65 56 70
rect 61 65 63 70
rect 68 65 70 70
rect 78 65 80 70
rect 85 65 87 70
rect 92 65 94 70
rect 99 65 101 70
rect 14 37 16 40
rect 9 35 16 37
rect 9 33 11 35
rect 13 33 16 35
rect 9 31 16 33
rect 10 18 12 31
rect 21 27 23 40
rect 17 25 23 27
rect 17 23 19 25
rect 21 23 23 25
rect 17 21 23 23
rect 28 27 30 40
rect 35 35 37 40
rect 47 35 49 38
rect 35 33 49 35
rect 38 31 40 33
rect 42 31 44 33
rect 38 29 44 31
rect 28 25 34 27
rect 28 23 30 25
rect 32 23 34 25
rect 28 21 34 23
rect 20 18 22 21
rect 32 18 34 21
rect 42 18 44 29
rect 54 27 56 38
rect 61 29 63 38
rect 68 35 70 38
rect 78 35 80 38
rect 68 33 81 35
rect 75 31 77 33
rect 79 31 81 33
rect 75 29 81 31
rect 61 27 71 29
rect 48 25 56 27
rect 48 23 50 25
rect 52 23 56 25
rect 65 25 67 27
rect 69 25 71 27
rect 85 25 87 38
rect 65 23 87 25
rect 48 21 56 23
rect 54 19 56 21
rect 92 19 94 38
rect 54 17 94 19
rect 99 19 101 38
rect 99 17 105 19
rect 99 15 101 17
rect 103 15 105 17
rect 99 13 105 15
rect 10 2 12 7
rect 20 2 22 7
rect 32 2 34 7
rect 42 2 44 7
<< ndif >>
rect 2 7 10 18
rect 12 16 20 18
rect 12 14 15 16
rect 17 14 20 16
rect 12 7 20 14
rect 22 7 32 18
rect 34 16 42 18
rect 34 14 37 16
rect 39 14 42 16
rect 34 7 42 14
rect 44 7 52 18
rect 2 5 4 7
rect 6 5 8 7
rect 2 3 8 5
rect 24 5 26 7
rect 28 5 30 7
rect 24 3 30 5
rect 46 5 48 7
rect 50 5 52 7
rect 46 3 52 5
<< pdif >>
rect 39 67 45 69
rect 39 65 41 67
rect 43 65 45 67
rect 9 59 14 65
rect 7 57 14 59
rect 7 55 9 57
rect 11 55 14 57
rect 7 53 14 55
rect 9 40 14 53
rect 16 40 21 65
rect 23 40 28 65
rect 30 40 35 65
rect 37 40 47 65
rect 39 38 47 40
rect 49 38 54 65
rect 56 38 61 65
rect 63 38 68 65
rect 70 57 78 65
rect 70 55 73 57
rect 75 55 78 57
rect 70 38 78 55
rect 80 38 85 65
rect 87 38 92 65
rect 94 38 99 65
rect 101 63 108 65
rect 101 61 104 63
rect 106 61 108 63
rect 101 56 108 61
rect 101 54 104 56
rect 106 54 108 56
rect 101 38 108 54
<< alu1 >>
rect -2 67 114 72
rect -2 65 41 67
rect 43 65 114 67
rect -2 64 114 65
rect 2 57 79 58
rect 2 55 9 57
rect 11 55 73 57
rect 75 55 79 57
rect 2 54 79 55
rect 2 19 6 54
rect 10 46 80 50
rect 10 35 14 46
rect 10 33 11 35
rect 13 33 14 35
rect 10 29 14 33
rect 18 38 70 42
rect 18 25 22 38
rect 38 33 62 34
rect 38 31 40 33
rect 42 31 62 33
rect 38 30 62 31
rect 18 23 19 25
rect 21 23 22 25
rect 18 21 22 23
rect 28 25 54 26
rect 28 23 30 25
rect 32 23 50 25
rect 52 23 54 25
rect 28 22 54 23
rect 2 17 14 19
rect 33 17 41 18
rect 2 16 41 17
rect 2 14 15 16
rect 17 14 37 16
rect 39 14 41 16
rect 2 13 41 14
rect 50 13 54 22
rect 58 18 62 30
rect 66 27 70 38
rect 74 33 80 46
rect 74 31 77 33
rect 79 31 80 33
rect 74 29 80 31
rect 66 25 67 27
rect 69 25 70 27
rect 66 23 70 25
rect 58 17 105 18
rect 58 15 101 17
rect 103 15 105 17
rect 58 14 105 15
rect -2 7 114 8
rect -2 5 4 7
rect 6 5 26 7
rect 28 5 48 7
rect 50 5 65 7
rect 67 5 73 7
rect 75 5 81 7
rect 83 5 89 7
rect 91 5 97 7
rect 99 5 105 7
rect 107 5 114 7
rect -2 0 114 5
<< ptie >>
rect 63 7 109 9
rect 63 5 65 7
rect 67 5 73 7
rect 75 5 81 7
rect 83 5 89 7
rect 91 5 97 7
rect 99 5 105 7
rect 107 5 109 7
rect 63 3 109 5
<< nmos >>
rect 10 7 12 18
rect 20 7 22 18
rect 32 7 34 18
rect 42 7 44 18
<< pmos >>
rect 14 40 16 65
rect 21 40 23 65
rect 28 40 30 65
rect 35 40 37 65
rect 47 38 49 65
rect 54 38 56 65
rect 61 38 63 65
rect 68 38 70 65
rect 78 38 80 65
rect 85 38 87 65
rect 92 38 94 65
rect 99 38 101 65
<< polyct1 >>
rect 11 33 13 35
rect 19 23 21 25
rect 40 31 42 33
rect 30 23 32 25
rect 77 31 79 33
rect 50 23 52 25
rect 67 25 69 27
rect 101 15 103 17
<< ndifct1 >>
rect 15 14 17 16
rect 37 14 39 16
rect 4 5 6 7
rect 26 5 28 7
rect 48 5 50 7
<< ptiect1 >>
rect 65 5 67 7
rect 73 5 75 7
rect 81 5 83 7
rect 89 5 91 7
rect 97 5 99 7
rect 105 5 107 7
<< pdifct0 >>
rect 104 61 106 63
rect 104 54 106 56
<< pdifct1 >>
rect 41 65 43 67
rect 9 55 11 57
rect 73 55 75 57
<< alu0 >>
rect 102 63 108 64
rect 102 61 104 63
rect 106 61 108 63
rect 102 56 108 61
rect 102 54 104 56
rect 106 54 108 56
rect 102 53 108 54
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 36 12 36 6 d
rlabel alu1 12 56 12 56 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 36 24 36 24 6 b
rlabel alu1 20 28 20 28 6 c
rlabel alu1 28 40 28 40 6 c
rlabel alu1 36 40 36 40 6 c
rlabel alu1 20 48 20 48 6 d
rlabel alu1 28 48 28 48 6 d
rlabel alu1 36 48 36 48 6 d
rlabel alu1 28 56 28 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 56 4 56 4 6 vss
rlabel alu1 52 16 52 16 6 b
rlabel alu1 44 24 44 24 6 b
rlabel alu1 60 24 60 24 6 a
rlabel alu1 52 32 52 32 6 a
rlabel alu1 44 32 44 32 6 a
rlabel alu1 44 40 44 40 6 c
rlabel alu1 52 40 52 40 6 c
rlabel alu1 60 40 60 40 6 c
rlabel alu1 44 48 44 48 6 d
rlabel alu1 52 48 52 48 6 d
rlabel alu1 60 48 60 48 6 d
rlabel alu1 52 56 52 56 6 z
rlabel alu1 60 56 60 56 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 56 68 56 68 6 vdd
rlabel alu1 76 16 76 16 6 a
rlabel alu1 84 16 84 16 6 a
rlabel alu1 68 16 68 16 6 a
rlabel alu1 68 32 68 32 6 c
rlabel alu1 76 40 76 40 6 d
rlabel alu1 68 48 68 48 6 d
rlabel alu1 76 56 76 56 6 z
rlabel alu1 68 56 68 56 6 z
rlabel alu1 100 16 100 16 6 a
rlabel alu1 92 16 92 16 6 a
<< end >>
