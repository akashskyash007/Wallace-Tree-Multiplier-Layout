magic
tech scmos
timestamp 1199202824
<< ab >>
rect 0 0 144 80
<< nwell >>
rect -5 36 149 88
<< pwell >>
rect -5 -8 149 36
<< poly >>
rect 20 69 22 74
rect 30 69 32 74
rect 40 69 42 74
rect 50 69 52 74
rect 70 69 72 74
rect 80 69 82 74
rect 100 69 102 74
rect 110 69 112 74
rect 120 69 122 74
rect 20 39 22 42
rect 30 39 32 42
rect 40 39 42 42
rect 10 37 42 39
rect 10 35 12 37
rect 14 35 19 37
rect 21 35 42 37
rect 10 33 42 35
rect 10 30 12 33
rect 20 30 22 33
rect 30 30 32 33
rect 40 30 42 33
rect 50 39 52 42
rect 70 39 72 42
rect 80 39 82 42
rect 100 39 102 42
rect 110 39 112 42
rect 120 39 122 42
rect 50 37 92 39
rect 50 35 52 37
rect 54 35 59 37
rect 61 35 92 37
rect 50 33 92 35
rect 50 30 52 33
rect 60 30 62 33
rect 70 30 72 33
rect 80 30 82 33
rect 90 30 92 33
rect 100 37 132 39
rect 100 35 120 37
rect 122 35 128 37
rect 130 35 132 37
rect 100 33 132 35
rect 100 30 102 33
rect 110 30 112 33
rect 120 30 122 33
rect 130 30 132 33
rect 80 15 82 20
rect 90 15 92 20
rect 10 6 12 10
rect 20 6 22 10
rect 30 6 32 10
rect 40 6 42 10
rect 50 6 52 10
rect 60 6 62 10
rect 70 6 72 10
rect 100 6 102 10
rect 110 6 112 10
rect 120 6 122 10
rect 130 6 132 10
<< ndif >>
rect 3 28 10 30
rect 3 26 5 28
rect 7 26 10 28
rect 3 21 10 26
rect 3 19 5 21
rect 7 19 10 21
rect 3 17 10 19
rect 5 10 10 17
rect 12 21 20 30
rect 12 19 15 21
rect 17 19 20 21
rect 12 14 20 19
rect 12 12 15 14
rect 17 12 20 14
rect 12 10 20 12
rect 22 28 30 30
rect 22 26 25 28
rect 27 26 30 28
rect 22 21 30 26
rect 22 19 25 21
rect 27 19 30 21
rect 22 10 30 19
rect 32 14 40 30
rect 32 12 35 14
rect 37 12 40 14
rect 32 10 40 12
rect 42 21 50 30
rect 42 19 45 21
rect 47 19 50 21
rect 42 10 50 19
rect 52 28 60 30
rect 52 26 55 28
rect 57 26 60 28
rect 52 10 60 26
rect 62 21 70 30
rect 62 19 65 21
rect 67 19 70 21
rect 62 10 70 19
rect 72 28 80 30
rect 72 26 75 28
rect 77 26 80 28
rect 72 20 80 26
rect 82 24 90 30
rect 82 22 85 24
rect 87 22 90 24
rect 82 20 90 22
rect 92 28 100 30
rect 92 26 95 28
rect 97 26 100 28
rect 92 20 100 26
rect 72 10 77 20
rect 95 10 100 20
rect 102 28 110 30
rect 102 26 105 28
rect 107 26 110 28
rect 102 10 110 26
rect 112 20 120 30
rect 112 18 115 20
rect 117 18 120 20
rect 112 10 120 18
rect 122 28 130 30
rect 122 26 125 28
rect 127 26 130 28
rect 122 10 130 26
rect 132 28 139 30
rect 132 26 135 28
rect 137 26 139 28
rect 132 21 139 26
rect 132 19 135 21
rect 137 19 139 21
rect 132 17 139 19
rect 132 10 137 17
<< pdif >>
rect 13 67 20 69
rect 13 65 15 67
rect 17 65 20 67
rect 13 60 20 65
rect 13 58 15 60
rect 17 58 20 60
rect 13 42 20 58
rect 22 53 30 69
rect 22 51 25 53
rect 27 51 30 53
rect 22 46 30 51
rect 22 44 25 46
rect 27 44 30 46
rect 22 42 30 44
rect 32 67 40 69
rect 32 65 35 67
rect 37 65 40 67
rect 32 60 40 65
rect 32 58 35 60
rect 37 58 40 60
rect 32 42 40 58
rect 42 53 50 69
rect 42 51 45 53
rect 47 51 50 53
rect 42 46 50 51
rect 42 44 45 46
rect 47 44 50 46
rect 42 42 50 44
rect 52 67 70 69
rect 52 65 55 67
rect 57 65 65 67
rect 67 65 70 67
rect 52 60 70 65
rect 52 58 55 60
rect 57 58 65 60
rect 67 58 70 60
rect 52 42 70 58
rect 72 53 80 69
rect 72 51 75 53
rect 77 51 80 53
rect 72 46 80 51
rect 72 44 75 46
rect 77 44 80 46
rect 72 42 80 44
rect 82 67 89 69
rect 82 65 85 67
rect 87 65 89 67
rect 82 60 89 65
rect 82 58 85 60
rect 87 58 89 60
rect 82 42 89 58
rect 95 55 100 69
rect 93 53 100 55
rect 93 51 95 53
rect 97 51 100 53
rect 93 46 100 51
rect 93 44 95 46
rect 97 44 100 46
rect 93 42 100 44
rect 102 67 110 69
rect 102 65 105 67
rect 107 65 110 67
rect 102 60 110 65
rect 102 58 105 60
rect 107 58 110 60
rect 102 42 110 58
rect 112 53 120 69
rect 112 51 115 53
rect 117 51 120 53
rect 112 46 120 51
rect 112 44 115 46
rect 117 44 120 46
rect 112 42 120 44
rect 122 67 130 69
rect 122 65 125 67
rect 127 65 130 67
rect 122 60 130 65
rect 122 58 125 60
rect 127 58 130 60
rect 122 42 130 58
<< alu1 >>
rect -2 81 146 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 146 81
rect -2 68 146 79
rect 2 38 6 55
rect 24 53 28 55
rect 24 51 25 53
rect 27 51 28 53
rect 24 46 28 51
rect 44 53 48 55
rect 44 51 45 53
rect 47 51 48 53
rect 44 46 48 51
rect 74 53 78 63
rect 74 51 75 53
rect 77 51 78 53
rect 74 46 78 51
rect 94 53 98 55
rect 94 51 95 53
rect 97 51 98 53
rect 94 46 98 51
rect 114 53 118 55
rect 114 51 115 53
rect 117 51 118 53
rect 114 46 118 51
rect 24 44 25 46
rect 27 44 45 46
rect 47 44 75 46
rect 77 44 95 46
rect 97 44 115 46
rect 117 44 118 46
rect 24 42 118 44
rect 2 37 23 38
rect 2 35 12 37
rect 14 35 19 37
rect 21 35 23 37
rect 2 33 23 35
rect 41 37 63 38
rect 41 35 52 37
rect 54 35 59 37
rect 61 35 63 37
rect 41 34 63 35
rect 41 26 47 34
rect 106 30 110 42
rect 129 38 135 46
rect 118 37 135 38
rect 118 35 120 37
rect 122 35 128 37
rect 130 35 135 37
rect 118 34 135 35
rect 103 28 129 30
rect 103 26 105 28
rect 107 26 125 28
rect 127 26 129 28
rect 103 25 129 26
rect -2 1 146 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 146 1
rect -2 -2 146 -1
<< ptie >>
rect 0 1 144 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 144 1
rect 0 -3 144 -1
<< ntie >>
rect 0 81 144 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 144 81
rect 0 77 144 79
<< nmos >>
rect 10 10 12 30
rect 20 10 22 30
rect 30 10 32 30
rect 40 10 42 30
rect 50 10 52 30
rect 60 10 62 30
rect 70 10 72 30
rect 80 20 82 30
rect 90 20 92 30
rect 100 10 102 30
rect 110 10 112 30
rect 120 10 122 30
rect 130 10 132 30
<< pmos >>
rect 20 42 22 69
rect 30 42 32 69
rect 40 42 42 69
rect 50 42 52 69
rect 70 42 72 69
rect 80 42 82 69
rect 100 42 102 69
rect 110 42 112 69
rect 120 42 122 69
<< polyct1 >>
rect 12 35 14 37
rect 19 35 21 37
rect 52 35 54 37
rect 59 35 61 37
rect 120 35 122 37
rect 128 35 130 37
<< ndifct0 >>
rect 5 26 7 28
rect 5 19 7 21
rect 15 19 17 21
rect 15 12 17 14
rect 25 26 27 28
rect 25 19 27 21
rect 35 12 37 14
rect 45 19 47 21
rect 55 26 57 28
rect 65 19 67 21
rect 75 26 77 28
rect 85 22 87 24
rect 95 26 97 28
rect 115 18 117 20
rect 135 26 137 28
rect 135 19 137 21
<< ndifct1 >>
rect 105 26 107 28
rect 125 26 127 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
<< pdifct0 >>
rect 15 65 17 67
rect 15 58 17 60
rect 35 65 37 67
rect 35 58 37 60
rect 55 65 57 67
rect 65 65 67 67
rect 55 58 57 60
rect 65 58 67 60
rect 85 65 87 67
rect 85 58 87 60
rect 105 65 107 67
rect 105 58 107 60
rect 125 65 127 67
rect 125 58 127 60
<< pdifct1 >>
rect 25 51 27 53
rect 25 44 27 46
rect 45 51 47 53
rect 45 44 47 46
rect 75 51 77 53
rect 75 44 77 46
rect 95 51 97 53
rect 95 44 97 46
rect 115 51 117 53
rect 115 44 117 46
<< alu0 >>
rect 14 67 18 68
rect 14 65 15 67
rect 17 65 18 67
rect 14 60 18 65
rect 14 58 15 60
rect 17 58 18 60
rect 14 56 18 58
rect 34 67 38 68
rect 34 65 35 67
rect 37 65 38 67
rect 34 60 38 65
rect 34 58 35 60
rect 37 58 38 60
rect 34 56 38 58
rect 54 67 58 68
rect 54 65 55 67
rect 57 65 58 67
rect 54 60 58 65
rect 54 58 55 60
rect 57 58 58 60
rect 54 56 58 58
rect 64 67 68 68
rect 64 65 65 67
rect 67 65 68 67
rect 64 60 68 65
rect 84 67 88 68
rect 84 65 85 67
rect 87 65 88 67
rect 64 58 65 60
rect 67 58 68 60
rect 64 56 68 58
rect 84 60 88 65
rect 84 58 85 60
rect 87 58 88 60
rect 84 56 88 58
rect 104 67 108 68
rect 104 65 105 67
rect 107 65 108 67
rect 104 60 108 65
rect 104 58 105 60
rect 107 58 108 60
rect 104 56 108 58
rect 124 67 128 68
rect 124 65 125 67
rect 127 65 128 67
rect 124 60 128 65
rect 124 58 125 60
rect 127 58 128 60
rect 124 56 128 58
rect 4 28 28 30
rect 4 26 5 28
rect 7 26 25 28
rect 27 26 28 28
rect 75 30 98 34
rect 75 29 79 30
rect 53 28 79 29
rect 53 26 55 28
rect 57 26 75 28
rect 77 26 79 28
rect 94 28 98 30
rect 94 26 95 28
rect 97 26 98 28
rect 4 21 8 26
rect 24 22 28 26
rect 53 25 79 26
rect 84 24 88 26
rect 84 22 85 24
rect 87 22 88 24
rect 4 19 5 21
rect 7 19 8 21
rect 4 17 8 19
rect 13 21 19 22
rect 13 19 15 21
rect 17 19 19 21
rect 13 14 19 19
rect 24 21 88 22
rect 24 19 25 21
rect 27 19 45 21
rect 47 19 65 21
rect 67 19 88 21
rect 24 18 88 19
rect 94 21 98 26
rect 134 28 138 30
rect 134 26 135 28
rect 137 26 138 28
rect 134 21 138 26
rect 94 20 135 21
rect 94 18 115 20
rect 117 19 135 20
rect 137 19 138 21
rect 117 18 138 19
rect 94 17 138 18
rect 13 12 15 14
rect 17 12 19 14
rect 33 14 39 15
rect 33 12 35 14
rect 37 12 39 14
<< labels >>
rlabel alu0 6 23 6 23 6 n1
rlabel alu0 26 24 26 24 6 n1
rlabel alu0 66 27 66 27 6 n2
rlabel alu0 56 20 56 20 6 n1
rlabel alu0 96 25 96 25 6 n2
rlabel ndifct0 116 19 116 19 6 n2
rlabel alu0 136 23 136 23 6 n2
rlabel alu1 4 44 4 44 6 a
rlabel alu1 12 36 12 36 6 a
rlabel polyct1 20 36 20 36 6 a
rlabel alu1 44 32 44 32 6 b
rlabel alu1 28 44 28 44 6 z
rlabel alu1 44 44 44 44 6 z
rlabel alu1 52 44 52 44 6 z
rlabel alu1 52 36 52 36 6 b
rlabel alu1 36 44 36 44 6 z
rlabel alu1 72 6 72 6 6 vss
rlabel alu1 60 44 60 44 6 z
rlabel polyct1 60 36 60 36 6 b
rlabel alu1 84 44 84 44 6 z
rlabel alu1 68 44 68 44 6 z
rlabel pdifct1 76 52 76 52 6 z
rlabel alu1 72 74 72 74 6 vdd
rlabel alu1 92 44 92 44 6 z
rlabel alu1 100 44 100 44 6 z
rlabel alu1 108 36 108 36 6 z
rlabel alu1 116 28 116 28 6 z
rlabel alu1 124 28 124 28 6 z
rlabel alu1 132 40 132 40 6 c
rlabel alu1 124 36 124 36 6 c
rlabel pdifct1 116 52 116 52 6 z
<< end >>
