magic
tech scmos
timestamp 1199201865
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 41 70 43 74
rect 9 33 11 43
rect 19 40 21 43
rect 19 38 25 40
rect 19 36 21 38
rect 23 36 25 38
rect 19 34 25 36
rect 29 39 31 43
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 9 27 15 29
rect 12 23 14 27
rect 20 23 22 34
rect 29 33 35 35
rect 30 23 32 33
rect 41 32 43 43
rect 41 30 47 32
rect 41 28 43 30
rect 45 28 47 30
rect 38 26 47 28
rect 38 23 40 26
rect 12 6 14 11
rect 20 6 22 11
rect 30 6 32 11
rect 38 6 40 11
<< ndif >>
rect 3 11 12 23
rect 14 11 20 23
rect 22 20 30 23
rect 22 18 25 20
rect 27 18 30 20
rect 22 11 30 18
rect 32 11 38 23
rect 40 15 48 23
rect 40 13 43 15
rect 45 13 48 15
rect 40 11 48 13
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 57 9 59
rect 4 43 9 57
rect 11 54 19 70
rect 11 52 14 54
rect 16 52 19 54
rect 11 43 19 52
rect 21 61 29 70
rect 21 59 24 61
rect 26 59 29 61
rect 21 43 29 59
rect 31 68 41 70
rect 31 66 35 68
rect 37 66 41 68
rect 31 43 41 66
rect 43 63 48 70
rect 43 61 50 63
rect 43 59 46 61
rect 48 59 50 61
rect 43 57 50 59
rect 43 43 48 57
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 54 18 55
rect 2 52 14 54
rect 16 52 18 54
rect 2 51 18 52
rect 2 23 6 51
rect 26 47 30 55
rect 10 31 14 47
rect 18 41 30 47
rect 34 50 47 54
rect 34 33 38 50
rect 10 29 11 31
rect 13 29 22 31
rect 10 27 22 29
rect 18 25 22 27
rect 26 29 30 31
rect 42 30 46 39
rect 42 29 43 30
rect 26 28 43 29
rect 45 28 46 30
rect 26 25 46 28
rect 2 17 14 23
rect 34 17 38 25
rect -2 11 58 12
rect -2 9 6 11
rect 8 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 12 11 14 23
rect 20 11 22 23
rect 30 11 32 23
rect 38 11 40 23
<< pmos >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 41 43 43 70
<< polyct0 >>
rect 21 36 23 38
rect 31 35 33 37
<< polyct1 >>
rect 11 29 13 31
rect 43 28 45 30
<< ndifct0 >>
rect 25 18 27 20
rect 43 13 45 15
<< ndifct1 >>
rect 6 9 8 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 59 6 61
rect 24 59 26 61
rect 35 66 37 68
rect 46 59 48 61
<< pdifct1 >>
rect 14 52 16 54
<< alu0 >>
rect 33 66 35 68
rect 37 66 39 68
rect 33 65 39 66
rect 2 61 50 62
rect 2 59 4 61
rect 6 59 24 61
rect 26 59 46 61
rect 48 59 50 61
rect 2 58 50 59
rect 20 38 24 41
rect 20 36 21 38
rect 23 36 24 38
rect 20 34 24 36
rect 29 37 34 38
rect 29 35 31 37
rect 33 35 34 37
rect 29 34 34 35
rect 14 20 29 21
rect 14 18 25 20
rect 27 18 29 20
rect 14 17 29 18
rect 42 15 46 17
rect 42 13 43 15
rect 45 13 46 15
rect 42 12 46 13
<< labels >>
rlabel alu0 26 60 26 60 6 n3
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 28 20 28 6 b1
rlabel alu1 20 44 20 44 6 b2
rlabel alu1 12 40 12 40 6 b1
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 20 36 20 6 a1
rlabel alu1 28 28 28 28 6 a1
rlabel alu1 36 40 36 40 6 a2
rlabel alu1 28 48 28 48 6 b2
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 44 52 44 52 6 a2
<< end >>
