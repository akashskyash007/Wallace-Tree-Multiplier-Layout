magic
tech scmos
timestamp 1199203407
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 9 66 11 70
rect 27 66 29 70
rect 37 66 39 70
rect 44 66 46 70
rect 57 66 59 70
rect 67 66 69 70
rect 9 35 11 38
rect 27 35 29 38
rect 9 33 29 35
rect 9 31 11 33
rect 13 31 15 33
rect 37 31 39 38
rect 44 35 46 38
rect 57 35 59 38
rect 9 29 15 31
rect 33 29 39 31
rect 43 33 49 35
rect 43 31 45 33
rect 47 31 49 33
rect 57 33 63 35
rect 57 31 59 33
rect 61 31 63 33
rect 43 29 52 31
rect 57 29 63 31
rect 67 32 69 38
rect 67 30 73 32
rect 11 22 13 29
rect 33 27 35 29
rect 37 27 39 29
rect 21 25 39 27
rect 21 22 23 25
rect 50 23 52 29
rect 60 23 62 29
rect 67 28 69 30
rect 71 28 73 30
rect 67 26 73 28
rect 67 23 69 26
rect 11 4 13 9
rect 21 4 23 9
rect 50 2 52 6
rect 60 2 62 6
rect 67 2 69 6
<< ndif >>
rect 4 13 11 22
rect 4 11 6 13
rect 8 11 11 13
rect 4 9 11 11
rect 13 20 21 22
rect 13 18 16 20
rect 18 18 21 20
rect 13 9 21 18
rect 23 20 31 22
rect 23 18 27 20
rect 29 18 31 20
rect 45 19 50 23
rect 23 16 31 18
rect 42 17 50 19
rect 23 9 28 16
rect 42 15 44 17
rect 46 15 50 17
rect 42 13 50 15
rect 45 6 50 13
rect 52 21 60 23
rect 52 19 55 21
rect 57 19 60 21
rect 52 6 60 19
rect 62 6 67 23
rect 69 10 76 23
rect 69 8 72 10
rect 74 8 76 10
rect 69 6 76 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 44 16 66
rect 22 59 27 66
rect 20 57 27 59
rect 20 55 22 57
rect 24 55 27 57
rect 20 53 27 55
rect 11 42 18 44
rect 11 40 14 42
rect 16 40 18 42
rect 11 38 18 40
rect 22 38 27 53
rect 29 42 37 66
rect 29 40 32 42
rect 34 40 37 42
rect 29 38 37 40
rect 39 38 44 66
rect 46 64 57 66
rect 46 62 50 64
rect 52 62 57 64
rect 46 38 57 62
rect 59 57 67 66
rect 59 55 62 57
rect 64 55 67 57
rect 59 50 67 55
rect 59 48 62 50
rect 64 48 67 50
rect 59 38 67 48
rect 69 64 77 66
rect 69 62 72 64
rect 74 62 77 64
rect 69 57 77 62
rect 69 55 72 57
rect 74 55 77 57
rect 69 38 77 55
<< alu1 >>
rect -2 64 82 72
rect 2 35 6 43
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 2 21 6 29
rect 26 22 30 42
rect 58 37 78 43
rect 58 33 62 37
rect 58 31 59 33
rect 61 31 62 33
rect 58 29 62 31
rect 66 25 78 27
rect 65 21 78 25
rect 34 14 38 18
rect 42 17 46 18
rect 42 15 44 17
rect 42 14 46 15
rect 65 14 71 21
rect -2 7 82 8
rect -2 5 34 7
rect 36 5 82 7
rect -2 0 82 5
<< ptie >>
rect 32 7 38 9
rect 32 5 34 7
rect 36 5 38 7
rect 32 3 38 5
<< nmos >>
rect 11 9 13 22
rect 21 9 23 22
rect 50 6 52 23
rect 60 6 62 23
rect 67 6 69 23
<< pmos >>
rect 9 38 11 66
rect 27 38 29 66
rect 37 38 39 66
rect 44 38 46 66
rect 57 38 59 66
rect 67 38 69 66
<< polyct0 >>
rect 45 31 47 33
rect 35 27 37 29
rect 69 28 71 30
<< polyct1 >>
rect 11 31 13 33
rect 59 31 61 33
<< ndifct0 >>
rect 6 11 8 13
rect 16 18 18 20
rect 27 18 29 20
rect 55 19 57 21
rect 72 8 74 10
<< ndifct1 >>
rect 44 15 46 17
<< ptiect1 >>
rect 34 5 36 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 22 55 24 57
rect 14 40 16 42
rect 32 40 34 42
rect 50 62 52 64
rect 62 55 64 57
rect 62 48 64 50
rect 72 62 74 64
rect 72 55 74 57
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 48 62 50 64
rect 52 62 54 64
rect 48 61 54 62
rect 70 62 72 64
rect 74 62 76 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 20 57 55 58
rect 20 55 22 57
rect 24 55 55 57
rect 20 54 55 55
rect 51 51 55 54
rect 61 57 66 59
rect 61 55 62 57
rect 64 55 66 57
rect 61 51 66 55
rect 70 57 76 62
rect 70 55 72 57
rect 74 55 76 57
rect 70 54 76 55
rect 51 50 66 51
rect 18 46 46 50
rect 18 43 22 46
rect 12 42 22 43
rect 12 40 14 42
rect 16 40 22 42
rect 12 39 22 40
rect 18 21 22 39
rect 14 20 22 21
rect 14 18 16 20
rect 18 18 22 20
rect 14 17 22 18
rect 26 42 36 43
rect 30 40 32 42
rect 34 40 36 42
rect 30 39 36 40
rect 42 35 46 46
rect 51 48 62 50
rect 64 48 66 50
rect 51 47 66 48
rect 42 33 48 35
rect 42 31 45 33
rect 47 31 48 33
rect 34 29 38 31
rect 42 29 48 31
rect 34 27 35 29
rect 37 27 38 29
rect 34 26 38 27
rect 51 26 55 47
rect 68 30 72 32
rect 68 28 69 30
rect 71 28 72 30
rect 68 27 72 28
rect 34 22 55 26
rect 26 20 30 22
rect 26 18 27 20
rect 29 18 30 20
rect 51 21 59 22
rect 51 19 55 21
rect 57 19 59 21
rect 51 18 59 19
rect 5 13 9 15
rect 26 14 34 18
rect 38 14 42 18
rect 46 14 48 18
rect 5 11 6 13
rect 8 11 9 13
rect 5 8 9 11
rect 70 10 76 11
rect 70 8 72 10
rect 74 8 76 10
<< labels >>
rlabel alu0 36 26 36 26 6 an
rlabel alu0 20 33 20 33 6 bn
rlabel alu0 17 41 17 41 6 bn
rlabel alu0 44 39 44 39 6 bn
rlabel alu0 37 56 37 56 6 an
rlabel alu0 53 38 53 38 6 an
rlabel alu0 63 53 63 53 6 an
rlabel alu1 4 32 4 32 6 b
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 36 16 36 16 6 z
rlabel alu1 28 32 28 32 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 44 16 44 16 6 z
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 68 20 68 20 6 a1
rlabel alu1 76 24 76 24 6 a1
rlabel alu1 68 40 68 40 6 a2
rlabel alu1 76 40 76 40 6 a2
rlabel alu1 60 36 60 36 6 a2
<< end >>
