magic
tech scmos
timestamp 1199541661
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 55 94 57 98
rect 67 94 69 98
rect 11 85 13 89
rect 23 86 25 90
rect 33 85 35 89
rect 45 85 47 89
rect 11 53 13 65
rect 23 63 25 66
rect 33 63 35 66
rect 45 63 47 66
rect 19 61 25 63
rect 31 61 35 63
rect 41 61 47 63
rect 19 53 21 61
rect 31 53 33 61
rect 7 51 13 53
rect 7 49 9 51
rect 11 49 13 51
rect 7 47 13 49
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 11 34 13 47
rect 19 34 21 47
rect 27 34 29 47
rect 41 43 43 61
rect 55 53 57 56
rect 67 53 69 56
rect 47 51 69 53
rect 47 49 49 51
rect 51 49 69 51
rect 47 47 69 49
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 35 37 43 39
rect 35 34 37 37
rect 55 25 57 47
rect 67 25 69 47
rect 11 11 13 15
rect 19 11 21 15
rect 27 11 29 15
rect 35 11 37 15
rect 55 2 57 6
rect 67 2 69 6
<< ndif >>
rect 3 15 11 34
rect 13 15 19 34
rect 21 15 27 34
rect 29 15 35 34
rect 37 23 43 34
rect 37 21 45 23
rect 37 19 41 21
rect 43 19 45 21
rect 37 17 45 19
rect 37 15 42 17
rect 3 11 9 15
rect 50 11 55 25
rect 3 9 5 11
rect 7 9 9 11
rect 47 9 55 11
rect 3 7 9 9
rect 47 7 49 9
rect 51 7 55 9
rect 47 6 55 7
rect 57 21 67 25
rect 57 19 61 21
rect 63 19 67 21
rect 57 6 67 19
rect 69 21 77 25
rect 69 19 73 21
rect 75 19 77 21
rect 69 11 77 19
rect 69 9 73 11
rect 75 9 77 11
rect 69 6 77 9
rect 47 5 53 6
<< pdif >>
rect 27 95 33 97
rect 27 93 29 95
rect 31 93 33 95
rect 3 91 9 93
rect 3 89 5 91
rect 7 89 9 91
rect 27 91 33 93
rect 47 95 53 97
rect 47 93 49 95
rect 51 94 53 95
rect 51 93 55 94
rect 47 91 55 93
rect 3 85 9 89
rect 27 86 31 91
rect 15 85 23 86
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 65 11 79
rect 13 81 23 85
rect 13 79 17 81
rect 19 79 23 81
rect 13 66 23 79
rect 25 85 31 86
rect 49 85 55 91
rect 25 66 33 85
rect 35 81 45 85
rect 35 79 39 81
rect 41 79 45 81
rect 35 66 45 79
rect 47 66 55 85
rect 13 65 18 66
rect 49 56 55 66
rect 57 81 67 94
rect 57 79 61 81
rect 63 79 67 81
rect 57 71 67 79
rect 57 69 61 71
rect 63 69 67 71
rect 57 61 67 69
rect 57 59 61 61
rect 63 59 67 61
rect 57 56 67 59
rect 69 91 77 94
rect 69 89 73 91
rect 75 89 77 91
rect 69 81 77 89
rect 69 79 73 81
rect 75 79 77 81
rect 69 71 77 79
rect 69 69 73 71
rect 75 69 77 71
rect 69 61 77 69
rect 69 59 73 61
rect 75 59 77 61
rect 69 56 77 59
<< alu1 >>
rect -2 95 82 100
rect -2 93 29 95
rect 31 93 49 95
rect 51 93 82 95
rect -2 91 82 93
rect -2 89 5 91
rect 7 89 73 91
rect 75 89 82 91
rect -2 88 82 89
rect 4 81 8 88
rect 58 82 62 83
rect 4 79 5 81
rect 7 79 8 81
rect 4 77 8 79
rect 15 81 53 82
rect 15 79 17 81
rect 19 79 39 81
rect 41 79 53 81
rect 15 78 53 79
rect 8 51 12 73
rect 8 49 9 51
rect 11 49 12 51
rect 8 17 12 49
rect 18 51 22 73
rect 18 49 19 51
rect 21 49 22 51
rect 18 17 22 49
rect 28 51 32 73
rect 28 49 29 51
rect 31 49 32 51
rect 28 17 32 49
rect 38 41 42 73
rect 49 52 53 78
rect 47 51 53 52
rect 47 49 49 51
rect 51 49 53 51
rect 47 48 53 49
rect 38 39 39 41
rect 41 39 42 41
rect 38 27 42 39
rect 49 22 53 48
rect 39 21 53 22
rect 39 19 41 21
rect 43 19 53 21
rect 39 18 53 19
rect 58 81 65 82
rect 58 79 61 81
rect 63 79 65 81
rect 58 78 65 79
rect 72 81 76 88
rect 72 79 73 81
rect 75 79 76 81
rect 58 72 62 78
rect 58 71 65 72
rect 58 69 61 71
rect 63 69 65 71
rect 58 68 65 69
rect 72 71 76 79
rect 72 69 73 71
rect 75 69 76 71
rect 58 62 62 68
rect 58 61 65 62
rect 58 59 61 61
rect 63 59 65 61
rect 58 58 65 59
rect 72 61 76 69
rect 72 59 73 61
rect 75 59 76 61
rect 58 22 62 58
rect 72 57 76 59
rect 58 21 65 22
rect 58 19 61 21
rect 63 19 65 21
rect 58 18 65 19
rect 72 21 76 23
rect 72 19 73 21
rect 75 19 76 21
rect 58 17 62 18
rect 72 12 76 19
rect -2 11 82 12
rect -2 9 5 11
rect 7 9 73 11
rect 75 9 82 11
rect -2 7 49 9
rect 51 7 82 9
rect -2 5 19 7
rect 21 5 35 7
rect 37 5 82 7
rect -2 0 82 5
<< ptie >>
rect 17 7 39 9
rect 17 5 19 7
rect 21 5 35 7
rect 37 5 39 7
rect 17 3 39 5
<< nmos >>
rect 11 15 13 34
rect 19 15 21 34
rect 27 15 29 34
rect 35 15 37 34
rect 55 6 57 25
rect 67 6 69 25
<< pmos >>
rect 11 65 13 85
rect 23 66 25 86
rect 33 66 35 85
rect 45 66 47 85
rect 55 56 57 94
rect 67 56 69 94
<< polyct1 >>
rect 9 49 11 51
rect 19 49 21 51
rect 29 49 31 51
rect 49 49 51 51
rect 39 39 41 41
<< ndifct1 >>
rect 41 19 43 21
rect 5 9 7 11
rect 49 7 51 9
rect 61 19 63 21
rect 73 19 75 21
rect 73 9 75 11
<< ptiect1 >>
rect 19 5 21 7
rect 35 5 37 7
<< pdifct1 >>
rect 29 93 31 95
rect 5 89 7 91
rect 49 93 51 95
rect 5 79 7 81
rect 17 79 19 81
rect 39 79 41 81
rect 61 79 63 81
rect 61 69 63 71
rect 61 59 63 61
rect 73 89 75 91
rect 73 79 75 81
rect 73 69 75 71
rect 73 59 75 61
<< labels >>
rlabel alu1 10 45 10 45 6 i0
rlabel alu1 20 45 20 45 6 i1
rlabel alu1 30 45 30 45 6 i2
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 40 50 40 50 6 i3
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 60 50 60 50 6 q
<< end >>
