magic
tech scmos
timestamp 1199469309
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -2 48 82 104
<< pwell >>
rect -2 -4 82 48
<< poly >>
rect 11 83 13 88
rect 23 83 25 88
rect 31 83 33 88
rect 43 83 45 88
rect 55 83 57 88
rect 67 83 69 88
rect 11 53 13 63
rect 23 53 25 63
rect 11 51 27 53
rect 11 49 17 51
rect 19 49 27 51
rect 11 47 27 49
rect 13 26 15 47
rect 25 33 27 47
rect 31 42 33 63
rect 43 54 45 63
rect 43 52 49 54
rect 43 50 45 52
rect 47 50 49 52
rect 43 48 49 50
rect 31 40 41 42
rect 31 38 37 40
rect 39 38 41 40
rect 31 36 41 38
rect 33 33 35 36
rect 45 33 47 48
rect 55 42 57 63
rect 67 52 69 57
rect 63 50 69 52
rect 63 48 65 50
rect 67 48 69 50
rect 63 46 69 48
rect 53 40 59 42
rect 53 38 55 40
rect 57 38 59 40
rect 53 36 59 38
rect 67 37 69 46
rect 57 33 59 36
rect 25 19 27 24
rect 33 19 35 24
rect 45 19 47 24
rect 57 19 59 24
rect 13 12 15 17
rect 67 19 69 24
<< ndif >>
rect 61 33 67 37
rect 17 26 25 33
rect 8 23 13 26
rect 5 21 13 23
rect 5 19 7 21
rect 9 19 13 21
rect 5 17 13 19
rect 15 24 25 26
rect 27 24 33 33
rect 35 31 45 33
rect 35 29 39 31
rect 41 29 45 31
rect 35 24 45 29
rect 47 28 57 33
rect 47 26 51 28
rect 53 26 57 28
rect 47 24 57 26
rect 59 24 67 33
rect 69 35 77 37
rect 69 33 73 35
rect 75 33 77 35
rect 69 31 77 33
rect 69 24 74 31
rect 15 17 23 24
rect 17 11 23 17
rect 61 17 65 24
rect 61 15 67 17
rect 61 13 63 15
rect 65 13 67 15
rect 61 11 67 13
rect 17 9 19 11
rect 21 9 23 11
rect 17 7 23 9
<< pdif >>
rect 3 81 11 83
rect 3 79 5 81
rect 7 79 11 81
rect 3 73 11 79
rect 3 71 5 73
rect 7 71 11 73
rect 3 69 11 71
rect 6 63 11 69
rect 13 81 23 83
rect 13 79 17 81
rect 19 79 23 81
rect 13 63 23 79
rect 25 63 31 83
rect 33 71 43 83
rect 33 69 37 71
rect 39 69 43 71
rect 33 63 43 69
rect 45 81 55 83
rect 45 79 49 81
rect 51 79 55 81
rect 45 63 55 79
rect 57 81 67 83
rect 57 79 61 81
rect 63 79 67 81
rect 57 63 67 79
rect 59 57 67 63
rect 69 63 74 83
rect 69 61 77 63
rect 69 59 73 61
rect 75 59 77 61
rect 69 57 77 59
<< alu1 >>
rect -2 95 82 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 82 95
rect -2 88 82 93
rect 4 81 8 83
rect 4 79 5 81
rect 7 79 8 81
rect 4 73 8 79
rect 16 81 20 88
rect 16 79 17 81
rect 19 79 20 81
rect 16 77 20 79
rect 26 81 53 82
rect 26 79 49 81
rect 51 79 53 81
rect 26 78 53 79
rect 60 81 64 88
rect 60 79 61 81
rect 63 79 64 81
rect 4 71 5 73
rect 7 72 8 73
rect 26 72 30 78
rect 60 77 64 79
rect 7 71 30 72
rect 4 68 30 71
rect 36 71 42 73
rect 36 69 37 71
rect 39 69 42 71
rect 36 63 42 69
rect 8 53 12 63
rect 28 57 42 63
rect 8 51 22 53
rect 8 49 17 51
rect 19 49 22 51
rect 8 47 22 49
rect 8 37 12 47
rect 28 32 32 57
rect 48 53 52 73
rect 38 52 52 53
rect 38 50 45 52
rect 47 50 52 52
rect 38 47 52 50
rect 58 67 72 73
rect 58 52 62 67
rect 72 61 76 63
rect 72 59 73 61
rect 75 59 76 61
rect 58 50 68 52
rect 58 48 65 50
rect 67 48 68 50
rect 58 46 68 48
rect 72 42 76 59
rect 36 40 76 42
rect 36 38 37 40
rect 39 38 55 40
rect 57 38 76 40
rect 36 36 76 38
rect 72 35 76 36
rect 72 33 73 35
rect 75 33 76 35
rect 28 31 43 32
rect 72 31 76 33
rect 28 29 39 31
rect 41 29 43 31
rect 28 27 43 29
rect 49 28 55 29
rect 49 26 51 28
rect 53 26 55 28
rect 49 22 55 26
rect 5 21 55 22
rect 5 19 7 21
rect 9 19 55 21
rect 5 18 55 19
rect 62 15 66 17
rect 62 13 63 15
rect 65 13 66 15
rect 62 12 66 13
rect -2 11 82 12
rect -2 9 19 11
rect 21 9 82 11
rect -2 7 82 9
rect -2 5 39 7
rect 41 5 49 7
rect 51 5 82 7
rect -2 0 82 5
<< ptie >>
rect 37 7 53 9
rect 37 5 39 7
rect 41 5 49 7
rect 51 5 53 7
rect 37 3 53 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 13 17 15 26
rect 25 24 27 33
rect 33 24 35 33
rect 45 24 47 33
rect 57 24 59 33
rect 67 24 69 37
<< pmos >>
rect 11 63 13 83
rect 23 63 25 83
rect 31 63 33 83
rect 43 63 45 83
rect 55 63 57 83
rect 67 57 69 83
<< polyct1 >>
rect 17 49 19 51
rect 45 50 47 52
rect 37 38 39 40
rect 65 48 67 50
rect 55 38 57 40
<< ndifct1 >>
rect 7 19 9 21
rect 39 29 41 31
rect 51 26 53 28
rect 73 33 75 35
rect 63 13 65 15
rect 19 9 21 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 39 5 41 7
rect 49 5 51 7
<< pdifct1 >>
rect 5 79 7 81
rect 5 71 7 73
rect 17 79 19 81
rect 37 69 39 71
rect 49 79 51 81
rect 61 79 63 81
rect 73 59 75 61
<< labels >>
rlabel alu1 10 50 10 50 6 b
rlabel alu1 6 75 6 75 6 n2
rlabel alu1 20 50 20 50 6 b
rlabel alu1 17 70 17 70 6 n2
rlabel ptiect1 40 6 40 6 6 vss
rlabel ndifct1 40 30 40 30 6 z
rlabel alu1 30 45 30 45 6 z
rlabel alu1 40 50 40 50 6 c
rlabel alu1 40 65 40 65 6 z
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 52 23 52 23 6 n4
rlabel alu1 30 20 30 20 6 n4
rlabel alu1 60 60 60 60 6 a
rlabel alu1 50 60 50 60 6 c
rlabel alu1 39 80 39 80 6 n2
rlabel polyct1 56 39 56 39 6 an
rlabel alu1 74 47 74 47 6 an
rlabel alu1 70 70 70 70 6 a
<< end >>
