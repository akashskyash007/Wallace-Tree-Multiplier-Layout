magic
tech scmos
timestamp 1199202116
<< ab >>
rect 0 0 152 80
<< nwell >>
rect -5 36 157 88
<< pwell >>
rect -5 -8 157 36
<< poly >>
rect 19 69 21 74
rect 29 69 31 74
rect 39 69 41 74
rect 49 69 51 74
rect 59 69 61 74
rect 71 69 73 74
rect 78 69 80 74
rect 88 69 90 74
rect 95 69 97 74
rect 107 69 109 74
rect 117 69 119 74
rect 127 69 129 74
rect 9 59 11 64
rect 137 59 139 64
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 71 39 73 42
rect 78 39 80 42
rect 88 39 90 42
rect 95 39 97 42
rect 9 37 21 39
rect 9 35 11 37
rect 13 35 21 37
rect 9 33 21 35
rect 25 37 32 39
rect 25 35 27 37
rect 29 35 32 37
rect 25 33 32 35
rect 39 37 52 39
rect 39 35 48 37
rect 50 35 52 37
rect 39 33 52 35
rect 59 37 73 39
rect 59 35 67 37
rect 69 35 73 37
rect 59 33 73 35
rect 77 37 90 39
rect 77 35 86 37
rect 88 35 90 37
rect 77 33 90 35
rect 94 37 102 39
rect 94 35 98 37
rect 100 35 102 37
rect 94 33 102 35
rect 107 33 109 42
rect 117 33 119 42
rect 127 38 129 42
rect 137 38 139 42
rect 9 30 11 33
rect 19 30 21 33
rect 30 30 32 33
rect 40 30 42 33
rect 50 30 52 33
rect 60 30 62 33
rect 70 30 72 33
rect 77 30 79 33
rect 87 30 89 33
rect 94 30 96 33
rect 106 31 119 33
rect 9 15 11 19
rect 19 15 21 19
rect 30 11 32 16
rect 40 11 42 16
rect 50 11 52 16
rect 60 11 62 16
rect 70 15 72 19
rect 77 14 79 19
rect 106 29 115 31
rect 117 29 119 31
rect 106 27 119 29
rect 126 36 139 38
rect 126 34 135 36
rect 137 34 139 36
rect 126 32 139 34
rect 106 24 108 27
rect 116 24 118 27
rect 126 24 128 32
rect 136 24 138 32
rect 87 12 89 17
rect 94 12 96 17
rect 106 6 108 10
rect 116 6 118 10
rect 126 8 128 13
rect 136 8 138 13
<< ndif >>
rect 2 19 9 30
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 19 19 26
rect 21 20 30 30
rect 21 19 25 20
rect 2 13 7 19
rect 23 18 25 19
rect 27 18 30 20
rect 23 16 30 18
rect 32 21 40 30
rect 32 19 35 21
rect 37 19 40 21
rect 32 16 40 19
rect 42 28 50 30
rect 42 26 45 28
rect 47 26 50 28
rect 42 16 50 26
rect 52 21 60 30
rect 52 19 55 21
rect 57 19 60 21
rect 52 16 60 19
rect 62 19 70 30
rect 72 19 77 30
rect 79 28 87 30
rect 79 26 82 28
rect 84 26 87 28
rect 79 19 87 26
rect 62 16 68 19
rect 2 11 8 13
rect 64 13 68 16
rect 82 17 87 19
rect 89 17 94 30
rect 96 24 104 30
rect 96 17 106 24
rect 64 11 70 13
rect 98 14 106 17
rect 98 12 100 14
rect 102 12 106 14
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
rect 64 9 66 11
rect 68 9 70 11
rect 98 10 106 12
rect 108 21 116 24
rect 108 19 111 21
rect 113 19 116 21
rect 108 10 116 19
rect 118 17 126 24
rect 118 15 121 17
rect 123 15 126 17
rect 118 13 126 15
rect 128 22 136 24
rect 128 20 131 22
rect 133 20 136 22
rect 128 13 136 20
rect 138 17 146 24
rect 138 15 141 17
rect 143 15 146 17
rect 138 13 146 15
rect 118 10 124 13
rect 64 7 70 9
<< pdif >>
rect 99 71 105 73
rect 99 69 101 71
rect 103 69 105 71
rect 14 59 19 69
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 49 9 55
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 11 53 19 59
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 60 39 69
rect 31 58 34 60
rect 36 58 39 60
rect 31 42 39 58
rect 41 46 49 69
rect 41 44 44 46
rect 46 44 49 46
rect 41 42 49 44
rect 51 60 59 69
rect 51 58 54 60
rect 56 58 59 60
rect 51 42 59 58
rect 61 67 71 69
rect 61 65 65 67
rect 67 65 71 67
rect 61 42 71 65
rect 73 42 78 69
rect 80 46 88 69
rect 80 44 83 46
rect 85 44 88 46
rect 80 42 88 44
rect 90 42 95 69
rect 97 42 107 69
rect 109 60 117 69
rect 109 58 112 60
rect 114 58 117 60
rect 109 53 117 58
rect 109 51 112 53
rect 114 51 117 53
rect 109 42 117 51
rect 119 67 127 69
rect 119 65 122 67
rect 124 65 127 67
rect 119 59 127 65
rect 119 57 122 59
rect 124 57 127 59
rect 119 42 127 57
rect 129 59 134 69
rect 129 54 137 59
rect 129 52 132 54
rect 134 52 137 54
rect 129 47 137 52
rect 129 45 132 47
rect 134 45 137 47
rect 129 42 137 45
rect 139 57 146 59
rect 139 55 142 57
rect 144 55 146 57
rect 139 49 146 55
rect 139 47 142 49
rect 144 47 146 49
rect 139 42 146 47
<< alu1 >>
rect -2 81 154 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 154 81
rect -2 71 154 79
rect -2 69 101 71
rect 103 69 154 71
rect -2 68 154 69
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 2 17 6 33
rect 34 46 48 47
rect 34 44 44 46
rect 46 44 48 46
rect 34 42 48 44
rect 34 30 38 42
rect 57 38 63 46
rect 46 37 63 38
rect 46 35 48 37
rect 50 35 63 37
rect 46 34 63 35
rect 74 46 87 47
rect 74 44 83 46
rect 85 44 87 46
rect 74 42 87 44
rect 74 30 78 42
rect 34 28 87 30
rect 34 26 45 28
rect 47 26 82 28
rect 84 26 87 28
rect 74 25 87 26
rect 130 36 142 39
rect 130 34 135 36
rect 137 34 142 36
rect 130 33 142 34
rect 138 25 142 33
rect -2 11 154 12
rect -2 9 4 11
rect 6 9 66 11
rect 68 9 154 11
rect -2 1 154 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 154 1
rect -2 -2 154 -1
<< ptie >>
rect 0 1 152 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 152 1
rect 0 -3 152 -1
<< ntie >>
rect 0 81 152 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 152 81
rect 0 77 152 79
<< nmos >>
rect 9 19 11 30
rect 19 19 21 30
rect 30 16 32 30
rect 40 16 42 30
rect 50 16 52 30
rect 60 16 62 30
rect 70 19 72 30
rect 77 19 79 30
rect 87 17 89 30
rect 94 17 96 30
rect 106 10 108 24
rect 116 10 118 24
rect 126 13 128 24
rect 136 13 138 24
<< pmos >>
rect 9 42 11 59
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 49 42 51 69
rect 59 42 61 69
rect 71 42 73 69
rect 78 42 80 69
rect 88 42 90 69
rect 95 42 97 69
rect 107 42 109 69
rect 117 42 119 69
rect 127 42 129 69
rect 137 42 139 59
<< polyct0 >>
rect 27 35 29 37
rect 67 35 69 37
rect 86 35 88 37
rect 98 35 100 37
rect 115 29 117 31
<< polyct1 >>
rect 11 35 13 37
rect 48 35 50 37
rect 135 34 137 36
<< ndifct0 >>
rect 14 26 16 28
rect 25 18 27 20
rect 35 19 37 21
rect 55 19 57 21
rect 100 12 102 14
rect 111 19 113 21
rect 121 15 123 17
rect 131 20 133 22
rect 141 15 143 17
<< ndifct1 >>
rect 45 26 47 28
rect 82 26 84 28
rect 4 9 6 11
rect 66 9 68 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
<< pdifct0 >>
rect 4 55 6 57
rect 4 47 6 49
rect 14 51 16 53
rect 14 44 16 46
rect 24 65 26 67
rect 24 58 26 60
rect 34 58 36 60
rect 54 58 56 60
rect 65 65 67 67
rect 112 58 114 60
rect 112 51 114 53
rect 122 65 124 67
rect 122 57 124 59
rect 132 52 134 54
rect 132 45 134 47
rect 142 55 144 57
rect 142 47 144 49
<< pdifct1 >>
rect 101 69 103 71
rect 44 44 46 46
rect 83 44 85 46
<< alu0 >>
rect 3 57 7 68
rect 22 67 28 68
rect 22 65 24 67
rect 26 65 28 67
rect 22 60 28 65
rect 63 67 69 68
rect 63 65 65 67
rect 67 65 69 67
rect 63 64 69 65
rect 121 67 125 68
rect 121 65 122 67
rect 124 65 125 67
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 32 60 116 61
rect 32 58 34 60
rect 36 58 54 60
rect 56 58 112 60
rect 114 58 116 60
rect 32 57 116 58
rect 3 55 4 57
rect 6 55 7 57
rect 3 49 7 55
rect 3 47 4 49
rect 6 47 7 49
rect 3 45 7 47
rect 12 53 101 54
rect 12 51 14 53
rect 16 51 101 53
rect 12 50 101 51
rect 110 53 116 57
rect 121 59 125 65
rect 121 57 122 59
rect 124 57 125 59
rect 121 55 125 57
rect 141 57 145 68
rect 110 51 112 53
rect 114 51 116 53
rect 110 50 116 51
rect 131 54 135 56
rect 131 52 132 54
rect 134 52 135 54
rect 12 46 18 50
rect 12 44 14 46
rect 16 44 18 46
rect 12 43 18 44
rect 26 37 30 50
rect 26 35 27 37
rect 29 35 30 37
rect 26 29 30 35
rect 12 28 30 29
rect 12 26 14 28
rect 16 26 30 28
rect 66 37 70 50
rect 66 35 67 37
rect 69 35 70 37
rect 66 33 70 35
rect 84 37 94 38
rect 84 35 86 37
rect 88 35 94 37
rect 84 34 94 35
rect 12 25 30 26
rect 43 25 49 26
rect 90 29 94 34
rect 97 37 101 50
rect 131 47 135 52
rect 97 35 98 37
rect 100 35 101 37
rect 97 33 101 35
rect 114 45 132 47
rect 134 45 135 47
rect 141 55 142 57
rect 144 55 145 57
rect 141 49 145 55
rect 141 47 142 49
rect 144 47 145 49
rect 141 45 145 47
rect 114 43 135 45
rect 114 31 118 43
rect 114 29 115 31
rect 117 29 118 31
rect 90 25 134 29
rect 130 22 134 25
rect 33 21 115 22
rect 23 20 29 21
rect 23 18 25 20
rect 27 18 29 20
rect 33 19 35 21
rect 37 19 55 21
rect 57 19 111 21
rect 113 19 115 21
rect 130 20 131 22
rect 133 20 134 22
rect 33 18 115 19
rect 23 12 29 18
rect 120 17 124 19
rect 130 18 134 20
rect 120 15 121 17
rect 123 15 124 17
rect 98 14 104 15
rect 98 12 100 14
rect 102 12 104 14
rect 120 12 124 15
rect 140 17 144 19
rect 140 15 141 17
rect 143 15 144 17
rect 140 12 144 15
<< labels >>
rlabel alu0 21 27 21 27 6 an
rlabel alu0 15 48 15 48 6 an
rlabel alu0 28 39 28 39 6 an
rlabel alu0 68 43 68 43 6 an
rlabel alu0 74 20 74 20 6 n3
rlabel alu0 116 36 116 36 6 bn
rlabel alu0 89 36 89 36 6 bn
rlabel alu0 113 55 113 55 6 n1
rlabel alu0 99 43 99 43 6 an
rlabel alu0 74 59 74 59 6 n1
rlabel alu0 132 23 132 23 6 bn
rlabel alu0 133 49 133 49 6 bn
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 4 28 4 28 6 a
rlabel alu1 68 28 68 28 6 z
rlabel alu1 60 28 60 28 6 z
rlabel alu1 52 36 52 36 6 c
rlabel alu1 52 28 52 28 6 z
rlabel alu1 44 28 44 28 6 z
rlabel alu1 44 44 44 44 6 z
rlabel alu1 60 40 60 40 6 c
rlabel alu1 36 40 36 40 6 z
rlabel alu1 76 6 76 6 6 vss
rlabel alu1 76 36 76 36 6 z
rlabel alu1 84 28 84 28 6 z
rlabel alu1 84 44 84 44 6 z
rlabel alu1 76 74 76 74 6 vdd
rlabel alu1 132 36 132 36 6 b
rlabel alu1 140 32 140 32 6 b
<< end >>
