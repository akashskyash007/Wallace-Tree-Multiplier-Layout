magic
tech scmos
timestamp 1199202595
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 10 61 12 66
rect 20 61 22 65
rect 10 39 12 47
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 23 11 33
rect 20 32 22 47
rect 20 30 26 32
rect 20 28 22 30
rect 24 28 26 30
rect 16 26 26 28
rect 16 23 18 26
rect 9 6 11 11
rect 16 6 18 11
<< ndif >>
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 11 9 17
rect 11 11 16 23
rect 18 15 30 23
rect 18 13 26 15
rect 28 13 30 15
rect 18 11 30 13
<< pdif >>
rect 2 61 8 63
rect 2 59 4 61
rect 6 59 10 61
rect 2 47 10 59
rect 12 59 20 61
rect 12 57 15 59
rect 17 57 20 59
rect 12 52 20 57
rect 12 50 15 52
rect 17 50 20 52
rect 12 47 20 50
rect 22 59 30 61
rect 22 57 26 59
rect 28 57 30 59
rect 22 52 30 57
rect 22 50 26 52
rect 28 50 30 52
rect 22 47 30 50
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 50 15 54
rect 2 23 6 50
rect 17 42 23 46
rect 10 38 23 42
rect 10 37 14 38
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 18 30 30 31
rect 18 28 22 30
rect 24 28 30 30
rect 18 25 30 28
rect 2 21 7 23
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect 18 17 22 25
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 11 11 23
rect 16 11 18 23
<< pmos >>
rect 10 47 12 61
rect 20 47 22 61
<< polyct1 >>
rect 11 35 13 37
rect 22 28 24 30
<< ndifct0 >>
rect 26 13 28 15
<< ndifct1 >>
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 59 6 61
rect 15 57 17 59
rect 15 50 17 52
rect 26 57 28 59
rect 26 50 28 52
<< alu0 >>
rect 2 61 8 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 59 19 60
rect 13 57 15 59
rect 17 57 19 59
rect 13 54 19 57
rect 15 52 19 54
rect 17 50 19 52
rect 6 49 19 50
rect 24 59 30 68
rect 24 57 26 59
rect 28 57 30 59
rect 24 52 30 57
rect 24 50 26 52
rect 28 50 30 52
rect 24 49 30 50
rect 25 15 29 17
rect 25 13 26 15
rect 28 13 29 15
rect 25 12 29 13
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 24 20 24 6 a
rlabel alu1 20 44 20 44 6 b
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 28 28 28 6 a
<< end >>
