magic
tech scmos
timestamp 1199202174
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 26 67 44 69
rect 9 58 11 63
rect 19 58 21 63
rect 26 58 28 67
rect 42 63 44 67
rect 36 58 38 63
rect 42 61 48 63
rect 46 58 48 61
rect 9 37 11 42
rect 19 37 21 42
rect 9 35 21 37
rect 9 32 11 35
rect 5 30 11 32
rect 19 30 21 35
rect 26 30 28 42
rect 36 39 38 42
rect 32 37 38 39
rect 32 35 34 37
rect 36 35 38 37
rect 32 33 38 35
rect 36 30 38 33
rect 46 39 48 42
rect 46 37 53 39
rect 46 35 49 37
rect 51 35 53 37
rect 46 33 53 35
rect 46 30 48 33
rect 5 28 7 30
rect 9 28 11 30
rect 5 26 11 28
rect 9 23 11 26
rect 19 18 21 23
rect 26 18 28 23
rect 36 18 38 23
rect 46 19 48 23
rect 9 11 11 16
<< ndif >>
rect 13 23 19 30
rect 21 23 26 30
rect 28 28 36 30
rect 28 26 31 28
rect 33 26 36 28
rect 28 23 36 26
rect 38 27 46 30
rect 38 25 41 27
rect 43 25 46 27
rect 38 23 46 25
rect 48 23 54 30
rect 2 20 9 23
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 17 23
rect 50 17 54 23
rect 13 11 19 16
rect 48 15 54 17
rect 48 13 50 15
rect 52 13 54 15
rect 48 11 54 13
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 48 69 54 71
rect 13 65 19 69
rect 13 58 17 65
rect 48 67 50 69
rect 52 67 54 69
rect 48 65 54 67
rect 50 58 54 65
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 4 42 9 45
rect 11 42 19 58
rect 21 42 26 58
rect 28 54 36 58
rect 28 52 31 54
rect 33 52 36 54
rect 28 42 36 52
rect 38 56 46 58
rect 38 54 41 56
rect 43 54 46 56
rect 38 42 46 54
rect 48 42 54 58
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 15 71
rect 17 69 58 71
rect -2 68 50 69
rect 52 68 58 69
rect 10 54 35 55
rect 10 52 31 54
rect 33 52 35 54
rect 10 51 35 52
rect 10 49 22 51
rect 2 31 6 39
rect 2 30 14 31
rect 2 28 7 30
rect 9 28 14 30
rect 2 25 14 28
rect 18 30 22 49
rect 26 38 30 47
rect 50 46 54 55
rect 41 42 54 46
rect 26 37 39 38
rect 26 35 34 37
rect 36 35 39 37
rect 26 34 39 35
rect 48 37 54 42
rect 48 35 49 37
rect 51 35 54 37
rect 48 33 54 35
rect 18 28 35 30
rect 18 26 31 28
rect 33 26 35 28
rect 18 25 35 26
rect -2 11 58 12
rect -2 9 15 11
rect 17 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 19 23 21 30
rect 26 23 28 30
rect 36 23 38 30
rect 46 23 48 30
rect 9 16 11 23
<< pmos >>
rect 9 42 11 58
rect 19 42 21 58
rect 26 42 28 58
rect 36 42 38 58
rect 46 42 48 58
<< polyct1 >>
rect 34 35 36 37
rect 49 35 51 37
rect 7 28 9 30
<< ndifct0 >>
rect 41 25 43 27
rect 4 18 6 20
rect 50 13 52 15
<< ndifct1 >>
rect 31 26 33 28
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 50 67 52 68
rect 4 54 6 56
rect 4 47 6 49
rect 41 54 43 56
<< pdifct1 >>
rect 15 69 17 71
rect 50 68 52 69
rect 31 52 33 54
<< alu0 >>
rect 49 67 50 68
rect 52 67 53 68
rect 49 65 53 67
rect 3 59 44 63
rect 3 56 7 59
rect 3 54 4 56
rect 6 54 7 56
rect 40 56 44 59
rect 3 49 7 54
rect 40 54 41 56
rect 43 54 44 56
rect 40 52 44 54
rect 3 47 4 49
rect 6 47 7 49
rect 3 45 7 47
rect 40 27 44 29
rect 40 25 41 27
rect 43 25 44 27
rect 40 21 44 25
rect 2 20 44 21
rect 2 18 4 20
rect 6 18 44 20
rect 2 17 44 18
rect 49 15 53 17
rect 49 13 50 15
rect 52 13 53 15
rect 49 12 53 13
<< labels >>
rlabel alu0 5 54 5 54 6 n1
rlabel alu0 42 23 42 23 6 n3
rlabel alu0 23 19 23 19 6 n3
rlabel alu0 42 57 42 57 6 n1
rlabel alu1 4 32 4 32 6 a
rlabel alu1 12 28 12 28 6 a
rlabel alu1 20 40 20 40 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 28 28 28 6 z
rlabel alu1 36 36 36 36 6 c
rlabel alu1 28 44 28 44 6 c
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 52 44 52 44 6 b
rlabel alu1 44 44 44 44 6 b
<< end >>
