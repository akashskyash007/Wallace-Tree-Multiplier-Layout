magic
tech scmos
timestamp 1199202998
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 18 70 20 74
rect 25 70 27 74
rect 32 70 34 74
rect 45 66 47 71
rect 45 47 47 50
rect 41 45 47 47
rect 41 43 43 45
rect 45 43 47 45
rect 18 39 20 42
rect 9 37 20 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 25 11 33
rect 25 32 27 42
rect 32 33 34 42
rect 41 41 47 43
rect 22 30 28 32
rect 22 28 24 30
rect 26 28 28 30
rect 22 26 28 28
rect 32 31 40 33
rect 32 29 36 31
rect 38 29 40 31
rect 32 27 40 29
rect 22 22 24 26
rect 32 22 34 27
rect 45 24 47 41
rect 9 15 11 19
rect 22 11 24 16
rect 32 11 34 16
rect 45 11 47 16
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 22 19 25
rect 36 22 45 24
rect 11 19 22 22
rect 13 16 22 19
rect 24 20 32 22
rect 24 18 27 20
rect 29 18 32 20
rect 24 16 32 18
rect 34 20 45 22
rect 34 18 39 20
rect 41 18 45 20
rect 34 16 45 18
rect 47 22 54 24
rect 47 20 50 22
rect 52 20 54 22
rect 47 18 54 20
rect 47 16 52 18
rect 13 11 19 16
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 13 63 18 70
rect 11 61 18 63
rect 11 59 13 61
rect 15 59 18 61
rect 11 54 18 59
rect 11 52 13 54
rect 15 52 18 54
rect 11 50 18 52
rect 13 42 18 50
rect 20 42 25 70
rect 27 42 32 70
rect 34 68 43 70
rect 34 66 39 68
rect 41 66 43 68
rect 34 61 45 66
rect 34 59 39 61
rect 41 59 45 61
rect 34 50 45 59
rect 47 63 52 66
rect 47 61 54 63
rect 47 59 50 61
rect 52 59 54 61
rect 47 54 54 59
rect 47 52 50 54
rect 52 52 54 54
rect 47 50 54 52
rect 34 42 39 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 11 61 17 62
rect 11 59 13 61
rect 15 59 17 61
rect 11 55 17 59
rect 2 54 17 55
rect 2 52 13 54
rect 15 52 17 54
rect 2 51 17 52
rect 2 25 6 51
rect 34 47 38 55
rect 10 41 22 47
rect 34 45 46 47
rect 34 43 43 45
rect 45 43 46 45
rect 34 41 46 43
rect 10 37 14 41
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 26 31 30 39
rect 18 30 30 31
rect 18 28 24 30
rect 26 28 30 30
rect 18 25 30 28
rect 2 23 7 25
rect 2 21 4 23
rect 6 21 14 23
rect 2 20 31 21
rect 2 18 27 20
rect 29 18 31 20
rect 2 17 31 18
rect -2 11 58 12
rect -2 9 15 11
rect 17 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 19 11 25
rect 22 16 24 22
rect 32 16 34 22
rect 45 16 47 24
<< pmos >>
rect 18 42 20 70
rect 25 42 27 70
rect 32 42 34 70
rect 45 50 47 66
<< polyct0 >>
rect 36 29 38 31
<< polyct1 >>
rect 43 43 45 45
rect 11 35 13 37
rect 24 28 26 30
<< ndifct0 >>
rect 39 18 41 20
rect 50 20 52 22
<< ndifct1 >>
rect 4 21 6 23
rect 27 18 29 20
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 39 66 41 68
rect 39 59 41 61
rect 50 59 52 61
rect 50 52 52 54
<< pdifct1 >>
rect 13 59 15 61
rect 13 52 15 54
<< alu0 >>
rect 37 66 39 68
rect 41 66 43 68
rect 37 61 43 66
rect 37 59 39 61
rect 41 59 43 61
rect 37 58 43 59
rect 49 61 54 63
rect 49 59 50 61
rect 52 59 54 61
rect 49 54 54 59
rect 49 52 50 54
rect 52 52 54 54
rect 49 50 54 52
rect 50 32 54 50
rect 34 31 54 32
rect 34 29 36 31
rect 38 29 54 31
rect 34 28 54 29
rect 49 22 53 28
rect 37 20 43 21
rect 37 18 39 20
rect 41 18 43 20
rect 49 20 50 22
rect 52 20 53 22
rect 49 18 53 20
rect 37 12 43 18
<< labels >>
rlabel alu0 51 25 51 25 6 an
rlabel alu0 44 30 44 30 6 an
rlabel alu0 52 45 52 45 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 44 20 44 6 c
rlabel alu1 12 40 12 40 6 c
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 32 28 32 6 b
rlabel alu1 36 48 36 48 6 a
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 44 44 44 6 a
<< end >>
