magic
tech scmos
timestamp 1199203206
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 22 70 24 74
rect 29 70 31 74
rect 9 61 11 65
rect 9 40 11 49
rect 22 47 24 52
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 19 41 25 43
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 9 25 11 34
rect 19 25 21 41
rect 29 39 31 52
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 29 25 31 33
rect 9 15 11 19
rect 19 15 21 19
rect 29 15 31 19
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 23 19 25
rect 11 21 14 23
rect 16 21 19 23
rect 11 19 19 21
rect 21 23 29 25
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 31 23 38 25
rect 31 21 34 23
rect 36 21 38 23
rect 31 19 38 21
<< pdif >>
rect 13 68 22 70
rect 13 66 16 68
rect 18 66 22 68
rect 13 61 22 66
rect 2 59 9 61
rect 2 57 4 59
rect 6 57 9 59
rect 2 55 9 57
rect 4 49 9 55
rect 11 52 22 61
rect 24 52 29 70
rect 31 63 36 70
rect 31 61 38 63
rect 31 59 34 61
rect 36 59 38 61
rect 31 57 38 59
rect 31 52 36 57
rect 11 49 19 52
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 59 15 62
rect 2 57 4 59
rect 6 58 15 59
rect 2 25 6 57
rect 26 46 30 55
rect 17 45 30 46
rect 17 43 21 45
rect 23 43 30 45
rect 17 42 30 43
rect 34 38 38 47
rect 25 37 38 38
rect 25 35 31 37
rect 33 35 38 37
rect 25 34 38 35
rect 34 33 38 34
rect 2 23 7 25
rect 2 21 4 23
rect 6 21 7 23
rect 2 17 7 21
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 19 31 25
<< pmos >>
rect 9 49 11 61
rect 22 52 24 70
rect 29 52 31 70
<< polyct0 >>
rect 11 36 13 38
<< polyct1 >>
rect 21 43 23 45
rect 31 35 33 37
<< ndifct0 >>
rect 14 21 16 23
rect 24 21 26 23
rect 34 21 36 23
<< ndifct1 >>
rect 4 21 6 23
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 16 66 18 68
rect 34 59 36 61
<< pdifct1 >>
rect 4 57 6 59
<< alu0 >>
rect 14 66 16 68
rect 18 66 20 68
rect 14 65 20 66
rect 18 61 38 62
rect 18 59 34 61
rect 36 59 38 61
rect 18 58 38 59
rect 6 55 7 58
rect 18 54 22 58
rect 10 50 22 54
rect 10 38 14 50
rect 10 36 11 38
rect 13 36 14 38
rect 10 31 14 36
rect 10 27 27 31
rect 12 23 18 24
rect 12 21 14 23
rect 16 21 18 23
rect 12 12 18 21
rect 23 23 27 27
rect 23 21 24 23
rect 26 21 27 23
rect 23 19 27 21
rect 32 23 38 24
rect 32 21 34 23
rect 36 21 38 23
rect 32 12 38 21
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 25 25 25 25 6 zn
rlabel alu0 28 60 28 60 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 44 20 44 6 a
rlabel alu1 28 52 28 52 6 a
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 40 36 40 6 b
<< end >>
