magic
tech scmos
timestamp 1199201714
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 62 11 67
rect 19 62 21 67
rect 29 62 31 67
rect 41 61 43 66
rect 9 39 11 44
rect 19 39 21 49
rect 29 46 31 49
rect 29 44 35 46
rect 29 42 31 44
rect 33 42 35 44
rect 29 40 35 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 29 11 33
rect 22 29 24 33
rect 29 29 31 40
rect 41 39 43 48
rect 41 37 47 39
rect 41 35 43 37
rect 45 35 47 37
rect 36 33 47 35
rect 36 29 38 33
rect 9 15 11 20
rect 22 11 24 16
rect 29 11 31 16
rect 36 11 38 16
<< ndif >>
rect 2 27 9 29
rect 2 25 4 27
rect 6 25 9 27
rect 2 23 9 25
rect 4 20 9 23
rect 11 20 22 29
rect 13 16 22 20
rect 24 16 29 29
rect 31 16 36 29
rect 38 22 43 29
rect 38 20 45 22
rect 38 18 41 20
rect 43 18 45 20
rect 38 16 45 18
rect 13 11 20 16
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 33 71 39 73
rect 33 69 35 71
rect 37 69 39 71
rect 33 62 39 69
rect 4 57 9 62
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 48 9 53
rect 2 46 4 48
rect 6 46 9 48
rect 2 44 9 46
rect 11 60 19 62
rect 11 58 14 60
rect 16 58 19 60
rect 11 49 19 58
rect 21 60 29 62
rect 21 58 24 60
rect 26 58 29 60
rect 21 53 29 58
rect 21 51 24 53
rect 26 51 29 53
rect 21 49 29 51
rect 31 61 39 62
rect 31 49 41 61
rect 11 44 17 49
rect 36 48 41 49
rect 43 59 50 61
rect 43 57 46 59
rect 48 57 50 59
rect 43 52 50 57
rect 43 50 46 52
rect 48 50 50 52
rect 43 48 50 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 35 71
rect 37 69 58 71
rect -2 68 58 69
rect 2 55 7 63
rect 2 53 4 55
rect 6 54 7 55
rect 6 53 15 54
rect 2 50 15 53
rect 2 48 6 50
rect 2 46 4 48
rect 2 27 6 46
rect 33 46 39 54
rect 25 44 47 46
rect 25 42 31 44
rect 33 42 47 44
rect 17 37 30 38
rect 17 35 21 37
rect 23 35 30 37
rect 17 34 30 35
rect 2 25 4 27
rect 2 17 6 25
rect 26 25 30 34
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 31 47 35
rect 34 25 47 31
rect -2 11 58 12
rect -2 9 15 11
rect 17 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 20 11 29
rect 22 16 24 29
rect 29 16 31 29
rect 36 16 38 29
<< pmos >>
rect 9 44 11 62
rect 19 49 21 62
rect 29 49 31 62
rect 41 48 43 61
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 42 33 44
rect 21 35 23 37
rect 43 35 45 37
<< ndifct0 >>
rect 41 18 43 20
<< ndifct1 >>
rect 4 25 6 27
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 14 58 16 60
rect 24 58 26 60
rect 24 51 26 53
rect 46 57 48 59
rect 46 50 48 52
<< pdifct1 >>
rect 35 69 37 71
rect 4 53 6 55
rect 4 46 6 48
<< alu0 >>
rect 12 60 18 68
rect 12 58 14 60
rect 16 58 18 60
rect 12 57 18 58
rect 23 60 50 62
rect 23 58 24 60
rect 26 59 50 60
rect 26 58 46 59
rect 23 53 27 58
rect 44 57 46 58
rect 48 57 50 59
rect 18 51 24 53
rect 26 51 27 53
rect 6 44 7 50
rect 18 49 27 51
rect 18 46 22 49
rect 44 52 50 57
rect 44 50 46 52
rect 48 50 50 52
rect 44 49 50 50
rect 10 42 22 46
rect 10 37 14 42
rect 29 41 35 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 6 23 7 29
rect 10 25 19 29
rect 15 21 19 25
rect 15 20 45 21
rect 15 18 41 20
rect 43 18 45 20
rect 15 17 45 18
<< labels >>
rlabel alu0 12 35 12 35 6 zn
rlabel alu0 25 55 25 55 6 zn
rlabel alu0 30 19 30 19 6 zn
rlabel alu0 47 55 47 55 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 36 20 36 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 28 28 28 6 a
rlabel alu1 36 28 36 28 6 c
rlabel alu1 28 44 28 44 6 b
rlabel alu1 36 48 36 48 6 b
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 c
rlabel polyct1 44 36 44 36 6 c
rlabel alu1 44 44 44 44 6 b
<< end >>
