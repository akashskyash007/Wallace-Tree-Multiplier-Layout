magic
tech scmos
timestamp 1199202693
<< ab >>
rect 0 0 112 72
<< nwell >>
rect -5 32 117 77
<< pwell >>
rect -5 -5 117 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 90 56 92 61
rect 100 56 102 61
rect 9 35 11 39
rect 19 35 21 39
rect 29 35 31 39
rect 39 35 41 39
rect 49 35 51 39
rect 59 35 61 39
rect 69 35 71 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 33 35
rect 19 31 27 33
rect 29 31 33 33
rect 19 29 33 31
rect 12 26 14 29
rect 19 26 21 29
rect 31 26 33 29
rect 38 33 51 35
rect 38 31 43 33
rect 45 31 51 33
rect 38 29 51 31
rect 55 33 71 35
rect 79 35 81 39
rect 90 35 92 39
rect 100 35 102 39
rect 79 33 92 35
rect 96 33 102 35
rect 55 31 59 33
rect 61 31 63 33
rect 55 29 63 31
rect 81 31 83 33
rect 85 31 87 33
rect 81 29 87 31
rect 96 31 98 33
rect 100 31 102 33
rect 96 29 102 31
rect 38 26 40 29
rect 48 26 50 29
rect 55 26 57 29
rect 12 7 14 12
rect 19 7 21 12
rect 31 2 33 7
rect 38 2 40 7
rect 48 2 50 7
rect 55 2 57 7
<< ndif >>
rect 5 24 12 26
rect 5 22 7 24
rect 9 22 12 24
rect 5 17 12 22
rect 5 15 7 17
rect 9 15 12 17
rect 5 12 12 15
rect 14 12 19 26
rect 21 12 31 26
rect 23 7 31 12
rect 33 7 38 26
rect 40 17 48 26
rect 40 15 43 17
rect 45 15 48 17
rect 40 7 48 15
rect 50 7 55 26
rect 57 7 66 26
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
rect 59 5 61 7
rect 63 5 66 7
rect 59 3 66 5
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 39 9 55
rect 11 56 19 66
rect 11 54 14 56
rect 16 54 19 56
rect 11 49 19 54
rect 11 47 14 49
rect 16 47 19 49
rect 11 39 19 47
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 39 29 55
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 49 39 55
rect 31 47 34 49
rect 36 47 39 49
rect 31 39 39 47
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 39 49 55
rect 51 56 59 66
rect 51 54 54 56
rect 56 54 59 56
rect 51 49 59 54
rect 51 47 54 49
rect 56 47 59 49
rect 51 39 59 47
rect 61 64 69 66
rect 61 62 64 64
rect 66 62 69 64
rect 61 57 69 62
rect 61 55 64 57
rect 66 55 69 57
rect 61 39 69 55
rect 71 57 79 66
rect 71 55 74 57
rect 76 55 79 57
rect 71 49 79 55
rect 71 47 74 49
rect 76 47 79 49
rect 71 39 79 47
rect 81 64 88 66
rect 81 62 84 64
rect 86 62 88 64
rect 81 57 88 62
rect 81 55 84 57
rect 86 56 88 57
rect 86 55 90 56
rect 81 39 90 55
rect 92 49 100 56
rect 92 47 95 49
rect 97 47 100 49
rect 92 39 100 47
rect 102 54 110 56
rect 102 52 105 54
rect 107 52 110 54
rect 102 46 110 52
rect 102 44 105 46
rect 107 44 110 46
rect 102 39 110 44
<< alu1 >>
rect -2 67 114 72
rect -2 65 97 67
rect 99 65 105 67
rect 107 65 114 67
rect -2 64 114 65
rect 33 57 38 59
rect 33 55 34 57
rect 36 55 38 57
rect 33 50 38 55
rect 73 57 78 59
rect 73 55 74 57
rect 76 55 78 57
rect 73 50 78 55
rect 2 49 99 50
rect 2 47 14 49
rect 16 47 34 49
rect 36 47 54 49
rect 56 47 74 49
rect 76 47 95 49
rect 97 47 99 49
rect 2 46 99 47
rect 2 25 6 46
rect 25 38 97 42
rect 10 33 20 35
rect 10 31 11 33
rect 13 31 20 33
rect 10 29 20 31
rect 25 33 31 38
rect 25 31 27 33
rect 29 31 31 33
rect 25 30 31 31
rect 41 33 47 34
rect 41 31 43 33
rect 45 31 47 33
rect 16 26 20 29
rect 41 26 47 31
rect 57 33 63 38
rect 93 34 97 38
rect 57 31 59 33
rect 61 31 63 33
rect 57 30 63 31
rect 81 33 87 34
rect 81 31 83 33
rect 85 31 87 33
rect 81 26 87 31
rect 93 33 103 34
rect 93 31 98 33
rect 100 31 103 33
rect 93 30 103 31
rect 2 24 11 25
rect 2 22 7 24
rect 9 22 11 24
rect 16 22 87 26
rect 2 21 11 22
rect 7 18 11 21
rect 7 17 47 18
rect 9 15 43 17
rect 45 15 47 17
rect 7 14 47 15
rect -2 7 114 8
rect -2 5 25 7
rect 27 5 61 7
rect 63 5 83 7
rect 85 5 91 7
rect 93 5 114 7
rect -2 0 114 5
<< ptie >>
rect 81 7 95 24
rect 81 5 83 7
rect 85 5 91 7
rect 93 5 95 7
rect 81 3 95 5
<< ntie >>
rect 95 67 109 69
rect 95 65 97 67
rect 99 65 105 67
rect 107 65 109 67
rect 95 63 109 65
<< nmos >>
rect 12 12 14 26
rect 19 12 21 26
rect 31 7 33 26
rect 38 7 40 26
rect 48 7 50 26
rect 55 7 57 26
<< pmos >>
rect 9 39 11 66
rect 19 39 21 66
rect 29 39 31 66
rect 39 39 41 66
rect 49 39 51 66
rect 59 39 61 66
rect 69 39 71 66
rect 79 39 81 66
rect 90 39 92 56
rect 100 39 102 56
<< polyct1 >>
rect 11 31 13 33
rect 27 31 29 33
rect 43 31 45 33
rect 59 31 61 33
rect 83 31 85 33
rect 98 31 100 33
<< ndifct1 >>
rect 7 22 9 24
rect 7 15 9 17
rect 43 15 45 17
rect 25 5 27 7
rect 61 5 63 7
<< ntiect1 >>
rect 97 65 99 67
rect 105 65 107 67
<< ptiect1 >>
rect 83 5 85 7
rect 91 5 93 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 54 16 56
rect 24 62 26 64
rect 24 55 26 57
rect 44 62 46 64
rect 44 55 46 57
rect 54 54 56 56
rect 64 62 66 64
rect 64 55 66 57
rect 84 62 86 64
rect 84 55 86 57
rect 105 52 107 54
rect 105 44 107 46
<< pdifct1 >>
rect 14 47 16 49
rect 34 55 36 57
rect 34 47 36 49
rect 54 47 56 49
rect 74 55 76 57
rect 74 47 76 49
rect 95 47 97 49
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 56 17 58
rect 13 54 14 56
rect 16 54 17 56
rect 22 57 28 62
rect 42 62 44 64
rect 46 62 48 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 13 50 17 54
rect 42 57 48 62
rect 62 62 64 64
rect 66 62 68 64
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 53 56 57 58
rect 53 54 54 56
rect 56 54 57 56
rect 62 57 68 62
rect 82 62 84 64
rect 86 62 88 64
rect 62 55 64 57
rect 66 55 68 57
rect 62 54 68 55
rect 53 50 57 54
rect 82 57 88 62
rect 82 55 84 57
rect 86 55 88 57
rect 82 54 88 55
rect 104 54 108 64
rect 104 52 105 54
rect 107 52 108 54
rect 104 46 108 52
rect 104 44 105 46
rect 107 44 108 46
rect 104 42 108 44
rect 5 14 7 21
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 24 20 24 6 b
rlabel alu1 28 24 28 24 6 b
rlabel alu1 36 24 36 24 6 b
rlabel polyct1 28 32 28 32 6 a
rlabel alu1 36 40 36 40 6 a
rlabel alu1 28 36 28 36 6 a
rlabel alu1 20 48 20 48 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 56 4 56 4 6 vss
rlabel ndifct1 44 16 44 16 6 z
rlabel alu1 52 24 52 24 6 b
rlabel alu1 60 24 60 24 6 b
rlabel alu1 44 28 44 28 6 b
rlabel alu1 44 40 44 40 6 a
rlabel alu1 52 40 52 40 6 a
rlabel alu1 60 36 60 36 6 a
rlabel alu1 44 48 44 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 56 68 56 68 6 vdd
rlabel alu1 68 24 68 24 6 b
rlabel alu1 76 24 76 24 6 b
rlabel alu1 84 28 84 28 6 b
rlabel alu1 68 40 68 40 6 a
rlabel alu1 76 40 76 40 6 a
rlabel alu1 84 40 84 40 6 a
rlabel alu1 68 48 68 48 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 84 48 84 48 6 z
rlabel alu1 100 32 100 32 6 a
rlabel alu1 92 40 92 40 6 a
rlabel alu1 92 48 92 48 6 z
<< end >>
