magic
tech scmos
timestamp 1199542936
<< ab >>
rect 0 0 130 100
<< nwell >>
rect -2 48 132 104
<< pwell >>
rect -2 -4 132 48
<< poly >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 69 95 71 98
rect 81 95 83 98
rect 93 95 95 98
rect 105 95 107 98
rect 117 75 119 78
rect 11 53 13 55
rect 23 53 25 55
rect 35 53 37 55
rect 47 53 49 55
rect 69 53 71 55
rect 81 53 83 55
rect 11 51 19 53
rect 23 51 29 53
rect 35 51 43 53
rect 17 43 19 51
rect 27 43 29 51
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 67 51 73 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 77 51 83 53
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 17 29 19 37
rect 27 29 29 37
rect 37 29 39 47
rect 47 29 49 47
rect 15 27 19 29
rect 23 27 29 29
rect 35 27 39 29
rect 43 27 49 29
rect 69 29 71 47
rect 69 27 75 29
rect 15 25 17 27
rect 23 25 25 27
rect 35 25 37 27
rect 43 25 45 27
rect 73 25 75 27
rect 81 25 83 47
rect 93 41 95 55
rect 105 43 107 55
rect 105 41 113 43
rect 93 39 109 41
rect 111 39 113 41
rect 93 25 95 39
rect 105 37 113 39
rect 105 25 107 37
rect 117 33 119 55
rect 111 31 119 33
rect 111 29 113 31
rect 115 29 119 31
rect 111 27 119 29
rect 117 25 119 27
rect 117 12 119 15
rect 15 2 17 5
rect 23 2 25 5
rect 35 2 37 5
rect 43 2 45 5
rect 73 2 75 5
rect 81 2 83 5
rect 93 2 95 5
rect 105 2 107 5
<< ndif >>
rect 97 31 103 33
rect 97 29 99 31
rect 101 29 103 31
rect 97 25 103 29
rect 7 11 15 25
rect 7 9 9 11
rect 11 9 15 11
rect 7 5 15 9
rect 17 5 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 5 35 19
rect 37 5 43 25
rect 45 11 53 25
rect 45 9 49 11
rect 51 9 53 11
rect 45 5 53 9
rect 65 21 73 25
rect 65 19 67 21
rect 69 19 73 21
rect 65 5 73 19
rect 75 5 81 25
rect 83 11 93 25
rect 83 9 87 11
rect 89 9 93 11
rect 83 5 93 9
rect 95 5 105 25
rect 107 15 117 25
rect 119 21 127 25
rect 119 19 123 21
rect 125 19 127 21
rect 119 15 127 19
rect 107 11 115 15
rect 107 9 111 11
rect 113 9 115 11
rect 107 5 115 9
<< pdif >>
rect 3 81 11 95
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 71 23 95
rect 13 69 17 71
rect 19 69 23 71
rect 13 55 23 69
rect 25 81 35 95
rect 25 79 29 81
rect 31 79 35 81
rect 25 55 35 79
rect 37 71 47 95
rect 37 69 41 71
rect 43 69 47 71
rect 37 55 47 69
rect 49 83 53 95
rect 61 93 69 95
rect 61 91 63 93
rect 65 91 69 93
rect 61 89 69 91
rect 49 81 57 83
rect 49 79 53 81
rect 55 79 57 81
rect 49 55 57 79
rect 63 55 69 89
rect 71 81 81 95
rect 71 79 75 81
rect 77 79 81 81
rect 71 55 81 79
rect 83 91 93 95
rect 83 89 87 91
rect 89 89 93 91
rect 83 81 93 89
rect 83 79 87 81
rect 89 79 93 81
rect 83 71 93 79
rect 83 69 87 71
rect 89 69 93 71
rect 83 55 93 69
rect 95 81 105 95
rect 95 79 99 81
rect 101 79 105 81
rect 95 71 105 79
rect 95 69 99 71
rect 101 69 105 71
rect 95 61 105 69
rect 95 59 99 61
rect 101 59 105 61
rect 95 55 105 59
rect 107 91 115 95
rect 107 89 111 91
rect 113 89 115 91
rect 107 81 115 89
rect 107 79 111 81
rect 113 79 115 81
rect 107 75 115 79
rect 107 71 117 75
rect 107 69 111 71
rect 113 69 117 71
rect 107 55 117 69
rect 119 71 127 75
rect 119 69 123 71
rect 125 69 127 71
rect 119 61 127 69
rect 119 59 123 61
rect 125 59 127 61
rect 119 55 127 59
<< alu1 >>
rect -2 93 132 100
rect -2 91 63 93
rect 65 91 123 93
rect 125 91 132 93
rect -2 89 87 91
rect 89 89 111 91
rect 113 89 132 91
rect -2 88 132 89
rect 4 81 8 82
rect 28 81 32 82
rect 52 81 56 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 53 81
rect 55 79 56 81
rect 4 78 8 79
rect 28 78 32 79
rect 52 78 56 79
rect 74 81 78 82
rect 74 79 75 81
rect 77 79 78 81
rect 74 78 78 79
rect 86 81 90 88
rect 86 79 87 81
rect 89 79 90 81
rect 16 71 20 72
rect 16 70 17 71
rect 9 69 17 70
rect 19 69 20 71
rect 9 68 20 69
rect 9 21 11 68
rect 18 41 22 62
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 28 41 32 72
rect 40 71 44 72
rect 75 71 77 78
rect 40 69 41 71
rect 43 69 77 71
rect 86 71 90 79
rect 86 69 87 71
rect 89 69 90 71
rect 40 68 44 69
rect 86 68 90 69
rect 98 81 102 82
rect 98 79 99 81
rect 101 79 102 81
rect 98 71 102 79
rect 98 69 99 71
rect 101 69 102 71
rect 28 39 29 41
rect 31 39 32 41
rect 28 28 32 39
rect 38 51 42 62
rect 38 49 39 51
rect 41 49 42 51
rect 38 28 42 49
rect 48 51 52 62
rect 48 49 49 51
rect 51 49 52 51
rect 48 28 52 49
rect 68 51 72 62
rect 68 49 69 51
rect 71 49 72 51
rect 68 28 72 49
rect 78 51 82 62
rect 78 49 79 51
rect 81 49 82 51
rect 78 28 82 49
rect 98 61 102 69
rect 110 81 114 88
rect 110 79 111 81
rect 113 79 114 81
rect 110 71 114 79
rect 110 69 111 71
rect 113 69 114 71
rect 110 68 114 69
rect 122 71 126 72
rect 122 69 123 71
rect 125 69 126 71
rect 122 68 126 69
rect 123 62 125 68
rect 98 59 99 61
rect 101 59 102 61
rect 98 31 102 59
rect 122 61 126 62
rect 122 59 123 61
rect 125 59 126 61
rect 122 58 126 59
rect 108 41 112 42
rect 123 41 125 58
rect 108 39 109 41
rect 111 39 125 41
rect 108 38 112 39
rect 98 29 99 31
rect 101 29 102 31
rect 98 28 102 29
rect 112 31 116 32
rect 112 29 113 31
rect 115 29 116 31
rect 112 28 116 29
rect 28 21 32 22
rect 66 21 70 22
rect 113 21 115 28
rect 123 22 125 39
rect 9 19 29 21
rect 31 19 67 21
rect 69 19 115 21
rect 122 21 126 22
rect 122 19 123 21
rect 125 19 126 21
rect 28 18 32 19
rect 66 18 70 19
rect 122 18 126 19
rect -2 11 132 12
rect -2 9 9 11
rect 11 9 49 11
rect 51 9 87 11
rect 89 9 111 11
rect 113 9 132 11
rect -2 0 132 9
<< ntie >>
rect 121 93 127 95
rect 121 91 123 93
rect 125 91 127 93
rect 121 83 127 91
<< nmos >>
rect 15 5 17 25
rect 23 5 25 25
rect 35 5 37 25
rect 43 5 45 25
rect 73 5 75 25
rect 81 5 83 25
rect 93 5 95 25
rect 105 5 107 25
rect 117 15 119 25
<< pmos >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 69 55 71 95
rect 81 55 83 95
rect 93 55 95 95
rect 105 55 107 95
rect 117 55 119 75
<< polyct1 >>
rect 39 49 41 51
rect 49 49 51 51
rect 69 49 71 51
rect 79 49 81 51
rect 19 39 21 41
rect 29 39 31 41
rect 109 39 111 41
rect 113 29 115 31
<< ndifct1 >>
rect 99 29 101 31
rect 9 9 11 11
rect 29 19 31 21
rect 49 9 51 11
rect 67 19 69 21
rect 87 9 89 11
rect 123 19 125 21
rect 111 9 113 11
<< ntiect1 >>
rect 123 91 125 93
<< pdifct1 >>
rect 5 79 7 81
rect 17 69 19 71
rect 29 79 31 81
rect 41 69 43 71
rect 63 91 65 93
rect 53 79 55 81
rect 75 79 77 81
rect 87 89 89 91
rect 87 79 89 81
rect 87 69 89 71
rect 99 79 101 81
rect 99 69 101 71
rect 99 59 101 61
rect 111 89 113 91
rect 111 79 113 81
rect 111 69 113 71
rect 123 69 125 71
rect 123 59 125 61
<< labels >>
rlabel alu1 20 45 20 45 6 i5
rlabel alu1 40 45 40 45 6 i3
rlabel alu1 30 50 30 50 6 i4
rlabel alu1 65 6 65 6 6 vss
rlabel alu1 70 45 70 45 6 i1
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 65 94 65 94 6 vdd
rlabel alu1 80 45 80 45 6 i0
rlabel alu1 100 55 100 55 6 nq
<< end >>
