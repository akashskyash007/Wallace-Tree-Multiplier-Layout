magic
tech scmos
timestamp 1199202288
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 70 11 74
rect 9 39 11 42
rect 9 37 16 39
rect 9 35 12 37
rect 14 35 16 37
rect 9 33 16 35
rect 9 30 11 33
rect 9 6 11 11
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 11 9 17
rect 11 23 19 30
rect 11 21 14 23
rect 16 21 19 23
rect 11 15 19 21
rect 11 13 14 15
rect 16 13 19 15
rect 11 11 19 13
<< pdif >>
rect 4 56 9 70
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 42 9 45
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 42 19 59
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 68 26 79
rect 2 54 14 55
rect 2 52 4 54
rect 6 52 14 54
rect 2 49 14 52
rect 2 47 6 49
rect 2 45 4 47
rect 2 29 6 45
rect 18 39 22 55
rect 10 37 22 39
rect 10 35 12 37
rect 14 35 22 37
rect 10 33 22 35
rect 2 28 8 29
rect 2 26 4 28
rect 6 26 8 28
rect 2 21 8 26
rect 2 19 4 21
rect 6 19 8 21
rect 2 17 8 19
rect -2 1 26 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 11 11 30
<< pmos >>
rect 9 42 11 70
<< polyct1 >>
rect 12 35 14 37
<< ndifct0 >>
rect 14 21 16 23
rect 14 13 16 15
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct0 >>
rect 14 66 16 68
rect 14 59 16 61
<< pdifct1 >>
rect 4 52 6 54
rect 4 45 6 47
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 61 18 66
rect 12 59 14 61
rect 16 59 18 61
rect 12 58 18 59
rect 6 43 7 49
rect 13 23 17 25
rect 13 21 14 23
rect 16 21 17 23
rect 13 15 17 21
rect 13 13 14 15
rect 16 13 17 15
rect 13 12 17 13
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 36 12 36 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 44 20 44 6 a
<< end >>
