magic
tech scmos
timestamp 1199202671
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 14 58 16 63
rect 24 58 26 63
rect 35 58 37 63
rect 45 58 47 63
rect 14 39 16 42
rect 24 39 26 42
rect 35 39 37 42
rect 45 39 47 42
rect 9 37 26 39
rect 9 35 11 37
rect 13 35 26 37
rect 9 33 26 35
rect 24 30 26 33
rect 31 37 47 39
rect 31 35 43 37
rect 45 35 47 37
rect 31 33 47 35
rect 31 30 33 33
rect 24 12 26 17
rect 31 12 33 17
<< ndif >>
rect 17 28 24 30
rect 17 26 19 28
rect 21 26 24 28
rect 17 21 24 26
rect 17 19 19 21
rect 21 19 24 21
rect 17 17 24 19
rect 26 17 31 30
rect 33 28 41 30
rect 33 26 36 28
rect 38 26 41 28
rect 33 21 41 26
rect 33 19 36 21
rect 38 19 41 21
rect 33 17 41 19
<< pdif >>
rect 6 56 14 58
rect 6 54 9 56
rect 11 54 14 56
rect 6 42 14 54
rect 16 53 24 58
rect 16 51 19 53
rect 21 51 24 53
rect 16 46 24 51
rect 16 44 19 46
rect 21 44 24 46
rect 16 42 24 44
rect 26 56 35 58
rect 26 54 29 56
rect 31 54 35 56
rect 26 42 35 54
rect 37 53 45 58
rect 37 51 40 53
rect 42 51 45 53
rect 37 46 45 51
rect 37 44 40 46
rect 42 44 45 46
rect 37 42 45 44
rect 47 56 54 58
rect 47 54 50 56
rect 52 54 54 56
rect 47 49 54 54
rect 47 47 50 49
rect 52 47 54 49
rect 47 42 54 47
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 18 53 22 55
rect 18 51 19 53
rect 21 51 22 53
rect 39 53 43 55
rect 2 39 6 47
rect 18 46 22 51
rect 39 51 40 53
rect 42 51 43 53
rect 39 46 43 51
rect 18 44 19 46
rect 21 44 40 46
rect 42 44 43 46
rect 18 42 43 44
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 18 28 22 42
rect 41 37 54 38
rect 41 35 43 37
rect 45 35 54 37
rect 41 34 54 35
rect 18 26 19 28
rect 21 26 22 28
rect 18 21 22 26
rect 18 19 19 21
rect 21 19 22 21
rect 18 17 22 19
rect 50 25 54 34
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 24 17 26 30
rect 31 17 33 30
<< pmos >>
rect 14 42 16 58
rect 24 42 26 58
rect 35 42 37 58
rect 45 42 47 58
<< polyct1 >>
rect 11 35 13 37
rect 43 35 45 37
<< ndifct0 >>
rect 36 26 38 28
rect 36 19 38 21
<< ndifct1 >>
rect 19 26 21 28
rect 19 19 21 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 9 54 11 56
rect 29 54 31 56
rect 50 54 52 56
rect 50 47 52 49
<< pdifct1 >>
rect 19 51 21 53
rect 19 44 21 46
rect 40 51 42 53
rect 40 44 42 46
<< alu0 >>
rect 8 56 12 68
rect 8 54 9 56
rect 11 54 12 56
rect 28 56 32 68
rect 8 52 12 54
rect 28 54 29 56
rect 31 54 32 56
rect 49 56 53 68
rect 28 52 32 54
rect 49 54 50 56
rect 52 54 53 56
rect 49 49 53 54
rect 49 47 50 49
rect 52 47 53 49
rect 49 45 53 47
rect 35 28 39 30
rect 35 26 36 28
rect 38 26 39 28
rect 35 21 39 26
rect 35 19 36 21
rect 38 19 39 21
rect 35 12 39 19
<< labels >>
rlabel alu1 4 40 4 40 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 36 20 36 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 44 36 44 6 z
rlabel alu1 28 44 28 44 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 36 44 36 6 a
rlabel alu1 52 28 52 28 6 a
<< end >>
