magic
tech scmos
timestamp 1199973108
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -5 40 101 97
<< pwell >>
rect -5 -9 101 40
<< poly >>
rect 2 81 11 83
rect 2 79 7 81
rect 9 79 11 81
rect 2 77 11 79
rect 9 74 11 77
rect 21 81 30 83
rect 21 79 26 81
rect 28 79 30 81
rect 21 77 30 79
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 81 75 83
rect 66 79 68 81
rect 70 79 75 81
rect 66 77 75 79
rect 53 74 55 77
rect 73 74 75 77
rect 85 77 94 83
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 37 14 43
rect 18 41 30 43
rect 18 39 20 41
rect 22 39 30 41
rect 18 37 30 39
rect 34 41 46 43
rect 34 39 36 41
rect 38 39 46 41
rect 34 37 46 39
rect 50 41 62 43
rect 50 39 56 41
rect 58 39 62 41
rect 50 37 62 39
rect 66 37 78 43
rect 82 41 94 43
rect 82 39 87 41
rect 89 39 94 41
rect 82 37 94 39
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 5 62 11
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndif >>
rect 2 14 9 34
rect 11 25 21 34
rect 11 23 15 25
rect 17 23 21 25
rect 11 18 21 23
rect 11 16 15 18
rect 17 16 21 18
rect 11 14 21 16
rect 23 32 30 34
rect 23 30 26 32
rect 28 30 30 32
rect 23 25 30 30
rect 23 23 26 25
rect 28 23 30 25
rect 23 14 30 23
rect 34 26 41 34
rect 34 24 36 26
rect 38 24 41 26
rect 34 18 41 24
rect 34 16 36 18
rect 38 16 41 18
rect 34 14 41 16
rect 43 14 53 34
rect 55 18 62 34
rect 55 16 58 18
rect 60 16 62 18
rect 55 14 62 16
rect 66 28 73 34
rect 66 26 68 28
rect 70 26 73 28
rect 66 21 73 26
rect 66 19 68 21
rect 70 19 73 21
rect 66 14 73 19
rect 75 32 85 34
rect 75 30 79 32
rect 81 30 85 32
rect 75 25 85 30
rect 75 23 79 25
rect 81 23 85 25
rect 75 14 85 23
rect 87 25 94 34
rect 87 23 90 25
rect 92 23 94 25
rect 87 18 94 23
rect 87 16 90 18
rect 92 16 94 18
rect 87 14 94 16
rect 13 2 19 14
rect 45 2 51 14
rect 77 2 83 14
<< pdif >>
rect 13 74 19 86
rect 45 74 51 86
rect 77 76 83 86
rect 77 74 79 76
rect 81 74 83 76
rect 2 46 9 74
rect 11 72 21 74
rect 11 70 15 72
rect 17 70 21 72
rect 11 65 21 70
rect 11 63 15 65
rect 17 63 21 65
rect 11 46 21 63
rect 23 61 30 74
rect 23 59 26 61
rect 28 59 30 61
rect 23 54 30 59
rect 23 52 26 54
rect 28 52 30 54
rect 23 46 30 52
rect 34 61 41 74
rect 34 59 36 61
rect 38 59 41 61
rect 34 46 41 59
rect 43 50 53 74
rect 43 48 47 50
rect 49 48 53 50
rect 43 46 53 48
rect 55 69 62 74
rect 55 67 58 69
rect 60 67 62 69
rect 55 46 62 67
rect 66 68 73 74
rect 66 66 68 68
rect 70 66 73 68
rect 66 61 73 66
rect 66 59 68 61
rect 70 59 73 61
rect 66 46 73 59
rect 75 69 85 74
rect 75 67 79 69
rect 81 67 85 69
rect 75 46 85 67
rect 87 69 94 74
rect 87 67 90 69
rect 92 67 94 69
rect 87 62 94 67
rect 87 60 90 62
rect 92 60 94 62
rect 87 46 94 60
<< alu1 >>
rect -2 89 98 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 73 87 87 89
rect 89 87 91 89
rect 93 87 98 89
rect -2 86 98 87
rect 6 81 10 86
rect 6 79 7 81
rect 9 79 10 81
rect 6 77 10 79
rect 14 81 18 86
rect 14 79 15 81
rect 17 79 18 81
rect 14 72 18 79
rect 78 81 82 86
rect 78 79 79 81
rect 81 79 82 81
rect 14 70 15 72
rect 17 70 18 72
rect 78 76 82 79
rect 78 74 79 76
rect 81 74 82 76
rect 14 65 18 70
rect 14 63 15 65
rect 17 63 18 65
rect 14 61 18 63
rect 14 33 18 55
rect 46 50 50 55
rect 46 48 47 50
rect 49 48 50 50
rect 14 25 18 27
rect 14 23 15 25
rect 17 23 18 25
rect 14 18 18 23
rect 46 30 50 48
rect 78 69 82 74
rect 78 67 79 69
rect 81 67 82 69
rect 78 65 82 67
rect 86 41 90 55
rect 86 39 87 41
rect 89 39 90 41
rect 86 33 90 39
rect 46 28 71 30
rect 46 27 68 28
rect 34 26 68 27
rect 70 26 71 28
rect 34 24 36 26
rect 38 24 50 26
rect 34 23 50 24
rect 38 19 42 23
rect 67 21 71 26
rect 89 25 93 27
rect 89 23 90 25
rect 92 23 93 25
rect 14 16 15 18
rect 17 16 18 18
rect 14 9 18 16
rect 34 18 42 19
rect 34 16 36 18
rect 38 16 42 18
rect 34 15 42 16
rect 57 18 61 20
rect 57 16 58 18
rect 60 16 61 18
rect 67 19 68 21
rect 70 19 71 21
rect 67 17 71 19
rect 89 18 93 23
rect 14 7 15 9
rect 17 7 18 9
rect 14 2 18 7
rect 57 9 61 16
rect 57 7 58 9
rect 60 7 61 9
rect 57 2 61 7
rect 89 16 90 18
rect 92 16 93 18
rect 89 9 93 16
rect 89 7 90 9
rect 92 7 93 9
rect 89 2 93 7
rect -2 1 98 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 73 -1 87 1
rect 89 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< alu2 >>
rect -2 89 98 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 71 89
rect 73 87 87 89
rect 89 87 98 89
rect -2 81 98 87
rect -2 79 15 81
rect 17 79 79 81
rect 81 79 98 81
rect -2 76 98 79
rect -2 9 98 12
rect -2 7 15 9
rect 17 7 58 9
rect 60 7 90 9
rect 92 7 98 9
rect -2 1 98 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 71 1
rect 73 -1 87 1
rect 89 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 71 3
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 57 -3 71 -1
rect 89 1 96 3
rect 89 -1 91 1
rect 93 -1 96 1
rect 89 -3 96 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 71 91
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 57 85 71 87
rect 89 89 96 91
rect 89 87 91 89
rect 93 87 96 89
rect 89 85 96 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polyct0 >>
rect 26 79 28 81
rect 68 79 70 81
rect 20 39 22 41
rect 36 39 38 41
rect 56 39 58 41
<< polyct1 >>
rect 7 79 9 81
rect 87 39 89 41
<< ndifct0 >>
rect 26 30 28 32
rect 26 23 28 25
rect 79 30 81 32
rect 79 23 81 25
<< ndifct1 >>
rect 15 23 17 25
rect 15 16 17 18
rect 36 24 38 26
rect 36 16 38 18
rect 58 16 60 18
rect 68 26 70 28
rect 68 19 70 21
rect 90 23 92 25
rect 90 16 92 18
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
rect 67 87 69 89
rect 91 87 93 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 91 -1 93 1
<< pdifct0 >>
rect 26 59 28 61
rect 26 52 28 54
rect 36 59 38 61
rect 58 67 60 69
rect 68 66 70 68
rect 68 59 70 61
rect 90 67 92 69
rect 90 60 92 62
<< pdifct1 >>
rect 79 74 81 76
rect 15 70 17 72
rect 15 63 17 65
rect 47 48 49 50
rect 79 67 81 69
<< alu0 >>
rect 24 81 72 82
rect 24 79 26 81
rect 28 79 68 81
rect 70 79 72 81
rect 24 78 72 79
rect 25 69 71 70
rect 25 67 58 69
rect 60 68 71 69
rect 60 67 68 68
rect 25 66 68 67
rect 70 66 71 68
rect 25 61 29 66
rect 25 59 26 61
rect 28 59 29 61
rect 25 54 29 59
rect 34 61 58 62
rect 34 59 36 61
rect 38 59 58 61
rect 34 58 58 59
rect 25 52 26 54
rect 28 52 39 54
rect 25 50 39 52
rect 18 41 24 42
rect 18 39 20 41
rect 22 39 24 41
rect 18 38 24 39
rect 35 41 39 50
rect 35 39 36 41
rect 38 39 39 41
rect 35 35 39 39
rect 25 32 39 35
rect 25 30 26 32
rect 28 31 39 32
rect 28 30 29 31
rect 25 25 29 30
rect 54 42 58 58
rect 67 61 71 66
rect 89 69 93 71
rect 89 67 90 69
rect 92 67 93 69
rect 89 62 93 67
rect 67 59 68 61
rect 70 59 71 61
rect 67 57 71 59
rect 78 60 90 62
rect 92 60 93 62
rect 78 58 93 60
rect 78 42 82 58
rect 54 41 82 42
rect 54 39 56 41
rect 58 39 82 41
rect 54 38 82 39
rect 78 32 82 38
rect 78 30 79 32
rect 81 30 82 32
rect 25 23 26 25
rect 28 23 29 25
rect 25 21 29 23
rect 78 25 82 30
rect 78 23 79 25
rect 81 23 82 25
rect 78 21 82 23
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 71 87 73 89
rect 87 87 89 89
rect 15 79 17 81
rect 79 79 81 81
rect 15 7 17 9
rect 58 7 60 9
rect 90 7 92 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
rect 71 -1 73 1
rect 87 -1 89 1
<< labels >>
rlabel alu1 16 44 16 44 6 b
rlabel alu1 40 20 40 20 6 z
rlabel alu1 48 40 48 40 6 z
rlabel alu1 64 28 64 28 6 z
rlabel alu1 56 28 56 28 6 z
rlabel alu1 88 44 88 44 6 a
rlabel alu2 48 6 48 6 6 vss
rlabel alu2 48 82 48 82 6 vdd
<< end >>
