magic
tech scmos
timestamp 1199202888
<< ab >>
rect 0 0 136 80
<< nwell >>
rect -5 36 141 88
<< pwell >>
rect -5 -8 141 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 84 70 86 74
rect 94 70 96 74
rect 101 70 103 74
rect 111 70 113 74
rect 121 61 123 65
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 67 39 69 42
rect 77 39 79 42
rect 16 37 29 39
rect 33 37 45 39
rect 23 35 25 37
rect 27 35 29 37
rect 23 33 29 35
rect 9 31 19 33
rect 13 29 15 31
rect 17 29 19 31
rect 13 27 19 29
rect 17 24 19 27
rect 27 24 29 33
rect 39 35 41 37
rect 43 35 45 37
rect 39 33 45 35
rect 49 37 63 39
rect 49 35 51 37
rect 53 35 63 37
rect 49 33 63 35
rect 67 37 79 39
rect 84 39 86 42
rect 94 39 96 42
rect 101 39 103 42
rect 111 39 113 42
rect 121 39 123 42
rect 84 37 96 39
rect 100 37 106 39
rect 67 35 69 37
rect 71 35 73 37
rect 67 33 73 35
rect 84 35 86 37
rect 88 35 90 37
rect 84 33 90 35
rect 100 35 102 37
rect 104 35 106 37
rect 100 33 106 35
rect 110 37 123 39
rect 110 35 116 37
rect 118 35 123 37
rect 110 33 123 35
rect 39 30 41 33
rect 49 30 51 33
rect 61 30 63 33
rect 71 30 73 33
rect 110 27 112 33
rect 120 27 122 33
rect 17 8 19 13
rect 27 8 29 13
rect 39 8 41 13
rect 49 8 51 13
rect 61 8 63 13
rect 71 8 73 13
rect 110 10 112 15
rect 120 10 122 15
<< ndif >>
rect 31 24 39 30
rect 8 13 17 24
rect 19 21 27 24
rect 19 19 22 21
rect 24 19 27 21
rect 19 13 27 19
rect 29 13 39 24
rect 41 21 49 30
rect 41 19 44 21
rect 46 19 49 21
rect 41 13 49 19
rect 51 13 61 30
rect 63 21 71 30
rect 63 19 66 21
rect 68 19 71 21
rect 63 13 71 19
rect 73 17 81 30
rect 73 15 76 17
rect 78 15 81 17
rect 103 19 110 27
rect 103 17 105 19
rect 107 17 110 19
rect 103 15 110 17
rect 112 25 120 27
rect 112 23 115 25
rect 117 23 120 25
rect 112 15 120 23
rect 122 19 130 27
rect 122 17 125 19
rect 127 17 130 19
rect 122 15 130 17
rect 73 13 81 15
rect 8 11 15 13
rect 8 9 11 11
rect 13 9 15 11
rect 8 7 15 9
rect 31 11 37 13
rect 31 9 33 11
rect 35 9 37 11
rect 31 7 37 9
rect 53 11 59 13
rect 53 9 55 11
rect 57 9 59 11
rect 53 7 59 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 42 16 70
rect 18 61 26 70
rect 18 59 21 61
rect 23 59 26 61
rect 18 53 26 59
rect 18 51 21 53
rect 23 51 26 53
rect 18 42 26 51
rect 28 42 33 70
rect 35 68 43 70
rect 35 66 38 68
rect 40 66 43 68
rect 35 61 43 66
rect 35 59 38 61
rect 40 59 43 61
rect 35 42 43 59
rect 45 42 50 70
rect 52 60 60 70
rect 52 58 55 60
rect 57 58 60 60
rect 52 53 60 58
rect 52 51 55 53
rect 57 51 60 53
rect 52 42 60 51
rect 62 42 67 70
rect 69 68 77 70
rect 69 66 72 68
rect 74 66 77 68
rect 69 61 77 66
rect 69 59 72 61
rect 74 59 77 61
rect 69 42 77 59
rect 79 42 84 70
rect 86 61 94 70
rect 86 59 89 61
rect 91 59 94 61
rect 86 53 94 59
rect 86 51 89 53
rect 91 51 94 53
rect 86 42 94 51
rect 96 42 101 70
rect 103 68 111 70
rect 103 66 106 68
rect 108 66 111 68
rect 103 61 111 66
rect 103 59 106 61
rect 108 59 111 61
rect 103 54 111 59
rect 103 52 106 54
rect 108 52 111 54
rect 103 42 111 52
rect 113 61 118 70
rect 113 53 121 61
rect 113 51 116 53
rect 118 51 121 53
rect 113 46 121 51
rect 113 44 116 46
rect 118 44 121 46
rect 113 42 121 44
rect 123 59 130 61
rect 123 57 126 59
rect 128 57 130 59
rect 123 52 130 57
rect 123 50 126 52
rect 128 50 130 52
rect 123 42 130 50
<< alu1 >>
rect -2 81 138 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 138 81
rect -2 68 138 79
rect 18 61 24 63
rect 18 59 21 61
rect 23 59 24 61
rect 18 54 24 59
rect 88 61 94 63
rect 88 59 89 61
rect 91 59 94 61
rect 88 54 94 59
rect 2 53 94 54
rect 2 51 21 53
rect 23 51 55 53
rect 57 51 89 53
rect 91 51 94 53
rect 2 50 94 51
rect 2 22 6 50
rect 25 42 87 46
rect 25 38 31 42
rect 23 37 31 38
rect 23 35 25 37
rect 27 35 31 37
rect 23 34 31 35
rect 49 37 55 42
rect 81 38 87 42
rect 49 35 51 37
rect 53 35 55 37
rect 49 34 55 35
rect 81 37 95 38
rect 81 35 86 37
rect 88 35 95 37
rect 81 34 95 35
rect 113 37 127 38
rect 113 35 116 37
rect 118 35 127 37
rect 113 34 127 35
rect 122 25 127 34
rect 2 21 71 22
rect 2 19 22 21
rect 24 19 44 21
rect 46 19 66 21
rect 68 19 71 21
rect 2 18 71 19
rect -2 11 138 12
rect -2 9 11 11
rect 13 9 33 11
rect 35 9 55 11
rect 57 9 138 11
rect -2 1 138 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 138 1
rect -2 -2 138 -1
<< ptie >>
rect 0 1 136 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 136 1
rect 0 -3 136 -1
<< ntie >>
rect 0 81 136 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 136 81
rect 0 77 136 79
<< nmos >>
rect 17 13 19 24
rect 27 13 29 24
rect 39 13 41 30
rect 49 13 51 30
rect 61 13 63 30
rect 71 13 73 30
rect 110 15 112 27
rect 120 15 122 27
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 84 42 86 70
rect 94 42 96 70
rect 101 42 103 70
rect 111 42 113 70
rect 121 42 123 61
<< polyct0 >>
rect 15 29 17 31
rect 41 35 43 37
rect 69 35 71 37
rect 102 35 104 37
<< polyct1 >>
rect 25 35 27 37
rect 51 35 53 37
rect 86 35 88 37
rect 116 35 118 37
<< ndifct0 >>
rect 76 15 78 17
rect 105 17 107 19
rect 115 23 117 25
rect 125 17 127 19
<< ndifct1 >>
rect 22 19 24 21
rect 44 19 46 21
rect 66 19 68 21
rect 11 9 13 11
rect 33 9 35 11
rect 55 9 57 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 38 66 40 68
rect 38 59 40 61
rect 55 58 57 60
rect 72 66 74 68
rect 72 59 74 61
rect 106 66 108 68
rect 106 59 108 61
rect 106 52 108 54
rect 116 51 118 53
rect 116 44 118 46
rect 126 57 128 59
rect 126 50 128 52
<< pdifct1 >>
rect 21 59 23 61
rect 21 51 23 53
rect 55 51 57 53
rect 89 59 91 61
rect 89 51 91 53
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 36 66 38 68
rect 40 66 42 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 36 61 42 66
rect 70 66 72 68
rect 74 66 76 68
rect 36 59 38 61
rect 40 59 42 61
rect 36 58 42 59
rect 54 60 58 62
rect 54 58 55 60
rect 57 58 58 60
rect 70 61 76 66
rect 105 66 106 68
rect 108 66 109 68
rect 70 59 72 61
rect 74 59 76 61
rect 70 58 76 59
rect 54 54 58 58
rect 105 61 109 66
rect 105 59 106 61
rect 108 59 109 61
rect 105 54 109 59
rect 124 59 130 68
rect 124 57 126 59
rect 128 57 130 59
rect 105 52 106 54
rect 108 52 109 54
rect 105 50 109 52
rect 115 53 119 55
rect 115 51 116 53
rect 118 51 119 53
rect 115 46 119 51
rect 124 52 130 57
rect 124 50 126 52
rect 128 50 130 52
rect 124 49 130 50
rect 39 37 45 38
rect 39 35 41 37
rect 43 35 45 37
rect 14 31 18 33
rect 14 29 15 31
rect 17 30 18 31
rect 39 30 45 35
rect 101 44 116 46
rect 118 44 119 46
rect 101 42 119 44
rect 67 37 73 38
rect 67 35 69 37
rect 71 35 73 37
rect 67 30 73 35
rect 101 37 105 42
rect 101 35 102 37
rect 104 35 105 37
rect 101 30 105 35
rect 17 29 118 30
rect 14 26 118 29
rect 114 25 118 26
rect 114 23 115 25
rect 117 23 118 25
rect 114 21 118 23
rect 104 19 108 21
rect 75 17 79 19
rect 75 15 76 17
rect 78 15 79 17
rect 75 12 79 15
rect 104 17 105 19
rect 107 17 108 19
rect 104 12 108 17
rect 124 19 128 21
rect 124 17 125 19
rect 127 17 128 19
rect 124 12 128 17
<< labels >>
rlabel alu0 42 32 42 32 6 an
rlabel alu0 70 32 70 32 6 an
rlabel polyct0 103 36 103 36 6 an
rlabel alu0 66 28 66 28 6 an
rlabel alu0 116 25 116 25 6 an
rlabel alu0 117 48 117 48 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 44 20 44 20 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 68 6 68 6 6 vss
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 52 40 52 40 6 b
rlabel alu1 60 44 60 44 6 b
rlabel alu1 68 44 68 44 6 b
rlabel alu1 76 44 76 44 6 b
rlabel alu1 60 52 60 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 68 74 68 74 6 vdd
rlabel alu1 84 40 84 40 6 b
rlabel alu1 92 36 92 36 6 b
rlabel alu1 84 52 84 52 6 z
rlabel alu1 92 60 92 60 6 z
rlabel alu1 124 32 124 32 6 a
rlabel alu1 116 36 116 36 6 a
<< end >>
