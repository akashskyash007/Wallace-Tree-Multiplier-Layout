magic
tech scmos
timestamp 1199201678
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 19 67 21 72
rect 29 67 31 72
rect 9 39 11 42
rect 19 39 21 50
rect 29 47 31 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 30 11 33
rect 22 30 24 33
rect 29 30 31 41
rect 9 11 11 16
rect 22 11 24 16
rect 29 11 31 16
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 20 9 26
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 22 30
rect 24 16 29 30
rect 31 22 36 30
rect 31 20 38 22
rect 31 18 34 20
rect 36 18 38 20
rect 31 16 38 18
rect 13 11 20 16
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 67 17 70
rect 11 65 19 67
rect 11 63 14 65
rect 16 63 19 65
rect 11 50 19 63
rect 21 61 29 67
rect 21 59 24 61
rect 26 59 29 61
rect 21 54 29 59
rect 21 52 24 54
rect 26 52 29 54
rect 21 50 29 52
rect 31 65 38 67
rect 31 63 34 65
rect 36 63 38 65
rect 31 50 38 63
rect 11 42 17 50
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 61 7 63
rect 2 59 4 61
rect 6 59 7 61
rect 2 54 7 59
rect 2 52 4 54
rect 6 52 7 54
rect 2 50 7 52
rect 2 28 6 50
rect 34 46 38 55
rect 25 45 38 46
rect 25 43 31 45
rect 33 43 38 45
rect 25 42 38 43
rect 17 37 31 38
rect 17 35 21 37
rect 23 35 31 37
rect 17 34 31 35
rect 2 26 4 28
rect 2 23 6 26
rect 2 20 14 23
rect 2 18 4 20
rect 6 18 14 20
rect 2 17 14 18
rect 26 25 31 34
rect -2 11 42 12
rect -2 9 15 11
rect 17 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 16 11 30
rect 22 16 24 30
rect 29 16 31 30
<< pmos >>
rect 9 42 11 70
rect 19 50 21 67
rect 29 50 31 67
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 21 35 23 37
<< ndifct0 >>
rect 34 18 36 20
<< ndifct1 >>
rect 4 26 6 28
rect 4 18 6 20
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 63 16 65
rect 24 59 26 61
rect 24 52 26 54
rect 34 63 36 65
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
<< alu0 >>
rect 13 65 17 68
rect 13 63 14 65
rect 16 63 17 65
rect 33 65 37 68
rect 33 63 34 65
rect 36 63 37 65
rect 13 61 17 63
rect 23 61 27 63
rect 33 61 37 63
rect 23 59 24 61
rect 26 59 27 61
rect 23 54 27 59
rect 10 52 24 54
rect 26 52 27 54
rect 10 50 27 52
rect 10 37 14 50
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 6 23 7 30
rect 10 26 22 30
rect 18 21 22 26
rect 18 20 38 21
rect 18 18 34 20
rect 36 18 38 20
rect 18 17 38 18
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 25 56 25 56 6 zn
rlabel alu0 28 19 28 19 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 52 36 52 6 b
<< end >>
