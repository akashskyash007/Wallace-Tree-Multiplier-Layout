magic
tech scmos
timestamp 1199203321
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 66 11 70
rect 28 66 30 70
rect 35 66 37 70
rect 42 66 44 70
rect 49 66 51 70
rect 9 35 11 38
rect 28 35 30 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 30 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 9 20 11 29
rect 20 18 22 29
rect 35 27 37 38
rect 30 25 37 27
rect 30 23 33 25
rect 35 23 37 25
rect 30 21 37 23
rect 42 27 44 38
rect 49 35 51 38
rect 49 33 59 35
rect 52 31 55 33
rect 57 31 59 33
rect 52 29 59 31
rect 42 25 48 27
rect 42 23 44 25
rect 46 23 48 25
rect 42 21 48 23
rect 30 18 32 21
rect 42 18 44 21
rect 52 18 54 29
rect 9 2 11 6
rect 20 5 22 10
rect 30 5 32 10
rect 42 5 44 10
rect 52 5 54 10
<< ndif >>
rect 2 18 9 20
rect 2 16 4 18
rect 6 16 9 18
rect 2 14 9 16
rect 4 6 9 14
rect 11 18 18 20
rect 11 17 20 18
rect 11 15 14 17
rect 16 15 20 17
rect 11 10 20 15
rect 22 16 30 18
rect 22 14 25 16
rect 27 14 30 16
rect 22 10 30 14
rect 32 10 42 18
rect 44 16 52 18
rect 44 14 47 16
rect 49 14 52 16
rect 44 10 52 14
rect 54 10 62 18
rect 11 8 14 10
rect 16 8 18 10
rect 11 6 18 8
rect 34 7 40 10
rect 34 5 36 7
rect 38 5 40 7
rect 56 7 62 10
rect 56 5 58 7
rect 60 5 62 7
rect 34 3 40 5
rect 56 3 62 5
<< pdif >>
rect 13 66 19 68
rect 4 52 9 66
rect 2 50 9 52
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 4 38 9 46
rect 11 65 19 66
rect 11 63 15 65
rect 17 63 19 65
rect 11 55 19 63
rect 11 38 17 55
rect 23 51 28 66
rect 21 49 28 51
rect 21 47 23 49
rect 25 47 28 49
rect 21 45 28 47
rect 23 38 28 45
rect 30 38 35 66
rect 37 38 42 66
rect 44 38 49 66
rect 51 64 59 66
rect 51 62 54 64
rect 56 62 59 64
rect 51 57 59 62
rect 51 55 54 57
rect 56 55 59 57
rect 51 38 59 55
<< alu1 >>
rect -2 65 66 72
rect -2 64 15 65
rect 17 64 66 65
rect 2 53 14 59
rect 2 50 6 53
rect 2 48 4 50
rect 2 20 6 48
rect 34 42 38 59
rect 19 38 38 42
rect 42 42 46 51
rect 42 38 59 42
rect 19 33 25 38
rect 19 31 21 33
rect 23 31 25 33
rect 19 30 25 31
rect 32 30 47 34
rect 53 33 59 38
rect 53 31 55 33
rect 57 31 59 33
rect 53 30 59 31
rect 2 18 7 20
rect 2 16 4 18
rect 6 16 7 18
rect 2 13 7 16
rect 32 25 38 30
rect 32 23 33 25
rect 35 23 38 25
rect 32 21 38 23
rect 42 25 62 26
rect 42 23 44 25
rect 46 23 62 25
rect 42 22 62 23
rect 58 13 62 22
rect -2 7 66 8
rect -2 5 36 7
rect 38 5 58 7
rect 60 5 66 7
rect -2 0 66 5
<< nmos >>
rect 9 6 11 20
rect 20 10 22 18
rect 30 10 32 18
rect 42 10 44 18
rect 52 10 54 18
<< pmos >>
rect 9 38 11 66
rect 28 38 30 66
rect 35 38 37 66
rect 42 38 44 66
rect 49 38 51 66
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 21 31 23 33
rect 33 23 35 25
rect 55 31 57 33
rect 44 23 46 25
<< ndifct0 >>
rect 14 15 16 17
rect 25 14 27 16
rect 47 14 49 16
rect 14 8 16 10
<< ndifct1 >>
rect 4 16 6 18
rect 36 5 38 7
rect 58 5 60 7
<< pdifct0 >>
rect 15 63 17 64
rect 23 47 25 49
rect 54 62 56 64
rect 54 55 56 57
<< pdifct1 >>
rect 4 48 6 50
rect 15 64 17 65
<< alu0 >>
rect 13 63 15 64
rect 17 63 19 64
rect 13 62 19 63
rect 52 62 54 64
rect 56 62 58 64
rect 6 46 7 53
rect 11 49 27 50
rect 11 47 23 49
rect 25 47 27 49
rect 11 46 27 47
rect 11 35 15 46
rect 52 57 58 62
rect 52 55 54 57
rect 56 55 58 57
rect 52 54 58 55
rect 10 33 15 35
rect 10 31 11 33
rect 13 31 15 33
rect 10 29 15 31
rect 11 26 15 29
rect 11 22 27 26
rect 12 17 18 18
rect 12 15 14 17
rect 16 15 18 17
rect 12 10 18 15
rect 23 17 27 22
rect 23 16 51 17
rect 23 14 25 16
rect 27 14 47 16
rect 49 14 51 16
rect 23 13 51 14
rect 12 8 14 10
rect 16 8 18 10
<< labels >>
rlabel alu0 13 36 13 36 6 zn
rlabel alu0 19 48 19 48 6 zn
rlabel alu0 37 15 37 15 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 40 28 40 6 d
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 28 36 28 6 c
rlabel alu1 44 32 44 32 6 c
rlabel alu1 36 52 36 52 6 d
rlabel alu1 44 48 44 48 6 a
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 60 16 60 16 6 b
rlabel alu1 52 24 52 24 6 b
rlabel alu1 52 40 52 40 6 a
<< end >>
