magic
tech scmos
timestamp 1199475724
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< alu1 >>
rect -2 96 72 102
rect -2 94 49 96
rect 51 94 72 96
rect -2 88 72 94
rect -2 6 72 12
rect -2 4 19 6
rect 21 4 72 6
rect -2 -2 72 4
<< alu2 >>
rect 7 96 63 102
rect 7 94 19 96
rect 21 94 49 96
rect 51 94 63 96
rect 7 88 63 94
rect 7 6 63 12
rect 7 4 19 6
rect 21 4 49 6
rect 51 4 63 6
rect 7 -2 63 4
<< alu3 >>
rect 8 96 32 102
rect 8 94 19 96
rect 21 94 32 96
rect 8 -2 32 94
rect 38 6 62 102
rect 38 4 49 6
rect 51 4 62 6
rect 38 -2 62 4
<< via1 >>
rect 49 94 51 96
rect 19 4 21 6
<< via2 >>
rect 19 94 21 96
rect 49 4 51 6
<< labels >>
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 35 94 35 94 6 vdd
rlabel alu2 35 6 35 6 6 vss
rlabel alu2 35 94 35 94 6 vdd
rlabel alu3 20 50 20 50 6 vdd
rlabel alu3 50 50 50 50 6 vss
<< end >>
