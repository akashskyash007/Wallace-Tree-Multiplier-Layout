magic
tech scmos
timestamp 1199202528
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 22 68 24 73
rect 32 68 34 73
rect 45 70 47 74
rect 9 61 11 65
rect 45 49 47 52
rect 41 47 47 49
rect 41 45 43 47
rect 45 45 47 47
rect 9 31 11 43
rect 22 41 24 44
rect 16 39 24 41
rect 32 41 34 44
rect 41 43 47 45
rect 32 39 37 41
rect 16 37 18 39
rect 20 37 24 39
rect 16 35 24 37
rect 35 37 41 39
rect 35 35 37 37
rect 39 35 41 37
rect 22 33 30 35
rect 9 29 16 31
rect 28 30 30 33
rect 35 33 41 35
rect 35 30 37 33
rect 45 30 47 43
rect 9 27 12 29
rect 14 27 16 29
rect 9 25 16 27
rect 9 22 11 25
rect 9 8 11 13
rect 45 16 47 21
rect 28 6 30 10
rect 35 6 37 10
<< ndif >>
rect 21 28 28 30
rect 21 26 23 28
rect 25 26 28 28
rect 21 24 28 26
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 4 13 9 16
rect 11 20 17 22
rect 11 13 19 20
rect 13 11 19 13
rect 13 9 15 11
rect 17 9 19 11
rect 23 10 28 24
rect 30 10 35 30
rect 37 25 45 30
rect 37 23 40 25
rect 42 23 45 25
rect 37 21 45 23
rect 47 28 54 30
rect 47 26 50 28
rect 52 26 54 28
rect 47 24 54 26
rect 47 21 52 24
rect 37 10 43 21
rect 13 7 19 9
<< pdif >>
rect 36 68 45 70
rect 14 61 22 68
rect 4 56 9 61
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 59 16 61
rect 18 59 22 61
rect 11 44 22 59
rect 24 56 32 68
rect 24 54 27 56
rect 29 54 32 56
rect 24 48 32 54
rect 24 46 27 48
rect 29 46 32 48
rect 24 44 32 46
rect 34 66 38 68
rect 40 66 45 68
rect 34 61 45 66
rect 34 59 38 61
rect 40 59 45 61
rect 34 52 45 59
rect 47 58 52 70
rect 47 56 54 58
rect 47 54 50 56
rect 52 54 54 56
rect 47 52 54 54
rect 34 44 39 52
rect 11 43 16 44
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 26 56 30 58
rect 26 54 27 56
rect 29 54 30 56
rect 17 50 30 54
rect 26 48 30 50
rect 34 49 46 55
rect 26 46 27 48
rect 29 46 30 48
rect 9 29 18 30
rect 9 27 12 29
rect 14 27 18 29
rect 9 26 18 27
rect 14 22 18 26
rect 26 26 30 46
rect 42 47 46 49
rect 42 45 43 47
rect 45 45 46 47
rect 42 41 46 45
rect 14 18 31 22
rect -2 11 58 12
rect -2 9 15 11
rect 17 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 13 11 22
rect 28 10 30 30
rect 35 10 37 30
rect 45 21 47 30
<< pmos >>
rect 9 43 11 61
rect 22 44 24 68
rect 32 44 34 68
rect 45 52 47 70
<< polyct0 >>
rect 18 37 20 39
rect 37 35 39 37
<< polyct1 >>
rect 43 45 45 47
rect 12 27 14 29
<< ndifct0 >>
rect 23 26 25 28
rect 4 18 6 20
rect 40 23 42 25
rect 50 26 52 28
<< ndifct1 >>
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 52 6 54
rect 4 45 6 47
rect 16 59 18 61
rect 38 66 40 68
rect 38 59 40 61
rect 50 54 52 56
<< pdifct1 >>
rect 27 54 29 56
rect 27 46 29 48
<< alu0 >>
rect 14 61 20 68
rect 14 59 16 61
rect 18 59 20 61
rect 14 58 20 59
rect 36 66 38 68
rect 40 66 42 68
rect 36 61 42 66
rect 36 59 38 61
rect 40 59 42 61
rect 36 58 42 59
rect 3 54 7 56
rect 49 56 53 58
rect 3 52 4 54
rect 6 52 7 54
rect 3 47 7 52
rect 3 45 4 47
rect 6 45 7 47
rect 3 40 7 45
rect 2 39 22 40
rect 2 37 18 39
rect 20 37 22 39
rect 2 36 22 37
rect 2 21 6 36
rect 21 28 26 30
rect 21 26 23 28
rect 25 26 26 28
rect 49 54 50 56
rect 52 54 53 56
rect 49 38 53 54
rect 35 37 53 38
rect 35 35 37 37
rect 39 35 53 37
rect 35 34 53 35
rect 49 28 53 34
rect 21 25 27 26
rect 39 25 43 27
rect 39 23 40 25
rect 42 23 43 25
rect 49 26 50 28
rect 52 26 53 28
rect 49 24 53 26
rect 2 20 8 21
rect 2 18 4 20
rect 6 18 8 20
rect 2 17 8 18
rect 39 12 43 23
<< labels >>
rlabel pdifct0 5 46 5 46 6 bn
rlabel alu0 4 28 4 28 6 bn
rlabel alu0 12 38 12 38 6 bn
rlabel alu0 44 36 44 36 6 an
rlabel alu0 51 41 51 41 6 an
rlabel alu1 20 20 20 20 6 b
rlabel alu1 12 28 12 28 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 20 28 20 6 b
rlabel alu1 28 44 28 44 6 z
rlabel alu1 36 52 36 52 6 a
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 48 44 48 6 a
<< end >>
