magic
tech scmos
timestamp 1199201739
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 67 21 72
rect 29 67 31 72
rect 41 67 43 72
rect 19 47 21 58
rect 29 55 31 58
rect 29 53 37 55
rect 29 51 33 53
rect 35 51 37 53
rect 29 49 37 51
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 9 39 11 42
rect 19 41 25 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 30 11 33
rect 22 26 24 41
rect 29 26 31 49
rect 41 35 43 58
rect 40 33 46 35
rect 40 31 42 33
rect 44 31 46 33
rect 36 29 46 31
rect 36 26 38 29
rect 9 12 11 16
rect 22 12 24 17
rect 29 12 31 17
rect 36 12 38 17
<< ndif >>
rect 4 23 9 30
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 16 9 19
rect 11 26 20 30
rect 11 17 22 26
rect 24 17 29 26
rect 31 17 36 26
rect 38 23 43 26
rect 38 21 45 23
rect 38 19 41 21
rect 43 19 45 21
rect 38 17 45 19
rect 11 16 20 17
rect 13 11 20 16
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 67 16 70
rect 33 71 39 73
rect 33 69 35 71
rect 37 69 39 71
rect 33 67 39 69
rect 11 65 19 67
rect 11 63 14 65
rect 16 63 19 65
rect 11 58 19 63
rect 21 62 29 67
rect 21 60 24 62
rect 26 60 29 62
rect 21 58 29 60
rect 31 58 41 67
rect 43 64 48 67
rect 43 62 50 64
rect 43 60 46 62
rect 48 60 50 62
rect 43 58 50 60
rect 11 42 17 58
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 35 71
rect 37 69 58 71
rect -2 68 58 69
rect 2 53 7 63
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 31 53 47 54
rect 31 51 33 53
rect 35 51 47 53
rect 31 50 47 51
rect 2 22 6 42
rect 17 45 31 46
rect 17 43 21 45
rect 23 43 31 45
rect 17 42 31 43
rect 41 42 47 50
rect 25 34 31 42
rect 41 33 47 38
rect 41 31 42 33
rect 44 31 47 33
rect 41 30 47 31
rect 25 26 47 30
rect 2 21 15 22
rect 2 19 4 21
rect 6 19 15 21
rect 2 18 15 19
rect -2 11 58 12
rect -2 9 15 11
rect 17 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 16 11 30
rect 22 17 24 26
rect 29 17 31 26
rect 36 17 38 26
<< pmos >>
rect 9 42 11 70
rect 19 58 21 67
rect 29 58 31 67
rect 41 58 43 67
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 33 51 35 53
rect 21 43 23 45
rect 42 31 44 33
<< ndifct0 >>
rect 41 19 43 21
<< ndifct1 >>
rect 4 19 6 21
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 14 63 16 65
rect 24 60 26 62
rect 46 60 48 62
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 35 69 37 71
<< alu0 >>
rect 13 65 17 68
rect 13 63 14 65
rect 16 63 17 65
rect 13 61 17 63
rect 22 62 50 63
rect 22 60 24 62
rect 26 60 46 62
rect 48 60 50 62
rect 22 59 50 60
rect 22 54 26 59
rect 10 50 26 54
rect 10 37 14 50
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 10 26 22 30
rect 18 22 22 26
rect 18 21 45 22
rect 18 19 41 21
rect 43 19 45 21
rect 18 18 45 19
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 31 20 31 20 6 zn
rlabel alu0 36 61 36 61 6 zn
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 44 20 44 6 a
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 28 28 28 6 c
rlabel alu1 36 28 36 28 6 c
rlabel alu1 28 40 28 40 6 a
rlabel alu1 36 52 36 52 6 b
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 c
rlabel alu1 44 48 44 48 6 b
<< end >>
