magic
tech scmos
timestamp 1199980664
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -8 40 72 97
<< pwell >>
rect -8 -9 72 40
<< poly >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 2 36 17 38
rect 2 34 7 36
rect 9 34 17 36
rect 2 32 17 34
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 2 14 8
rect 18 2 27 8
rect 37 6 46 8
rect 37 4 42 6
rect 44 4 46 6
rect 37 2 46 4
rect 50 6 59 8
rect 50 4 52 6
rect 54 4 59 6
rect 50 2 59 4
<< ndif >>
rect 2 23 9 29
rect 2 21 4 23
rect 6 21 9 23
rect 2 16 9 21
rect 2 14 4 16
rect 6 14 9 16
rect 2 11 9 14
rect 11 24 21 29
rect 11 22 15 24
rect 17 22 21 24
rect 11 17 21 22
rect 11 15 15 17
rect 17 15 21 17
rect 11 11 21 15
rect 23 16 30 29
rect 23 14 26 16
rect 28 14 30 16
rect 23 11 30 14
rect 34 24 41 29
rect 34 22 36 24
rect 38 22 41 24
rect 34 17 41 22
rect 34 15 36 17
rect 38 15 41 17
rect 34 11 41 15
rect 43 25 53 29
rect 43 23 47 25
rect 49 23 53 25
rect 43 11 53 23
rect 55 16 62 29
rect 55 14 58 16
rect 60 14 62 16
rect 55 11 62 14
<< pdif >>
rect 2 74 9 77
rect 2 72 4 74
rect 6 72 9 74
rect 2 67 9 72
rect 2 65 4 67
rect 6 65 9 67
rect 2 51 9 65
rect 11 65 21 77
rect 11 63 15 65
rect 17 63 21 65
rect 11 57 21 63
rect 11 55 15 57
rect 17 55 21 57
rect 11 51 21 55
rect 23 74 30 77
rect 23 72 26 74
rect 28 72 30 74
rect 23 67 30 72
rect 23 65 26 67
rect 28 65 30 67
rect 23 51 30 65
rect 34 74 41 77
rect 34 72 36 74
rect 38 72 41 74
rect 34 67 41 72
rect 34 65 36 67
rect 38 65 41 67
rect 34 51 41 65
rect 43 65 53 77
rect 43 63 47 65
rect 49 63 53 65
rect 43 58 53 63
rect 43 56 47 58
rect 49 56 53 58
rect 43 51 53 56
rect 55 74 62 77
rect 55 72 58 74
rect 60 72 62 74
rect 55 67 62 72
rect 55 65 58 67
rect 60 65 62 67
rect 55 51 62 65
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect 62 85 66 90
rect -2 83 -1 85
rect 1 83 7 85
rect -2 81 7 83
rect 3 74 7 81
rect 3 72 4 74
rect 6 72 7 74
rect 3 67 7 72
rect 25 83 31 85
rect 33 83 39 85
rect 25 81 39 83
rect 25 74 29 81
rect 25 72 26 74
rect 28 72 29 74
rect 25 67 29 72
rect 3 65 4 67
rect 6 65 7 67
rect 3 63 7 65
rect 13 65 18 67
rect 13 63 15 65
rect 17 63 18 65
rect 25 65 26 67
rect 28 65 29 67
rect 25 63 29 65
rect 35 74 39 81
rect 35 72 36 74
rect 38 72 39 74
rect 35 67 39 72
rect 57 83 63 85
rect 65 83 66 85
rect 57 81 66 83
rect 57 74 61 81
rect 57 72 58 74
rect 60 72 61 74
rect 57 67 61 72
rect 35 65 36 67
rect 38 65 39 67
rect 35 63 39 65
rect 46 65 50 67
rect 46 63 47 65
rect 49 63 50 65
rect 57 65 58 67
rect 60 65 61 67
rect 57 63 61 65
rect 13 58 18 63
rect 46 58 50 63
rect 13 57 47 58
rect 13 55 15 57
rect 17 56 47 57
rect 49 56 50 58
rect 17 55 50 56
rect 13 54 50 55
rect 6 46 10 48
rect 6 44 7 46
rect 9 44 10 46
rect 6 36 10 44
rect 6 34 7 36
rect 9 34 10 36
rect 21 46 27 50
rect 21 44 23 46
rect 25 44 27 46
rect 21 36 27 44
rect 21 34 23 36
rect 25 34 27 36
rect 6 30 27 34
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 16 7 21
rect 3 14 4 16
rect 6 14 7 16
rect 3 7 7 14
rect 25 16 29 18
rect 25 14 26 16
rect 28 14 29 16
rect 25 7 29 14
rect 46 25 50 54
rect 54 46 58 59
rect 54 44 55 46
rect 57 44 58 46
rect 54 36 58 44
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 46 23 47 25
rect 49 23 50 25
rect 46 21 50 23
rect -2 5 34 7
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 34 5
rect 62 5 66 7
rect 62 3 63 5
rect 65 3 66 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 -2 66 3
<< alu2 >>
rect -2 85 66 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 66 85
rect -2 80 66 83
rect -2 5 66 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 66 5
rect -2 -2 66 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polyct0 >>
rect 39 44 41 46
rect 39 34 41 36
rect 42 4 44 6
rect 52 4 54 6
<< polyct1 >>
rect 7 44 9 46
rect 23 44 25 46
rect 55 44 57 46
rect 7 34 9 36
rect 23 34 25 36
rect 55 34 57 36
<< ndifct0 >>
rect 15 22 17 24
rect 15 15 17 17
rect 36 22 38 24
rect 36 15 38 17
rect 58 14 60 16
<< ndifct1 >>
rect 4 21 6 23
rect 4 14 6 16
rect 26 14 28 16
rect 47 23 49 25
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< pdifct1 >>
rect 4 72 6 74
rect 4 65 6 67
rect 15 63 17 65
rect 15 55 17 57
rect 26 72 28 74
rect 26 65 28 67
rect 36 72 38 74
rect 36 65 38 67
rect 47 63 49 65
rect 47 56 49 58
rect 58 72 60 74
rect 58 65 60 67
<< alu0 >>
rect 38 46 42 48
rect 38 44 39 46
rect 41 44 42 46
rect 38 36 42 44
rect 38 34 39 36
rect 41 34 42 36
rect 38 32 42 34
rect 14 24 39 26
rect 14 22 15 24
rect 17 22 36 24
rect 38 22 39 24
rect 14 17 18 22
rect 14 15 15 17
rect 17 15 18 17
rect 14 13 18 15
rect 35 17 39 22
rect 35 15 36 17
rect 38 16 62 17
rect 38 15 58 16
rect 35 14 58 15
rect 60 14 62 16
rect 35 13 62 14
rect 40 6 56 7
rect 40 4 42 6
rect 44 4 52 6
rect 54 4 56 6
rect 40 3 56 4
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< labels >>
rlabel alu1 8 40 8 40 6 a
rlabel alu1 16 32 16 32 6 a
rlabel alu1 24 40 24 40 6 a
rlabel alu1 16 60 16 60 6 z
rlabel alu1 24 56 24 56 6 z
rlabel alu1 40 56 40 56 6 z
rlabel ndifct1 48 24 48 24 6 z
rlabel alu1 56 48 56 48 6 b
rlabel alu1 48 44 48 44 6 z
rlabel via1 32 4 32 4 6 vss
rlabel via1 32 84 32 84 6 vdd
<< end >>
