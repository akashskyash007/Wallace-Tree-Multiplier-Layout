magic
tech scmos
timestamp 1199202044
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 60 41 65
rect 49 60 51 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 9 37 31 39
rect 14 35 27 37
rect 29 35 31 37
rect 14 33 31 35
rect 37 37 51 39
rect 37 35 43 37
rect 45 35 47 37
rect 37 33 47 35
rect 14 30 16 33
rect 24 30 26 33
rect 37 30 39 33
rect 14 6 16 10
rect 24 6 26 10
rect 37 7 39 12
<< ndif >>
rect 6 21 14 30
rect 6 19 9 21
rect 11 19 14 21
rect 6 14 14 19
rect 6 12 9 14
rect 11 12 14 14
rect 6 10 14 12
rect 16 28 24 30
rect 16 26 19 28
rect 21 26 24 28
rect 16 21 24 26
rect 16 19 19 21
rect 21 19 24 21
rect 16 10 24 19
rect 26 21 37 30
rect 26 19 31 21
rect 33 19 37 21
rect 26 14 37 19
rect 26 12 31 14
rect 33 12 37 14
rect 39 28 46 30
rect 39 26 42 28
rect 44 26 46 28
rect 39 21 46 26
rect 39 19 42 21
rect 44 19 46 21
rect 39 17 46 19
rect 39 12 44 17
rect 26 10 35 12
<< pdif >>
rect 4 55 9 69
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 66 19 69
rect 11 64 14 66
rect 16 64 19 66
rect 11 58 19 64
rect 11 56 14 58
rect 16 56 19 58
rect 11 42 19 56
rect 21 53 29 69
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 60 37 69
rect 31 58 39 60
rect 31 56 34 58
rect 36 56 39 58
rect 31 42 39 56
rect 41 53 49 60
rect 41 51 44 53
rect 46 51 49 53
rect 41 46 49 51
rect 41 44 44 46
rect 46 44 49 46
rect 41 42 49 44
rect 51 58 58 60
rect 51 56 54 58
rect 56 56 58 58
rect 51 50 58 56
rect 51 48 54 50
rect 56 48 58 50
rect 51 42 58 48
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 23 53 27 55
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 2 44 4 46
rect 6 44 24 46
rect 26 44 27 46
rect 2 42 27 44
rect 2 41 14 42
rect 9 30 14 41
rect 41 37 55 38
rect 41 35 43 37
rect 45 35 55 37
rect 41 34 55 35
rect 9 28 23 30
rect 9 26 19 28
rect 21 26 23 28
rect 49 26 55 34
rect 18 21 23 26
rect 18 19 19 21
rect 21 19 23 21
rect 18 17 23 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 14 10 16 30
rect 24 10 26 30
rect 37 12 39 30
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 60
rect 49 42 51 60
<< polyct0 >>
rect 27 35 29 37
<< polyct1 >>
rect 43 35 45 37
<< ndifct0 >>
rect 9 19 11 21
rect 9 12 11 14
rect 31 19 33 21
rect 31 12 33 14
rect 42 26 44 28
rect 42 19 44 21
<< ndifct1 >>
rect 19 26 21 28
rect 19 19 21 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 14 64 16 66
rect 14 56 16 58
rect 34 56 36 58
rect 44 51 46 53
rect 44 44 46 46
rect 54 56 56 58
rect 54 48 56 50
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 51 26 53
rect 24 44 26 46
<< alu0 >>
rect 13 66 17 68
rect 13 64 14 66
rect 16 64 17 66
rect 13 58 17 64
rect 13 56 14 58
rect 16 56 17 58
rect 13 54 17 56
rect 33 58 37 68
rect 33 56 34 58
rect 36 56 37 58
rect 33 54 37 56
rect 53 58 57 68
rect 53 56 54 58
rect 56 56 57 58
rect 43 53 47 55
rect 43 51 44 53
rect 46 51 47 53
rect 43 46 47 51
rect 53 50 57 56
rect 53 48 54 50
rect 56 48 57 50
rect 53 46 57 48
rect 33 44 44 46
rect 46 44 47 46
rect 33 42 47 44
rect 33 38 37 42
rect 25 37 37 38
rect 25 35 27 37
rect 29 35 37 37
rect 25 34 37 35
rect 33 30 37 34
rect 33 28 45 30
rect 33 26 42 28
rect 44 26 45 28
rect 7 21 13 22
rect 7 19 9 21
rect 11 19 13 21
rect 7 14 13 19
rect 29 21 35 22
rect 29 19 31 21
rect 33 19 35 21
rect 7 12 9 14
rect 11 12 13 14
rect 29 14 35 19
rect 41 21 45 26
rect 41 19 42 21
rect 44 19 45 21
rect 41 17 45 19
rect 29 12 31 14
rect 33 12 35 14
<< labels >>
rlabel alu0 43 23 43 23 6 an
rlabel alu0 31 36 31 36 6 an
rlabel alu0 45 48 45 48 6 an
rlabel alu1 12 36 12 36 6 z
rlabel alu1 4 48 4 48 6 z
rlabel alu1 20 24 20 24 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel polyct1 44 36 44 36 6 a
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 32 52 32 6 a
<< end >>
