magic
tech scmos
timestamp 1199202686
<< ab >>
rect 0 0 96 72
<< nwell >>
rect -5 32 101 77
<< pwell >>
rect -5 -5 101 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 70 53 72 58
rect 80 53 82 58
rect 9 35 11 40
rect 19 35 21 40
rect 29 35 31 40
rect 39 35 41 40
rect 49 35 51 40
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 31 35
rect 19 31 27 33
rect 29 31 31 33
rect 19 29 31 31
rect 35 33 51 35
rect 59 35 61 40
rect 70 35 72 40
rect 80 35 82 40
rect 59 33 72 35
rect 76 33 82 35
rect 35 31 37 33
rect 39 31 41 33
rect 35 29 41 31
rect 59 31 61 33
rect 63 31 65 33
rect 59 29 65 31
rect 76 31 78 33
rect 80 31 82 33
rect 76 29 82 31
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 12 2 14 7
rect 19 2 21 7
rect 29 2 31 7
rect 36 2 38 7
<< ndif >>
rect 3 7 12 26
rect 14 7 19 26
rect 21 17 29 26
rect 21 15 24 17
rect 26 15 29 17
rect 21 7 29 15
rect 31 7 36 26
rect 38 7 47 26
rect 3 5 6 7
rect 8 5 10 7
rect 3 3 10 5
rect 40 5 42 7
rect 44 5 47 7
rect 40 3 47 5
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 40 9 55
rect 11 56 19 66
rect 11 54 14 56
rect 16 54 19 56
rect 11 49 19 54
rect 11 47 14 49
rect 16 47 19 49
rect 11 40 19 47
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 40 29 55
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 49 39 55
rect 31 47 34 49
rect 36 47 39 49
rect 31 40 39 47
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 40 49 55
rect 51 57 59 66
rect 51 55 54 57
rect 56 55 59 57
rect 51 49 59 55
rect 51 47 54 49
rect 56 47 59 49
rect 51 40 59 47
rect 61 64 68 66
rect 61 62 64 64
rect 66 62 68 64
rect 61 57 68 62
rect 61 55 64 57
rect 66 55 68 57
rect 61 53 68 55
rect 61 40 70 53
rect 72 51 80 53
rect 72 49 75 51
rect 77 49 80 51
rect 72 44 80 49
rect 72 42 75 44
rect 77 42 80 44
rect 72 40 80 42
rect 82 51 90 53
rect 82 49 85 51
rect 87 49 90 51
rect 82 40 90 49
<< alu1 >>
rect -2 67 98 72
rect -2 65 77 67
rect 79 65 85 67
rect 87 65 98 67
rect -2 64 98 65
rect 33 57 38 59
rect 33 55 34 57
rect 36 55 38 57
rect 33 50 38 55
rect 74 51 78 53
rect 74 50 75 51
rect 2 49 75 50
rect 77 49 78 51
rect 2 47 14 49
rect 16 47 34 49
rect 36 47 54 49
rect 56 47 78 49
rect 2 46 78 47
rect 2 18 6 46
rect 74 44 78 46
rect 74 42 75 44
rect 77 42 78 44
rect 25 38 49 42
rect 74 40 78 42
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 25 33 31 38
rect 45 34 49 38
rect 25 31 27 33
rect 29 31 31 33
rect 25 30 31 31
rect 45 33 65 34
rect 45 31 61 33
rect 63 31 65 33
rect 45 30 65 31
rect 73 33 87 34
rect 73 31 78 33
rect 80 31 87 33
rect 73 30 87 31
rect 73 26 79 30
rect 10 22 79 26
rect 2 17 31 18
rect 2 15 24 17
rect 26 15 31 17
rect 2 14 31 15
rect -2 7 98 8
rect -2 5 6 7
rect 8 5 42 7
rect 44 5 77 7
rect 79 5 85 7
rect 87 5 98 7
rect -2 0 98 5
<< ptie >>
rect 75 7 89 24
rect 75 5 77 7
rect 79 5 85 7
rect 87 5 89 7
rect 75 3 89 5
<< ntie >>
rect 75 67 89 69
rect 75 65 77 67
rect 79 65 85 67
rect 87 65 89 67
rect 75 61 89 65
<< nmos >>
rect 12 7 14 26
rect 19 7 21 26
rect 29 7 31 26
rect 36 7 38 26
<< pmos >>
rect 9 40 11 66
rect 19 40 21 66
rect 29 40 31 66
rect 39 40 41 66
rect 49 40 51 66
rect 59 40 61 66
rect 70 40 72 53
rect 80 40 82 53
<< polyct0 >>
rect 37 31 39 33
<< polyct1 >>
rect 11 31 13 33
rect 27 31 29 33
rect 61 31 63 33
rect 78 31 80 33
<< ndifct1 >>
rect 24 15 26 17
rect 6 5 8 7
rect 42 5 44 7
<< ntiect1 >>
rect 77 65 79 67
rect 85 65 87 67
<< ptiect1 >>
rect 77 5 79 7
rect 85 5 87 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 54 16 56
rect 24 62 26 64
rect 24 55 26 57
rect 44 62 46 64
rect 44 55 46 57
rect 54 55 56 57
rect 64 62 66 64
rect 64 55 66 57
rect 85 49 87 51
<< pdifct1 >>
rect 14 47 16 49
rect 34 55 36 57
rect 34 47 36 49
rect 54 47 56 49
rect 75 49 77 51
rect 75 42 77 44
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 56 17 58
rect 13 54 14 56
rect 16 54 17 56
rect 22 57 28 62
rect 42 62 44 64
rect 46 62 48 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 13 50 17 54
rect 42 57 48 62
rect 62 62 64 64
rect 66 62 68 64
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 53 57 57 59
rect 53 55 54 57
rect 56 55 57 57
rect 53 50 57 55
rect 62 57 68 62
rect 62 55 64 57
rect 66 55 68 57
rect 62 54 68 55
rect 84 51 88 64
rect 84 49 85 51
rect 87 49 88 51
rect 84 47 88 49
rect 35 33 41 34
rect 35 31 37 33
rect 39 31 41 33
rect 35 26 41 31
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 24 20 24 6 a
rlabel alu1 28 24 28 24 6 a
rlabel polyct1 28 32 28 32 6 b
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 48 4 48 4 6 vss
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 52 24 52 24 6 a
rlabel alu1 52 32 52 32 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 48 68 48 68 6 vdd
rlabel alu1 60 24 60 24 6 a
rlabel alu1 68 24 68 24 6 a
rlabel alu1 76 28 76 28 6 a
rlabel alu1 60 32 60 32 6 b
rlabel alu1 60 48 60 48 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 76 48 76 48 6 z
rlabel alu1 84 32 84 32 6 a
<< end >>
