magic
tech scmos
timestamp 1199202230
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 61 15 63
rect 9 59 11 61
rect 13 59 15 61
rect 9 57 15 59
rect 9 54 11 57
rect 9 30 11 42
rect 9 19 11 24
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 11 28 18 30
rect 11 26 14 28
rect 16 26 18 28
rect 11 24 18 26
<< pdif >>
rect 2 71 8 73
rect 2 69 4 71
rect 6 69 8 71
rect 2 65 8 69
rect 2 54 7 65
rect 2 42 9 54
rect 11 48 16 54
rect 11 46 18 48
rect 11 44 14 46
rect 16 44 18 46
rect 11 42 18 44
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 71 26 79
rect -2 69 4 71
rect 6 69 26 71
rect -2 68 26 69
rect 2 61 14 63
rect 2 59 11 61
rect 13 59 14 61
rect 2 57 14 59
rect 2 49 6 57
rect 10 46 18 47
rect 10 44 14 46
rect 16 44 18 46
rect 10 43 18 44
rect 10 39 14 43
rect 2 33 14 39
rect 2 28 8 33
rect 2 26 4 28
rect 6 26 8 28
rect 2 25 8 26
rect -2 1 26 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 24 11 30
<< pmos >>
rect 9 42 11 54
<< polyct1 >>
rect 11 59 13 61
<< ndifct0 >>
rect 14 26 16 28
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct1 >>
rect 4 69 6 71
rect 14 44 16 46
<< alu0 >>
rect 12 28 18 29
rect 12 26 14 28
rect 16 26 18 28
rect 12 12 18 26
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 4 56 4 56 6 a
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 40 12 40 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel polyct1 12 60 12 60 6 a
<< end >>
