magic
tech scmos
timestamp 1199202215
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 64 11 70
rect 20 67 26 69
rect 20 65 22 67
rect 24 65 26 67
rect 20 63 26 65
rect 9 43 11 46
rect 9 41 18 43
rect 12 39 14 41
rect 16 39 18 41
rect 12 26 18 39
rect 22 36 26 63
rect 36 57 38 62
rect 43 57 45 62
rect 36 46 38 49
rect 43 46 45 49
rect 32 44 38 46
rect 32 42 34 44
rect 36 42 38 44
rect 32 40 38 42
rect 42 44 48 46
rect 42 42 44 44
rect 46 42 48 44
rect 42 40 48 42
rect 22 34 37 36
rect 9 24 18 26
rect 23 28 29 30
rect 23 26 25 28
rect 27 26 29 28
rect 23 24 29 26
rect 33 28 37 34
rect 33 24 49 28
rect 9 21 11 24
rect 16 21 18 24
rect 26 21 28 24
rect 33 21 35 24
rect 40 21 42 24
rect 47 21 49 24
rect 26 10 28 15
rect 33 10 35 15
rect 40 10 42 15
rect 47 11 49 15
rect 9 2 11 6
rect 16 2 18 6
<< ndif >>
rect 2 19 9 21
rect 2 17 4 19
rect 6 17 9 19
rect 2 6 9 17
rect 11 6 16 21
rect 18 19 26 21
rect 18 17 21 19
rect 23 17 26 19
rect 18 15 26 17
rect 28 15 33 21
rect 35 15 40 21
rect 42 15 47 21
rect 49 19 56 21
rect 49 17 52 19
rect 54 17 56 19
rect 49 15 56 17
rect 18 6 24 15
<< pdif >>
rect 2 58 9 64
rect 2 56 4 58
rect 6 56 9 58
rect 2 50 9 56
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 11 62 18 64
rect 11 60 14 62
rect 16 60 18 62
rect 11 46 18 60
rect 28 67 34 69
rect 28 65 30 67
rect 32 65 34 67
rect 28 57 34 65
rect 28 49 36 57
rect 38 49 43 57
rect 45 53 56 57
rect 45 51 52 53
rect 54 51 56 53
rect 45 49 56 51
<< alu1 >>
rect -2 67 66 72
rect -2 65 22 67
rect 24 65 30 67
rect 32 65 53 67
rect 55 65 66 67
rect -2 64 66 65
rect 12 62 18 64
rect 12 60 14 62
rect 16 60 18 62
rect 2 58 8 59
rect 2 56 4 58
rect 6 56 8 58
rect 12 56 18 60
rect 2 52 8 56
rect 22 53 56 59
rect 2 50 18 52
rect 2 48 4 50
rect 6 48 18 50
rect 2 46 18 48
rect 2 34 8 46
rect 22 42 28 53
rect 50 51 52 53
rect 54 51 56 53
rect 12 41 28 42
rect 12 39 14 41
rect 16 39 28 41
rect 12 38 28 39
rect 33 44 39 46
rect 33 42 34 44
rect 36 42 39 44
rect 33 34 39 42
rect 2 28 19 34
rect 23 30 39 34
rect 23 28 29 30
rect 2 19 8 28
rect 23 26 25 28
rect 27 26 29 28
rect 23 24 29 26
rect 2 17 4 19
rect 6 17 8 19
rect 2 13 8 17
rect 19 19 25 20
rect 19 17 21 19
rect 23 17 25 19
rect 19 8 25 17
rect 50 19 56 51
rect 50 17 52 19
rect 54 17 56 19
rect 50 13 56 17
rect -2 7 66 8
rect -2 5 53 7
rect 55 5 66 7
rect -2 0 66 5
<< ptie >>
rect 51 7 57 9
rect 51 5 53 7
rect 55 5 57 7
rect 51 3 57 5
<< ntie >>
rect 51 67 57 69
rect 51 65 53 67
rect 55 65 57 67
rect 51 63 57 65
<< nmos >>
rect 9 6 11 21
rect 16 6 18 21
rect 26 15 28 21
rect 33 15 35 21
rect 40 15 42 21
rect 47 15 49 21
<< pmos >>
rect 9 46 11 64
rect 36 49 38 57
rect 43 49 45 57
<< polyct0 >>
rect 44 42 46 44
<< polyct1 >>
rect 22 65 24 67
rect 14 39 16 41
rect 34 42 36 44
rect 25 26 27 28
<< ndifct1 >>
rect 4 17 6 19
rect 21 17 23 19
rect 52 17 54 19
<< ntiect1 >>
rect 53 65 55 67
<< ptiect1 >>
rect 53 5 55 7
<< pdifct1 >>
rect 4 56 6 58
rect 4 48 6 50
rect 14 60 16 62
rect 30 65 32 67
rect 52 51 54 53
<< alu0 >>
rect 43 44 47 49
rect 43 42 44 44
rect 46 42 47 44
rect 43 8 47 42
<< labels >>
rlabel polyct1 15 40 15 40 6 an
rlabel ndifct1 53 18 53 18 6 an
rlabel pdifct1 53 52 53 52 6 an
rlabel alu1 12 32 12 32 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 32 28 32 6 a
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 36 36 36 6 a
rlabel alu1 32 68 32 68 6 vdd
<< end >>
