magic
tech scmos
timestamp 1199203438
<< ab >>
rect 0 0 176 72
<< nwell >>
rect -5 32 181 77
<< pwell >>
rect -5 -5 181 32
<< poly >>
rect 22 66 24 70
rect 32 66 34 70
rect 42 66 44 70
rect 52 66 54 70
rect 62 66 64 70
rect 72 66 74 70
rect 82 66 84 70
rect 92 66 94 70
rect 102 66 104 70
rect 112 66 114 70
rect 122 66 124 70
rect 132 66 134 70
rect 142 66 144 70
rect 152 66 154 70
rect 162 66 164 70
rect 22 31 24 38
rect 32 35 34 38
rect 42 35 44 38
rect 32 33 44 35
rect 52 35 54 38
rect 62 35 64 38
rect 72 35 74 38
rect 82 35 84 38
rect 92 35 94 38
rect 102 35 104 38
rect 112 35 114 38
rect 122 35 124 38
rect 132 35 134 38
rect 52 33 58 35
rect 62 33 74 35
rect 32 31 35 33
rect 37 31 40 33
rect 9 29 40 31
rect 56 29 58 33
rect 68 31 70 33
rect 72 31 74 33
rect 68 29 74 31
rect 78 33 94 35
rect 98 33 104 35
rect 110 33 116 35
rect 78 31 80 33
rect 82 31 90 33
rect 78 29 90 31
rect 98 29 100 33
rect 110 31 112 33
rect 114 31 116 33
rect 110 29 116 31
rect 9 26 11 29
rect 19 26 21 29
rect 38 26 40 29
rect 49 25 51 29
rect 56 27 64 29
rect 58 25 60 27
rect 62 25 64 27
rect 71 26 73 29
rect 78 26 80 29
rect 58 23 64 25
rect 9 2 11 6
rect 19 2 21 6
rect 38 4 40 7
rect 49 4 51 7
rect 88 20 90 29
rect 94 27 100 29
rect 94 25 96 27
rect 98 25 100 27
rect 114 26 116 29
rect 121 33 134 35
rect 121 31 127 33
rect 129 31 134 33
rect 142 35 144 38
rect 152 35 154 38
rect 142 33 154 35
rect 162 33 164 38
rect 142 31 145 33
rect 147 31 150 33
rect 121 29 134 31
rect 138 29 150 31
rect 161 31 167 33
rect 161 29 163 31
rect 165 29 167 31
rect 121 26 123 29
rect 131 26 133 29
rect 138 26 140 29
rect 94 23 100 25
rect 95 20 97 23
rect 148 24 150 29
rect 155 27 167 29
rect 155 24 157 27
rect 38 2 51 4
rect 71 2 73 6
rect 78 2 80 6
rect 88 2 90 6
rect 95 2 97 6
rect 114 2 116 6
rect 121 2 123 6
rect 131 2 133 6
rect 138 2 140 6
rect 148 2 150 6
rect 155 2 157 6
<< ndif >>
rect 4 18 9 26
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 4 6 9 12
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 6 19 22
rect 21 24 28 26
rect 21 22 24 24
rect 26 22 28 24
rect 21 20 28 22
rect 21 6 26 20
rect 32 16 38 26
rect 30 9 38 16
rect 30 7 32 9
rect 34 7 38 9
rect 40 25 47 26
rect 40 24 49 25
rect 40 22 43 24
rect 45 22 49 24
rect 40 7 49 22
rect 51 20 56 25
rect 66 20 71 26
rect 51 17 71 20
rect 51 15 60 17
rect 62 15 71 17
rect 51 10 71 15
rect 51 8 60 10
rect 62 8 71 10
rect 51 7 71 8
rect 30 5 36 7
rect 53 6 71 7
rect 73 6 78 26
rect 80 20 85 26
rect 102 20 114 26
rect 80 17 88 20
rect 80 15 83 17
rect 85 15 88 17
rect 80 6 88 15
rect 90 6 95 20
rect 97 10 114 20
rect 97 8 100 10
rect 102 8 109 10
rect 111 8 114 10
rect 97 6 114 8
rect 116 6 121 26
rect 123 17 131 26
rect 123 15 126 17
rect 128 15 131 17
rect 123 6 131 15
rect 133 6 138 26
rect 140 24 145 26
rect 140 10 148 24
rect 140 8 143 10
rect 145 8 148 10
rect 140 6 148 8
rect 150 6 155 24
rect 157 19 162 24
rect 157 17 164 19
rect 157 15 160 17
rect 162 15 164 17
rect 157 13 164 15
rect 157 6 162 13
<< pdif >>
rect 14 64 22 66
rect 14 62 17 64
rect 19 62 22 64
rect 14 38 22 62
rect 24 42 32 66
rect 24 40 27 42
rect 29 40 32 42
rect 24 38 32 40
rect 34 64 42 66
rect 34 62 37 64
rect 39 62 42 64
rect 34 38 42 62
rect 44 42 52 66
rect 44 40 47 42
rect 49 40 52 42
rect 44 38 52 40
rect 54 49 62 66
rect 54 47 57 49
rect 59 47 62 49
rect 54 38 62 47
rect 64 57 72 66
rect 64 55 67 57
rect 69 55 72 57
rect 64 38 72 55
rect 74 49 82 66
rect 74 47 77 49
rect 79 47 82 49
rect 74 38 82 47
rect 84 42 92 66
rect 84 40 87 42
rect 89 40 92 42
rect 84 38 92 40
rect 94 49 102 66
rect 94 47 97 49
rect 99 47 102 49
rect 94 42 102 47
rect 94 40 97 42
rect 99 40 102 42
rect 94 38 102 40
rect 104 57 112 66
rect 104 55 107 57
rect 109 55 112 57
rect 104 50 112 55
rect 104 48 107 50
rect 109 48 112 50
rect 104 38 112 48
rect 114 64 122 66
rect 114 62 117 64
rect 119 62 122 64
rect 114 57 122 62
rect 114 55 117 57
rect 119 55 122 57
rect 114 38 122 55
rect 124 56 132 66
rect 124 54 127 56
rect 129 54 132 56
rect 124 49 132 54
rect 124 47 127 49
rect 129 47 132 49
rect 124 38 132 47
rect 134 64 142 66
rect 134 62 137 64
rect 139 62 142 64
rect 134 57 142 62
rect 134 55 137 57
rect 139 55 142 57
rect 134 38 142 55
rect 144 56 152 66
rect 144 54 147 56
rect 149 54 152 56
rect 144 49 152 54
rect 144 47 147 49
rect 149 47 152 49
rect 144 38 152 47
rect 154 64 162 66
rect 154 62 157 64
rect 159 62 162 64
rect 154 57 162 62
rect 154 55 157 57
rect 159 55 162 57
rect 154 38 162 55
rect 164 58 169 66
rect 164 56 171 58
rect 164 54 167 56
rect 169 54 171 56
rect 164 49 171 54
rect 164 47 167 49
rect 169 47 171 49
rect 164 45 171 47
rect 164 38 169 45
<< alu1 >>
rect -2 67 178 72
rect -2 65 5 67
rect 7 65 178 67
rect -2 64 178 65
rect 10 49 101 50
rect 10 47 57 49
rect 59 47 77 49
rect 79 47 97 49
rect 99 47 101 49
rect 10 46 101 47
rect 10 25 14 46
rect 26 33 38 35
rect 26 31 35 33
rect 37 31 38 33
rect 26 29 38 31
rect 10 24 18 25
rect 10 22 14 24
rect 16 22 18 24
rect 10 21 18 22
rect 34 21 38 29
rect 96 42 101 46
rect 96 40 97 42
rect 99 40 107 42
rect 96 38 107 40
rect 103 18 107 38
rect 113 33 119 42
rect 129 38 166 42
rect 129 34 135 38
rect 114 31 119 33
rect 113 26 119 31
rect 125 33 135 34
rect 125 31 127 33
rect 129 31 135 33
rect 125 30 135 31
rect 139 33 151 34
rect 139 31 145 33
rect 147 31 151 33
rect 139 30 151 31
rect 162 31 166 38
rect 139 26 143 30
rect 113 22 143 26
rect 162 29 163 31
rect 165 29 166 31
rect 162 21 166 29
rect 81 17 111 18
rect 81 15 83 17
rect 85 15 111 17
rect 81 14 111 15
rect -2 7 32 8
rect 34 7 178 8
rect -2 5 169 7
rect 171 5 178 7
rect -2 0 178 5
<< ptie >>
rect 167 7 173 9
rect 167 5 169 7
rect 171 5 173 7
rect 167 3 173 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 40 9 65
<< nmos >>
rect 9 6 11 26
rect 19 6 21 26
rect 38 7 40 26
rect 49 7 51 25
rect 71 6 73 26
rect 78 6 80 26
rect 88 6 90 20
rect 95 6 97 20
rect 114 6 116 26
rect 121 6 123 26
rect 131 6 133 26
rect 138 6 140 26
rect 148 6 150 24
rect 155 6 157 24
<< pmos >>
rect 22 38 24 66
rect 32 38 34 66
rect 42 38 44 66
rect 52 38 54 66
rect 62 38 64 66
rect 72 38 74 66
rect 82 38 84 66
rect 92 38 94 66
rect 102 38 104 66
rect 112 38 114 66
rect 122 38 124 66
rect 132 38 134 66
rect 142 38 144 66
rect 152 38 154 66
rect 162 38 164 66
<< polyct0 >>
rect 70 31 72 33
rect 80 31 82 33
rect 112 31 113 33
rect 60 25 62 27
rect 96 25 98 27
<< polyct1 >>
rect 35 31 37 33
rect 113 31 114 33
rect 127 31 129 33
rect 145 31 147 33
rect 163 29 165 31
<< ndifct0 >>
rect 4 14 6 16
rect 24 22 26 24
rect 32 8 34 9
rect 43 22 45 24
rect 60 15 62 17
rect 60 8 62 10
rect 100 8 102 10
rect 109 8 111 10
rect 126 15 128 17
rect 143 8 145 10
rect 160 15 162 17
<< ndifct1 >>
rect 14 22 16 24
rect 32 7 34 8
rect 83 15 85 17
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 169 5 171 7
<< pdifct0 >>
rect 17 62 19 64
rect 27 40 29 42
rect 37 62 39 64
rect 47 40 49 42
rect 67 55 69 57
rect 87 40 89 42
rect 107 55 109 57
rect 107 48 109 50
rect 117 62 119 64
rect 117 55 119 57
rect 127 54 129 56
rect 127 47 129 49
rect 137 62 139 64
rect 137 55 139 57
rect 147 54 149 56
rect 147 47 149 49
rect 157 62 159 64
rect 157 55 159 57
rect 167 54 169 56
rect 167 47 169 49
<< pdifct1 >>
rect 57 47 59 49
rect 77 47 79 49
rect 97 47 99 49
rect 97 40 99 42
<< alu0 >>
rect 15 62 17 64
rect 19 62 21 64
rect 15 61 21 62
rect 35 62 37 64
rect 39 62 41 64
rect 35 61 41 62
rect 115 62 117 64
rect 119 62 121 64
rect 2 57 111 58
rect 2 55 67 57
rect 69 55 107 57
rect 109 55 111 57
rect 2 54 111 55
rect 115 57 121 62
rect 135 62 137 64
rect 139 62 141 64
rect 115 55 117 57
rect 119 55 121 57
rect 115 54 121 55
rect 126 56 130 58
rect 126 54 127 56
rect 129 54 130 56
rect 135 57 141 62
rect 155 62 157 64
rect 159 62 161 64
rect 135 55 137 57
rect 139 55 141 57
rect 135 54 141 55
rect 146 56 150 58
rect 146 54 147 56
rect 149 54 150 56
rect 155 57 161 62
rect 155 55 157 57
rect 159 55 161 57
rect 155 54 161 55
rect 166 56 170 58
rect 166 54 167 56
rect 169 54 170 56
rect 2 17 6 54
rect 106 50 111 54
rect 126 50 130 54
rect 146 50 150 54
rect 166 50 170 54
rect 106 48 107 50
rect 109 49 174 50
rect 109 48 127 49
rect 106 47 127 48
rect 129 47 147 49
rect 149 47 167 49
rect 169 47 174 49
rect 106 46 174 47
rect 25 42 92 43
rect 25 40 27 42
rect 29 40 47 42
rect 49 40 87 42
rect 89 40 92 42
rect 25 39 92 40
rect 23 24 27 26
rect 23 22 24 24
rect 26 22 27 24
rect 23 17 27 22
rect 42 24 46 39
rect 68 33 74 39
rect 68 31 70 33
rect 72 31 74 33
rect 68 30 74 31
rect 78 33 84 34
rect 78 31 80 33
rect 82 31 84 33
rect 59 27 63 29
rect 59 26 60 27
rect 42 22 43 24
rect 45 22 46 24
rect 42 20 46 22
rect 49 25 60 26
rect 62 26 63 27
rect 78 26 84 31
rect 62 25 84 26
rect 49 22 84 25
rect 88 29 92 39
rect 88 27 99 29
rect 88 25 96 27
rect 98 25 99 27
rect 88 23 99 25
rect 49 17 53 22
rect 111 33 113 35
rect 111 31 112 33
rect 111 29 113 31
rect 170 18 174 46
rect 2 16 53 17
rect 2 14 4 16
rect 6 14 53 16
rect 2 13 53 14
rect 58 17 64 18
rect 58 15 60 17
rect 62 15 64 17
rect 58 10 64 15
rect 124 17 174 18
rect 124 15 126 17
rect 128 15 160 17
rect 162 15 174 17
rect 124 14 174 15
rect 30 9 36 10
rect 30 8 32 9
rect 34 8 36 9
rect 58 8 60 10
rect 62 8 64 10
rect 97 10 113 11
rect 97 8 100 10
rect 102 8 109 10
rect 111 8 113 10
rect 141 10 147 11
rect 141 8 143 10
rect 145 8 147 10
<< labels >>
rlabel alu0 25 19 25 19 6 an
rlabel alu0 27 15 27 15 6 an
rlabel alu0 66 24 66 24 6 an
rlabel alu0 81 28 81 28 6 an
rlabel alu0 71 36 71 36 6 bn
rlabel alu0 44 31 44 31 6 bn
rlabel alu0 93 26 93 26 6 bn
rlabel alu0 58 41 58 41 6 bn
rlabel alu0 108 52 108 52 6 an
rlabel alu0 128 52 128 52 6 an
rlabel alu0 56 56 56 56 6 an
rlabel alu0 149 16 149 16 6 an
rlabel alu0 140 48 140 48 6 an
rlabel alu0 148 52 148 52 6 an
rlabel alu0 168 52 168 52 6 an
rlabel alu1 12 32 12 32 6 z
rlabel alu1 28 32 28 32 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 28 36 28 6 b
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 88 4 88 4 6 vss
rlabel alu1 100 16 100 16 6 z
rlabel ndifct1 84 16 84 16 6 z
rlabel alu1 92 16 92 16 6 z
rlabel alu1 100 40 100 40 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 76 48 76 48 6 z
rlabel alu1 84 48 84 48 6 z
rlabel alu1 92 48 92 48 6 z
rlabel alu1 88 68 88 68 6 vdd
rlabel alu1 108 16 108 16 6 z
rlabel alu1 124 24 124 24 6 a1
rlabel alu1 132 24 132 24 6 a1
rlabel alu1 140 24 140 24 6 a1
rlabel alu1 116 32 116 32 6 a1
rlabel alu1 140 40 140 40 6 a2
rlabel alu1 132 36 132 36 6 a2
rlabel alu1 148 32 148 32 6 a1
rlabel alu1 164 28 164 28 6 a2
rlabel alu1 148 40 148 40 6 a2
rlabel alu1 156 40 156 40 6 a2
<< end >>
