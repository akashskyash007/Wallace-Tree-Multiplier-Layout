magic
tech scmos
timestamp 1199202282
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 61 11 65
rect 9 39 11 43
rect 9 37 16 39
rect 9 35 12 37
rect 14 35 16 37
rect 9 33 16 35
rect 9 30 11 33
rect 9 14 11 18
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 18 9 24
rect 11 22 19 30
rect 11 20 14 22
rect 16 20 19 22
rect 11 18 19 20
<< pdif >>
rect 13 61 20 63
rect 4 56 9 61
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 59 15 61
rect 17 59 20 61
rect 11 43 20 59
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 68 26 79
rect 2 54 14 55
rect 2 52 4 54
rect 6 52 14 54
rect 2 49 14 52
rect 2 47 6 49
rect 2 45 4 47
rect 2 28 6 45
rect 18 39 22 55
rect 10 37 22 39
rect 10 35 12 37
rect 14 35 22 37
rect 10 33 22 35
rect 2 26 4 28
rect 2 17 6 26
rect -2 1 26 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 18 11 30
<< pmos >>
rect 9 43 11 61
<< polyct1 >>
rect 12 35 14 37
<< ndifct0 >>
rect 14 20 16 22
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct0 >>
rect 15 59 17 61
<< pdifct1 >>
rect 4 52 6 54
rect 4 45 6 47
<< alu0 >>
rect 13 61 19 68
rect 13 59 15 61
rect 17 59 19 61
rect 13 58 19 59
rect 6 43 7 49
rect 6 24 7 30
rect 13 22 17 24
rect 13 20 14 22
rect 16 20 17 22
rect 13 12 17 20
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 36 12 36 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 44 20 44 6 a
<< end >>
