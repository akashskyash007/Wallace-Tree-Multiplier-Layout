magic
tech scmos
timestamp 1199542123
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 13 94 15 98
rect 25 94 27 98
rect 37 94 39 98
rect 49 94 51 98
rect 13 33 15 55
rect 25 33 27 55
rect 37 33 39 55
rect 49 33 51 55
rect 7 31 51 33
rect 7 29 9 31
rect 11 29 51 31
rect 7 27 51 29
rect 13 24 15 27
rect 25 24 27 27
rect 37 24 39 27
rect 49 24 51 27
rect 13 2 15 6
rect 25 2 27 6
rect 37 2 39 6
rect 49 2 51 6
<< ndif >>
rect 5 11 13 24
rect 5 9 7 11
rect 9 9 13 11
rect 5 6 13 9
rect 15 21 25 24
rect 15 19 19 21
rect 21 19 25 21
rect 15 6 25 19
rect 27 21 37 24
rect 27 19 31 21
rect 33 19 37 21
rect 27 11 37 19
rect 27 9 31 11
rect 33 9 37 11
rect 27 6 37 9
rect 39 21 49 24
rect 39 19 43 21
rect 45 19 49 21
rect 39 6 49 19
rect 51 21 59 24
rect 51 19 55 21
rect 57 19 59 21
rect 51 11 59 19
rect 51 9 55 11
rect 57 9 59 11
rect 51 6 59 9
<< pdif >>
rect 5 91 13 94
rect 5 89 7 91
rect 9 89 13 91
rect 5 55 13 89
rect 15 81 25 94
rect 15 79 19 81
rect 21 79 25 81
rect 15 71 25 79
rect 15 69 19 71
rect 21 69 25 71
rect 15 61 25 69
rect 15 59 19 61
rect 21 59 25 61
rect 15 55 25 59
rect 27 91 37 94
rect 27 89 31 91
rect 33 89 37 91
rect 27 81 37 89
rect 27 79 31 81
rect 33 79 37 81
rect 27 71 37 79
rect 27 69 31 71
rect 33 69 37 71
rect 27 61 37 69
rect 27 59 31 61
rect 33 59 37 61
rect 27 55 37 59
rect 39 81 49 94
rect 39 79 43 81
rect 45 79 49 81
rect 39 71 49 79
rect 39 69 43 71
rect 45 69 49 71
rect 39 61 49 69
rect 39 59 43 61
rect 45 59 49 61
rect 39 55 49 59
rect 51 91 59 94
rect 51 89 55 91
rect 57 89 59 91
rect 51 81 59 89
rect 51 79 55 81
rect 57 79 59 81
rect 51 77 59 79
rect 51 55 56 77
<< alu1 >>
rect -2 91 72 100
rect -2 89 7 91
rect 9 89 31 91
rect 33 89 55 91
rect 57 89 72 91
rect -2 88 72 89
rect 8 31 12 83
rect 8 29 9 31
rect 11 29 12 31
rect 8 17 12 29
rect 18 81 22 83
rect 18 79 19 81
rect 21 79 22 81
rect 18 71 22 79
rect 18 69 19 71
rect 21 69 22 71
rect 18 61 22 69
rect 18 59 19 61
rect 21 59 22 61
rect 18 42 22 59
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 71 34 79
rect 30 69 31 71
rect 33 69 34 71
rect 30 61 34 69
rect 30 59 31 61
rect 33 59 34 61
rect 30 57 34 59
rect 42 81 46 83
rect 42 79 43 81
rect 45 79 46 81
rect 42 71 46 79
rect 42 69 43 71
rect 45 69 46 71
rect 42 61 46 69
rect 54 81 58 88
rect 54 79 55 81
rect 57 79 58 81
rect 54 70 58 79
rect 62 70 66 71
rect 54 69 66 70
rect 54 67 63 69
rect 65 67 66 69
rect 54 66 66 67
rect 42 59 43 61
rect 45 59 46 61
rect 42 42 46 59
rect 62 59 66 66
rect 62 57 63 59
rect 65 57 66 59
rect 62 55 66 57
rect 18 38 46 42
rect 18 21 22 38
rect 18 19 19 21
rect 21 19 22 21
rect 18 17 22 19
rect 30 21 34 23
rect 30 19 31 21
rect 33 19 34 21
rect 30 12 34 19
rect 42 21 46 38
rect 42 19 43 21
rect 45 19 46 21
rect 42 17 46 19
rect 54 36 58 37
rect 54 35 67 36
rect 54 33 55 35
rect 57 33 63 35
rect 65 33 67 35
rect 54 32 67 33
rect 54 21 58 32
rect 54 19 55 21
rect 57 19 58 21
rect 54 12 58 19
rect -2 11 72 12
rect -2 9 7 11
rect 9 9 31 11
rect 33 9 55 11
rect 57 9 72 11
rect -2 0 72 9
<< ptie >>
rect 53 35 67 37
rect 53 33 55 35
rect 57 33 63 35
rect 65 33 67 35
rect 53 31 67 33
<< ntie >>
rect 61 69 67 71
rect 61 67 63 69
rect 65 67 67 69
rect 61 59 67 67
rect 61 57 63 59
rect 65 57 67 59
rect 61 55 67 57
<< nmos >>
rect 13 6 15 24
rect 25 6 27 24
rect 37 6 39 24
rect 49 6 51 24
<< pmos >>
rect 13 55 15 94
rect 25 55 27 94
rect 37 55 39 94
rect 49 55 51 94
<< polyct1 >>
rect 9 29 11 31
<< ndifct1 >>
rect 7 9 9 11
rect 19 19 21 21
rect 31 19 33 21
rect 31 9 33 11
rect 43 19 45 21
rect 55 19 57 21
rect 55 9 57 11
<< ntiect1 >>
rect 63 67 65 69
rect 63 57 65 59
<< ptiect1 >>
rect 55 33 57 35
rect 63 33 65 35
<< pdifct1 >>
rect 7 89 9 91
rect 19 79 21 81
rect 19 69 21 71
rect 19 59 21 61
rect 31 89 33 91
rect 31 79 33 81
rect 31 69 33 71
rect 31 59 33 61
rect 43 79 45 81
rect 43 69 45 71
rect 43 59 45 61
rect 55 89 57 91
rect 55 79 57 81
<< labels >>
rlabel alu1 10 50 10 50 6 i
rlabel alu1 30 40 30 40 6 nq
rlabel alu1 20 50 20 50 6 nq
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 40 40 40 6 nq
rlabel alu1 35 94 35 94 6 vdd
<< end >>
