magic
tech scmos
timestamp 1199201751
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 20 66 22 71
rect 30 66 32 71
rect 42 66 44 71
rect 52 66 54 71
rect 9 60 11 65
rect 9 39 11 48
rect 20 39 22 56
rect 30 53 32 56
rect 30 51 38 53
rect 30 49 34 51
rect 36 49 38 51
rect 30 47 38 49
rect 42 47 44 56
rect 9 37 16 39
rect 9 35 12 37
rect 14 35 16 37
rect 9 33 16 35
rect 20 37 28 39
rect 20 35 24 37
rect 26 35 28 37
rect 20 33 28 35
rect 9 28 11 33
rect 25 30 27 33
rect 32 30 34 47
rect 42 45 48 47
rect 42 43 44 45
rect 46 43 48 45
rect 39 41 48 43
rect 39 30 41 41
rect 52 39 54 56
rect 52 37 58 39
rect 52 35 54 37
rect 56 35 58 37
rect 46 33 58 35
rect 46 30 48 33
rect 9 17 11 22
rect 25 13 27 18
rect 32 13 34 18
rect 39 13 41 18
rect 46 13 48 18
<< ndif >>
rect 13 28 25 30
rect 2 26 9 28
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 11 22 25 28
rect 13 18 25 22
rect 27 18 32 30
rect 34 18 39 30
rect 41 18 46 30
rect 48 24 53 30
rect 48 22 55 24
rect 48 20 51 22
rect 53 20 55 22
rect 48 18 55 20
rect 13 11 23 18
rect 13 9 17 11
rect 19 9 23 11
rect 13 7 23 9
<< pdif >>
rect 34 71 40 73
rect 34 69 36 71
rect 38 69 40 71
rect 34 66 40 69
rect 13 62 20 66
rect 13 60 15 62
rect 17 60 20 62
rect 4 54 9 60
rect 2 52 9 54
rect 2 50 4 52
rect 6 50 9 52
rect 2 48 9 50
rect 11 56 20 60
rect 22 62 30 66
rect 22 60 25 62
rect 27 60 30 62
rect 22 56 30 60
rect 32 56 42 66
rect 44 62 52 66
rect 44 60 47 62
rect 49 60 52 62
rect 44 56 52 60
rect 54 64 61 66
rect 54 62 57 64
rect 59 62 61 64
rect 54 56 61 62
rect 11 48 18 56
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 36 71
rect 38 69 66 71
rect -2 68 66 69
rect 2 52 7 63
rect 2 50 4 52
rect 6 50 7 52
rect 2 48 7 50
rect 33 51 47 54
rect 2 26 6 48
rect 33 49 34 51
rect 36 50 47 51
rect 36 49 37 50
rect 33 46 37 49
rect 58 46 62 55
rect 25 42 37 46
rect 41 45 62 46
rect 41 43 44 45
rect 46 43 62 45
rect 41 42 62 43
rect 22 37 31 38
rect 22 35 24 37
rect 26 35 31 37
rect 22 34 31 35
rect 41 37 62 38
rect 41 35 54 37
rect 56 35 62 37
rect 41 34 62 35
rect 2 24 4 26
rect 2 23 6 24
rect 2 17 14 23
rect 26 30 31 34
rect 26 26 39 30
rect 58 17 62 34
rect -2 11 66 12
rect -2 9 17 11
rect 19 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 22 11 28
rect 25 18 27 30
rect 32 18 34 30
rect 39 18 41 30
rect 46 18 48 30
<< pmos >>
rect 9 48 11 60
rect 20 56 22 66
rect 30 56 32 66
rect 42 56 44 66
rect 52 56 54 66
<< polyct0 >>
rect 12 35 14 37
<< polyct1 >>
rect 34 49 36 51
rect 24 35 26 37
rect 44 43 46 45
rect 54 35 56 37
<< ndifct0 >>
rect 51 20 53 22
<< ndifct1 >>
rect 4 24 6 26
rect 17 9 19 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 15 60 17 62
rect 25 60 27 62
rect 47 60 49 62
rect 57 62 59 64
<< pdifct1 >>
rect 36 69 38 71
rect 4 50 6 52
<< alu0 >>
rect 14 62 18 68
rect 56 64 60 68
rect 14 60 15 62
rect 17 60 18 62
rect 14 58 18 60
rect 23 62 51 63
rect 23 60 25 62
rect 27 60 47 62
rect 49 60 51 62
rect 56 62 57 64
rect 59 62 60 64
rect 56 60 60 62
rect 23 59 51 60
rect 23 54 27 59
rect 14 50 27 54
rect 14 38 18 50
rect 10 37 18 38
rect 10 35 12 37
rect 14 35 18 37
rect 10 34 18 35
rect 14 31 18 34
rect 6 23 7 28
rect 14 27 22 31
rect 18 21 22 27
rect 50 22 54 24
rect 50 21 51 22
rect 18 20 51 21
rect 53 20 54 22
rect 18 17 54 20
<< labels >>
rlabel alu0 16 40 16 40 6 zn
rlabel alu0 36 19 36 19 6 zn
rlabel alu0 37 61 37 61 6 zn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 36 28 36 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 36 44 36 6 d
rlabel alu1 44 44 44 44 6 c
rlabel alu1 36 52 36 52 6 b
rlabel alu1 44 52 44 52 6 b
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 36 52 36 6 d
rlabel alu1 60 24 60 24 6 d
rlabel alu1 52 44 52 44 6 c
rlabel alu1 60 52 60 52 6 c
<< end >>
