magic
tech scmos
timestamp 1199202472
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 19 72 53 74
rect 9 64 11 69
rect 19 64 21 72
rect 29 64 31 68
rect 40 64 42 68
rect 51 60 53 72
rect 51 46 53 50
rect 50 44 56 46
rect 50 42 52 44
rect 54 42 56 44
rect 9 39 11 42
rect 2 37 12 39
rect 19 37 21 42
rect 29 39 31 42
rect 25 37 32 39
rect 2 35 4 37
rect 6 35 12 37
rect 2 33 12 35
rect 10 30 12 33
rect 25 35 28 37
rect 30 35 32 37
rect 25 33 32 35
rect 40 36 42 42
rect 50 40 56 42
rect 40 34 46 36
rect 25 31 27 33
rect 21 29 27 31
rect 40 32 42 34
rect 44 32 46 34
rect 40 30 46 32
rect 53 30 55 40
rect 21 25 23 29
rect 31 25 33 29
rect 41 27 43 30
rect 10 15 12 19
rect 21 9 23 14
rect 31 8 33 14
rect 41 12 43 16
rect 53 8 55 23
rect 31 6 55 8
<< ndif >>
rect 2 23 10 30
rect 2 21 4 23
rect 6 21 10 23
rect 2 19 10 21
rect 12 25 17 30
rect 48 27 53 30
rect 36 25 41 27
rect 12 22 21 25
rect 12 20 16 22
rect 18 20 21 22
rect 12 19 21 20
rect 14 18 21 19
rect 16 14 21 18
rect 23 23 31 25
rect 23 21 26 23
rect 28 21 31 23
rect 23 14 31 21
rect 33 23 41 25
rect 33 21 36 23
rect 38 21 41 23
rect 33 16 41 21
rect 43 23 53 27
rect 55 28 62 30
rect 55 26 58 28
rect 60 26 62 28
rect 55 23 62 26
rect 43 16 51 23
rect 33 14 38 16
rect 45 14 51 16
rect 45 12 47 14
rect 49 12 51 14
rect 45 10 51 12
<< pdif >>
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 42 9 60
rect 11 46 19 64
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 61 29 64
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 46 40 64
rect 31 44 35 46
rect 37 44 40 46
rect 31 42 40 44
rect 42 62 49 64
rect 42 60 45 62
rect 47 60 49 62
rect 42 50 51 60
rect 53 56 58 60
rect 53 54 60 56
rect 53 52 56 54
rect 58 52 60 54
rect 53 50 60 52
rect 42 42 48 50
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 10 55 14 63
rect 2 51 14 55
rect 20 61 31 62
rect 20 59 24 61
rect 26 59 31 61
rect 20 58 31 59
rect 2 37 7 51
rect 2 35 4 37
rect 6 35 7 37
rect 2 33 7 35
rect 20 39 24 58
rect 18 33 24 39
rect 20 30 24 33
rect 20 26 31 30
rect 25 23 31 26
rect 25 21 26 23
rect 28 21 31 23
rect 25 18 31 21
rect 41 44 55 46
rect 41 42 52 44
rect 54 42 55 44
rect 50 40 55 42
rect 41 34 46 36
rect 41 32 42 34
rect 44 32 46 34
rect 50 33 54 40
rect 41 30 46 32
rect 42 22 46 30
rect 42 18 55 22
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 10 19 12 30
rect 21 14 23 25
rect 31 14 33 25
rect 41 16 43 27
rect 53 23 55 30
<< pmos >>
rect 9 42 11 64
rect 19 42 21 64
rect 29 42 31 64
rect 40 42 42 64
rect 51 50 53 60
<< polyct0 >>
rect 28 35 30 37
<< polyct1 >>
rect 52 42 54 44
rect 4 35 6 37
rect 42 32 44 34
<< ndifct0 >>
rect 4 21 6 23
rect 16 20 18 22
rect 36 21 38 23
rect 58 26 60 28
rect 47 12 49 14
<< ndifct1 >>
rect 26 21 28 23
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 60 6 62
rect 14 44 16 46
rect 35 44 37 46
rect 45 60 47 62
rect 56 52 58 54
<< pdifct1 >>
rect 24 59 26 61
<< alu0 >>
rect 3 62 7 68
rect 3 60 4 62
rect 6 60 7 62
rect 3 58 7 60
rect 43 62 49 68
rect 43 60 45 62
rect 47 60 49 62
rect 43 59 49 60
rect 11 46 17 48
rect 11 44 14 46
rect 16 44 17 46
rect 11 42 17 44
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 12 7 21
rect 11 23 15 42
rect 27 54 62 55
rect 27 52 56 54
rect 58 52 62 54
rect 27 51 62 52
rect 27 37 31 51
rect 27 35 28 37
rect 30 35 31 37
rect 27 33 31 35
rect 34 46 38 48
rect 34 44 35 46
rect 37 44 38 46
rect 11 22 20 23
rect 11 20 16 22
rect 18 20 20 22
rect 11 19 20 20
rect 34 25 38 44
rect 34 23 39 25
rect 34 21 36 23
rect 38 21 39 23
rect 34 19 39 21
rect 58 29 62 51
rect 56 28 62 29
rect 56 26 58 28
rect 60 26 62 28
rect 56 25 62 26
rect 45 14 51 15
rect 45 12 47 14
rect 49 12 51 14
<< labels >>
rlabel alu0 15 21 15 21 6 a0n
rlabel alu0 29 44 29 44 6 sn
rlabel alu0 14 45 14 45 6 a0n
rlabel alu0 36 33 36 33 6 a1n
rlabel alu0 60 40 60 40 6 sn
rlabel alu0 44 53 44 53 6 sn
rlabel alu1 4 44 4 44 6 a0
rlabel alu1 12 60 12 60 6 a0
rlabel alu1 20 36 20 36 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 28 44 28 6 a1
rlabel alu1 44 44 44 44 6 s
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 20 52 20 6 a1
rlabel alu1 52 40 52 40 6 s
<< end >>
