magic
tech scmos
timestamp 1199202447
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 66 11 71
rect 16 66 18 71
rect 26 66 28 71
rect 33 66 35 71
rect 45 62 51 64
rect 45 60 47 62
rect 49 60 51 62
rect 45 58 51 60
rect 45 55 47 58
rect 9 47 11 50
rect 2 45 11 47
rect 2 43 4 45
rect 6 43 8 45
rect 2 41 8 43
rect 16 41 18 50
rect 26 47 28 50
rect 23 45 29 47
rect 23 43 25 45
rect 27 43 29 45
rect 23 41 29 43
rect 6 27 8 41
rect 12 39 18 41
rect 12 37 14 39
rect 16 37 18 39
rect 33 40 35 50
rect 45 46 47 49
rect 45 44 52 46
rect 33 38 46 40
rect 12 35 28 37
rect 16 29 22 31
rect 16 27 18 29
rect 20 27 22 29
rect 6 25 11 27
rect 9 22 11 25
rect 16 25 22 27
rect 16 22 18 25
rect 26 22 28 35
rect 33 36 42 38
rect 44 36 46 38
rect 33 34 46 36
rect 33 22 35 34
rect 50 30 52 44
rect 45 28 52 30
rect 45 25 47 28
rect 45 15 47 19
rect 9 10 11 15
rect 16 10 18 15
rect 26 10 28 15
rect 33 10 35 15
<< ndif >>
rect 37 22 45 25
rect 2 19 9 22
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 15 16 22
rect 18 20 26 22
rect 18 18 21 20
rect 23 18 26 20
rect 18 15 26 18
rect 28 15 33 22
rect 35 19 45 22
rect 47 23 54 25
rect 47 21 50 23
rect 52 21 54 23
rect 47 19 54 21
rect 35 15 43 19
rect 37 11 43 15
rect 37 9 39 11
rect 41 9 43 11
rect 37 7 43 9
<< pdif >>
rect 37 71 43 73
rect 37 69 39 71
rect 41 69 43 71
rect 37 66 43 69
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 50 9 62
rect 11 50 16 66
rect 18 54 26 66
rect 18 52 21 54
rect 23 52 26 54
rect 18 50 26 52
rect 28 50 33 66
rect 35 55 43 66
rect 35 50 45 55
rect 37 49 45 50
rect 47 53 54 55
rect 47 51 50 53
rect 52 51 54 53
rect 47 49 54 51
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 39 71
rect 41 69 58 71
rect -2 68 58 69
rect 45 62 51 63
rect 11 60 47 62
rect 49 60 51 62
rect 11 58 51 60
rect 11 55 15 58
rect 2 50 15 55
rect 19 52 21 54
rect 23 52 38 54
rect 19 50 38 52
rect 2 45 8 50
rect 2 43 4 45
rect 6 43 8 45
rect 2 42 8 43
rect 23 45 30 46
rect 23 43 25 45
rect 27 43 30 45
rect 23 42 30 43
rect 12 39 18 40
rect 12 38 14 39
rect 2 37 14 38
rect 16 37 18 39
rect 2 34 18 37
rect 2 25 6 34
rect 26 30 30 42
rect 16 29 30 30
rect 16 27 18 29
rect 20 27 30 29
rect 16 26 30 27
rect 34 22 38 50
rect 17 20 38 22
rect 17 18 21 20
rect 23 18 38 20
rect 17 17 38 18
rect -2 11 58 12
rect -2 9 39 11
rect 41 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 15 11 22
rect 16 15 18 22
rect 26 15 28 22
rect 33 15 35 22
rect 45 19 47 25
<< pmos >>
rect 9 50 11 66
rect 16 50 18 66
rect 26 50 28 66
rect 33 50 35 66
rect 45 49 47 55
<< polyct0 >>
rect 42 36 44 38
<< polyct1 >>
rect 47 60 49 62
rect 4 43 6 45
rect 25 43 27 45
rect 14 37 16 39
rect 18 27 20 29
<< ndifct0 >>
rect 4 17 6 19
rect 50 21 52 23
<< ndifct1 >>
rect 21 18 23 20
rect 39 9 41 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 62 6 64
rect 50 51 52 53
<< pdifct1 >>
rect 39 69 41 71
rect 21 52 23 54
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 3 60 7 62
rect 19 54 25 55
rect 49 53 53 55
rect 49 51 50 53
rect 52 51 53 53
rect 49 40 53 51
rect 41 38 53 40
rect 41 36 42 38
rect 44 36 53 38
rect 41 34 53 36
rect 3 19 7 21
rect 3 17 4 19
rect 6 17 7 19
rect 49 23 53 34
rect 49 21 50 23
rect 52 21 53 23
rect 49 19 53 21
rect 3 12 7 17
<< labels >>
rlabel alu0 47 37 47 37 6 sn
rlabel alu0 51 37 51 37 6 sn
rlabel alu1 4 28 4 28 6 a0
rlabel alu1 4 52 4 52 6 s
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 36 12 36 6 a0
rlabel alu1 20 28 20 28 6 a1
rlabel alu1 12 52 12 52 6 s
rlabel alu1 20 60 20 60 6 s
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 36 28 36 6 a1
rlabel alu1 36 32 36 32 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 60 36 60 6 s
rlabel alu1 28 60 28 60 6 s
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 60 44 60 6 s
<< end >>
