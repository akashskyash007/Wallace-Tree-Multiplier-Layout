magic
tech scmos
timestamp 1199543719
<< ab >>
rect 0 0 110 100
<< nwell >>
rect -5 48 115 105
<< pwell >>
rect -5 -5 115 48
<< poly >>
rect 15 94 17 98
rect 27 85 29 89
rect 39 85 41 89
rect 51 85 53 89
rect 63 85 65 89
rect 77 85 79 89
rect 87 85 89 89
rect 97 85 99 89
rect 15 43 17 55
rect 27 43 29 63
rect 39 43 41 63
rect 51 43 53 63
rect 63 43 65 61
rect 15 41 23 43
rect 15 39 19 41
rect 21 39 23 41
rect 15 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 57 41 65 43
rect 57 39 59 41
rect 61 39 65 41
rect 77 53 79 56
rect 87 53 89 56
rect 77 51 83 53
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 87 51 93 53
rect 87 49 89 51
rect 91 49 93 51
rect 87 47 93 49
rect 77 39 79 47
rect 87 39 89 47
rect 57 37 65 39
rect 73 37 79 39
rect 85 37 89 39
rect 97 43 99 55
rect 97 41 103 43
rect 97 39 99 41
rect 101 39 103 41
rect 97 37 103 39
rect 15 34 17 37
rect 29 33 31 37
rect 39 33 41 37
rect 49 33 51 37
rect 61 29 63 37
rect 73 25 75 37
rect 85 25 87 37
rect 97 25 99 37
rect 15 10 17 14
rect 29 13 31 17
rect 39 13 41 17
rect 49 13 51 17
rect 61 13 63 17
rect 73 13 75 17
rect 85 13 87 17
rect 97 13 99 17
<< ndif >>
rect 7 31 15 34
rect 7 29 9 31
rect 11 29 15 31
rect 7 14 15 29
rect 17 33 27 34
rect 17 17 29 33
rect 31 17 39 33
rect 41 17 49 33
rect 51 29 56 33
rect 51 21 61 29
rect 51 19 55 21
rect 57 19 61 21
rect 51 17 61 19
rect 63 25 70 29
rect 63 21 73 25
rect 63 19 67 21
rect 69 19 73 21
rect 63 17 73 19
rect 75 17 85 25
rect 87 21 97 25
rect 87 19 91 21
rect 93 19 97 21
rect 87 17 97 19
rect 99 21 107 25
rect 99 19 103 21
rect 105 19 107 21
rect 99 17 107 19
rect 17 14 27 17
rect 21 11 27 14
rect 77 11 83 17
rect 21 9 23 11
rect 25 9 27 11
rect 21 7 27 9
rect 77 9 79 11
rect 81 9 83 11
rect 77 7 83 9
<< pdif >>
rect 7 81 15 94
rect 7 79 9 81
rect 11 79 15 81
rect 7 71 15 79
rect 7 69 9 71
rect 11 69 15 71
rect 7 61 15 69
rect 7 59 9 61
rect 11 59 15 61
rect 7 55 15 59
rect 17 85 24 94
rect 43 91 49 93
rect 43 89 45 91
rect 47 89 49 91
rect 43 85 49 89
rect 17 81 27 85
rect 17 79 21 81
rect 23 79 27 81
rect 17 63 27 79
rect 29 81 39 85
rect 29 79 33 81
rect 35 79 39 81
rect 29 63 39 79
rect 41 63 51 85
rect 53 81 63 85
rect 53 79 57 81
rect 59 79 63 81
rect 53 63 63 79
rect 17 55 24 63
rect 56 61 63 63
rect 65 71 77 85
rect 65 69 69 71
rect 71 69 77 71
rect 65 61 77 69
rect 67 59 69 61
rect 71 59 77 61
rect 67 57 77 59
rect 72 56 77 57
rect 79 56 87 85
rect 89 56 97 85
rect 92 55 97 56
rect 99 81 107 85
rect 99 79 103 81
rect 105 79 107 81
rect 99 55 107 79
<< alu1 >>
rect -2 95 112 100
rect -2 93 57 95
rect 59 93 69 95
rect 71 93 81 95
rect 83 93 93 95
rect 95 93 112 95
rect -2 91 112 93
rect -2 89 45 91
rect 47 89 112 91
rect -2 88 112 89
rect 8 81 12 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 71 12 79
rect 20 81 24 88
rect 20 79 21 81
rect 23 79 24 81
rect 20 77 24 79
rect 31 81 107 82
rect 31 79 33 81
rect 35 79 57 81
rect 59 79 103 81
rect 105 79 107 81
rect 31 78 107 79
rect 8 69 9 71
rect 11 69 12 71
rect 8 61 12 69
rect 8 59 9 61
rect 11 59 12 61
rect 8 31 12 59
rect 8 29 9 31
rect 11 29 12 31
rect 8 17 12 29
rect 18 41 22 43
rect 18 39 19 41
rect 21 39 22 41
rect 18 22 22 39
rect 28 41 32 73
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 41 42 73
rect 38 39 39 41
rect 41 39 42 41
rect 38 27 42 39
rect 48 41 52 73
rect 48 39 49 41
rect 51 39 52 41
rect 48 37 52 39
rect 58 41 62 73
rect 58 39 59 41
rect 61 39 62 41
rect 58 37 62 39
rect 68 71 72 73
rect 68 69 69 71
rect 71 69 72 71
rect 68 61 72 69
rect 68 59 69 61
rect 71 59 72 61
rect 68 32 72 59
rect 54 28 72 32
rect 78 51 82 73
rect 78 49 79 51
rect 81 49 82 51
rect 54 22 58 28
rect 78 27 82 49
rect 88 51 92 73
rect 88 49 89 51
rect 91 49 92 51
rect 88 27 92 49
rect 98 41 102 73
rect 98 39 99 41
rect 101 39 102 41
rect 98 27 102 39
rect 18 21 58 22
rect 18 19 55 21
rect 57 19 58 21
rect 18 18 58 19
rect 65 21 95 22
rect 65 19 67 21
rect 69 19 91 21
rect 93 19 95 21
rect 65 18 95 19
rect 102 21 106 23
rect 102 19 103 21
rect 105 19 106 21
rect 54 17 58 18
rect 102 12 106 19
rect -2 11 112 12
rect -2 9 23 11
rect 25 9 79 11
rect 81 9 112 11
rect -2 7 35 9
rect 37 7 45 9
rect 47 7 55 9
rect 57 7 66 9
rect 68 7 93 9
rect 95 7 101 9
rect 103 7 112 9
rect -2 0 112 7
<< ptie >>
rect 33 9 70 11
rect 33 7 35 9
rect 37 7 45 9
rect 47 7 55 9
rect 57 7 66 9
rect 68 7 70 9
rect 91 9 105 11
rect 91 7 93 9
rect 95 7 101 9
rect 103 7 105 9
rect 33 5 70 7
rect 91 5 105 7
<< ntie >>
rect 55 95 97 97
rect 55 93 57 95
rect 59 93 69 95
rect 71 93 81 95
rect 83 93 93 95
rect 95 93 97 95
rect 55 91 97 93
<< nmos >>
rect 15 14 17 34
rect 29 17 31 33
rect 39 17 41 33
rect 49 17 51 33
rect 61 17 63 29
rect 73 17 75 25
rect 85 17 87 25
rect 97 17 99 25
<< pmos >>
rect 15 55 17 94
rect 27 63 29 85
rect 39 63 41 85
rect 51 63 53 85
rect 63 61 65 85
rect 77 56 79 85
rect 87 56 89 85
rect 97 55 99 85
<< polyct1 >>
rect 19 39 21 41
rect 29 39 31 41
rect 39 39 41 41
rect 49 39 51 41
rect 59 39 61 41
rect 79 49 81 51
rect 89 49 91 51
rect 99 39 101 41
<< ndifct1 >>
rect 9 29 11 31
rect 55 19 57 21
rect 67 19 69 21
rect 91 19 93 21
rect 103 19 105 21
rect 23 9 25 11
rect 79 9 81 11
<< ntiect1 >>
rect 57 93 59 95
rect 69 93 71 95
rect 81 93 83 95
rect 93 93 95 95
<< ptiect1 >>
rect 35 7 37 9
rect 45 7 47 9
rect 55 7 57 9
rect 66 7 68 9
rect 93 7 95 9
rect 101 7 103 9
<< pdifct1 >>
rect 9 79 11 81
rect 9 69 11 71
rect 9 59 11 61
rect 45 89 47 91
rect 21 79 23 81
rect 33 79 35 81
rect 57 79 59 81
rect 69 69 71 71
rect 69 59 71 61
rect 103 79 105 81
<< labels >>
rlabel alu1 10 50 10 50 6 q
rlabel alu1 40 50 40 50 6 i1
rlabel alu1 30 50 30 50 6 i0
rlabel alu1 50 55 50 55 6 i2
rlabel alu1 55 6 55 6 6 vss
rlabel polyct1 80 50 80 50 6 i3
rlabel alu1 60 55 60 55 6 i6
rlabel alu1 55 94 55 94 6 vdd
rlabel polyct1 90 50 90 50 6 i4
rlabel alu1 100 50 100 50 6 i5
<< end >>
