magic
tech scmos
timestamp 1199203270
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 31 66 33 70
rect 38 66 40 70
rect 45 66 47 70
rect 55 66 57 70
rect 62 66 64 70
rect 69 66 71 70
rect 9 57 11 61
rect 19 59 21 64
rect 9 35 11 38
rect 19 35 21 38
rect 31 35 33 38
rect 9 33 21 35
rect 9 31 17 33
rect 19 31 21 33
rect 9 29 21 31
rect 28 33 34 35
rect 28 31 30 33
rect 32 31 34 33
rect 28 29 34 31
rect 9 26 11 29
rect 29 18 31 29
rect 38 27 40 38
rect 45 35 47 38
rect 55 35 57 38
rect 45 33 57 35
rect 51 31 53 33
rect 55 31 57 33
rect 51 29 57 31
rect 38 25 47 27
rect 38 23 43 25
rect 45 23 47 25
rect 38 21 47 23
rect 39 18 41 21
rect 52 18 54 29
rect 62 27 64 38
rect 69 35 71 38
rect 69 33 78 35
rect 72 31 74 33
rect 76 31 78 33
rect 72 29 78 31
rect 62 25 68 27
rect 62 23 64 25
rect 66 23 68 25
rect 62 21 68 23
rect 9 2 11 6
rect 29 3 31 8
rect 39 3 41 8
rect 52 3 54 8
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 6 9 13
rect 11 18 27 26
rect 11 16 14 18
rect 16 16 29 18
rect 11 12 29 16
rect 11 10 24 12
rect 26 10 29 12
rect 11 8 14 10
rect 16 8 29 10
rect 31 16 39 18
rect 31 14 34 16
rect 36 14 39 16
rect 31 8 39 14
rect 41 8 52 18
rect 54 16 61 18
rect 54 14 57 16
rect 59 14 61 16
rect 54 12 61 14
rect 54 8 59 12
rect 11 6 27 8
rect 43 7 50 8
rect 43 5 45 7
rect 47 5 50 7
rect 43 3 50 5
<< pdif >>
rect 23 64 31 66
rect 23 62 25 64
rect 27 62 31 64
rect 23 59 31 62
rect 14 57 19 59
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 48 9 53
rect 2 46 4 48
rect 6 46 9 48
rect 2 38 9 46
rect 11 49 19 57
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 57 31 59
rect 21 55 25 57
rect 27 55 31 57
rect 21 38 31 55
rect 33 38 38 66
rect 40 38 45 66
rect 47 57 55 66
rect 47 55 50 57
rect 52 55 55 57
rect 47 50 55 55
rect 47 48 50 50
rect 52 48 55 50
rect 47 38 55 48
rect 57 38 62 66
rect 64 38 69 66
rect 71 64 78 66
rect 71 62 74 64
rect 76 62 78 64
rect 71 56 78 62
rect 71 54 74 56
rect 76 54 78 56
rect 71 38 78 54
<< alu1 >>
rect -2 67 82 72
rect -2 65 7 67
rect 9 65 82 67
rect -2 64 82 65
rect 13 49 17 51
rect 13 47 14 49
rect 16 47 17 49
rect 13 42 17 47
rect 2 40 14 42
rect 16 40 17 42
rect 2 38 17 40
rect 2 26 6 38
rect 58 42 62 51
rect 33 38 78 42
rect 33 34 39 38
rect 28 33 39 34
rect 28 31 30 33
rect 32 31 39 33
rect 28 30 39 31
rect 49 33 63 34
rect 49 31 53 33
rect 55 31 63 33
rect 49 30 63 31
rect 74 33 78 38
rect 76 31 78 33
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 17 7 22
rect 74 29 78 31
rect 41 25 70 26
rect 41 23 43 25
rect 45 23 64 25
rect 66 23 70 25
rect 41 22 70 23
rect 2 15 4 17
rect 6 15 7 17
rect 2 13 7 15
rect 66 13 70 22
rect -2 7 82 8
rect -2 5 45 7
rect 47 5 73 7
rect 75 5 82 7
rect -2 0 82 5
<< ptie >>
rect 71 7 77 24
rect 71 5 73 7
rect 75 5 77 7
rect 71 3 77 5
<< ntie >>
rect 3 67 13 69
rect 3 65 7 67
rect 9 65 13 67
rect 3 63 13 65
<< nmos >>
rect 9 6 11 26
rect 29 8 31 18
rect 39 8 41 18
rect 52 8 54 18
<< pmos >>
rect 9 38 11 57
rect 19 38 21 59
rect 31 38 33 66
rect 38 38 40 66
rect 45 38 47 66
rect 55 38 57 66
rect 62 38 64 66
rect 69 38 71 66
<< polyct0 >>
rect 17 31 19 33
<< polyct1 >>
rect 30 31 32 33
rect 53 31 55 33
rect 43 23 45 25
rect 74 31 76 33
rect 64 23 66 25
<< ndifct0 >>
rect 14 16 16 18
rect 24 10 26 12
rect 14 8 16 10
rect 34 14 36 16
rect 57 14 59 16
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
rect 45 5 47 7
<< ntiect1 >>
rect 7 65 9 67
<< ptiect1 >>
rect 73 5 75 7
<< pdifct0 >>
rect 25 62 27 64
rect 4 53 6 55
rect 4 46 6 48
rect 25 55 27 57
rect 50 55 52 57
rect 50 48 52 50
rect 74 62 76 64
rect 74 54 76 56
<< pdifct1 >>
rect 14 47 16 49
rect 14 40 16 42
<< alu0 >>
rect 2 55 8 64
rect 2 53 4 55
rect 6 53 8 55
rect 23 62 25 64
rect 27 62 29 64
rect 23 57 29 62
rect 73 62 74 64
rect 76 62 77 64
rect 23 55 25 57
rect 27 55 29 57
rect 23 54 29 55
rect 49 57 53 59
rect 49 55 50 57
rect 52 55 53 57
rect 2 48 8 53
rect 2 46 4 48
rect 6 46 8 48
rect 2 45 8 46
rect 49 50 53 55
rect 73 56 77 62
rect 73 54 74 56
rect 76 54 77 56
rect 73 52 77 54
rect 21 48 50 50
rect 52 48 53 50
rect 21 46 53 48
rect 21 34 25 46
rect 15 33 25 34
rect 15 31 17 33
rect 19 31 25 33
rect 15 30 25 31
rect 72 30 74 38
rect 21 25 25 30
rect 21 21 36 25
rect 13 18 17 20
rect 13 16 14 18
rect 16 16 17 18
rect 13 10 17 16
rect 32 17 36 21
rect 32 16 61 17
rect 32 14 34 16
rect 36 14 57 16
rect 59 14 61 16
rect 13 8 14 10
rect 16 8 17 10
rect 23 12 27 14
rect 32 13 61 14
rect 23 10 24 12
rect 26 10 27 12
rect 23 8 27 10
<< labels >>
rlabel alu0 20 32 20 32 6 zn
rlabel alu0 51 52 51 52 6 zn
rlabel alu0 46 15 46 15 6 zn
rlabel alu1 4 24 4 24 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 36 36 36 36 6 a
rlabel alu1 40 4 40 4 6 vss
rlabel polyct1 44 24 44 24 6 b
rlabel alu1 52 24 52 24 6 b
rlabel alu1 52 32 52 32 6 c
rlabel alu1 52 40 52 40 6 a
rlabel alu1 44 40 44 40 6 a
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 68 16 68 16 6 b
rlabel alu1 60 24 60 24 6 b
rlabel alu1 60 32 60 32 6 c
rlabel alu1 76 32 76 32 6 a
rlabel alu1 68 40 68 40 6 a
rlabel alu1 60 44 60 44 6 a
<< end >>
