magic
tech scmos
timestamp 1199202491
<< ab >>
rect 0 0 224 80
<< nwell >>
rect -5 36 229 88
<< pwell >>
rect -5 -8 229 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 59 71 81 73
rect 59 65 61 71
rect 69 68 71 71
rect 79 68 81 71
rect 139 72 205 74
rect 139 69 141 72
rect 49 63 61 65
rect 49 60 51 63
rect 59 60 61 63
rect 89 64 91 69
rect 99 67 141 69
rect 99 64 101 67
rect 109 64 111 67
rect 119 64 121 67
rect 129 64 131 67
rect 139 64 141 67
rect 149 64 151 68
rect 163 64 165 68
rect 173 64 175 68
rect 183 64 185 68
rect 193 64 195 68
rect 203 64 205 72
rect 213 58 215 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 41 39
rect 49 38 51 42
rect 59 38 61 42
rect 69 38 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 9 35 11 37
rect 13 35 19 37
rect 21 35 41 37
rect 9 33 41 35
rect 79 37 91 39
rect 99 38 101 42
rect 109 38 111 42
rect 119 39 121 42
rect 79 35 85 37
rect 87 35 91 37
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 33
rect 49 30 51 34
rect 59 30 61 34
rect 69 30 71 34
rect 79 33 91 35
rect 119 37 125 39
rect 129 37 131 42
rect 139 37 141 42
rect 149 39 151 42
rect 163 39 165 42
rect 173 39 175 42
rect 183 39 185 42
rect 193 39 195 42
rect 149 37 195 39
rect 203 39 205 42
rect 213 39 215 42
rect 119 35 121 37
rect 123 35 125 37
rect 79 30 81 33
rect 89 30 91 33
rect 99 30 101 34
rect 109 30 111 34
rect 119 33 125 35
rect 149 35 151 37
rect 153 35 159 37
rect 161 35 181 37
rect 149 33 181 35
rect 79 13 81 17
rect 89 14 91 17
rect 99 14 101 17
rect 109 14 111 17
rect 89 12 111 14
rect 19 7 21 12
rect 29 7 31 12
rect 39 7 41 12
rect 49 8 51 12
rect 59 8 61 12
rect 69 8 71 12
rect 120 8 122 33
rect 149 30 151 33
rect 159 30 161 33
rect 169 30 171 33
rect 179 30 181 33
rect 203 33 215 39
rect 203 30 205 33
rect 213 30 215 33
rect 49 6 122 8
rect 149 11 151 16
rect 159 11 161 16
rect 169 11 171 16
rect 179 11 181 16
rect 203 14 205 19
rect 213 15 215 19
<< ndif >>
rect 11 24 19 30
rect 11 22 14 24
rect 16 22 19 24
rect 11 16 19 22
rect 11 14 14 16
rect 16 14 19 16
rect 11 12 19 14
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 21 29 26
rect 21 19 24 21
rect 26 19 29 21
rect 21 12 29 19
rect 31 16 39 30
rect 31 14 34 16
rect 36 14 39 16
rect 31 12 39 14
rect 41 28 49 30
rect 41 26 44 28
rect 46 26 49 28
rect 41 21 49 26
rect 41 19 44 21
rect 46 19 49 21
rect 41 12 49 19
rect 51 28 59 30
rect 51 26 54 28
rect 56 26 59 28
rect 51 12 59 26
rect 61 20 69 30
rect 61 18 64 20
rect 66 18 69 20
rect 61 12 69 18
rect 71 28 79 30
rect 71 26 74 28
rect 76 26 79 28
rect 71 21 79 26
rect 71 19 74 21
rect 76 19 79 21
rect 71 17 79 19
rect 81 21 89 30
rect 81 19 84 21
rect 86 19 89 21
rect 81 17 89 19
rect 91 28 99 30
rect 91 26 94 28
rect 96 26 99 28
rect 91 17 99 26
rect 101 21 109 30
rect 101 19 104 21
rect 106 19 109 21
rect 101 17 109 19
rect 111 28 118 30
rect 111 26 114 28
rect 116 26 118 28
rect 111 24 118 26
rect 111 17 116 24
rect 71 12 76 17
rect 141 16 149 30
rect 151 28 159 30
rect 151 26 154 28
rect 156 26 159 28
rect 151 21 159 26
rect 151 19 154 21
rect 156 19 159 21
rect 151 16 159 19
rect 161 20 169 30
rect 161 18 164 20
rect 166 18 169 20
rect 161 16 169 18
rect 171 28 179 30
rect 171 26 174 28
rect 176 26 179 28
rect 171 21 179 26
rect 171 19 174 21
rect 176 19 179 21
rect 171 16 179 19
rect 181 28 189 30
rect 181 26 184 28
rect 186 26 189 28
rect 181 20 189 26
rect 181 18 184 20
rect 186 18 189 20
rect 195 23 203 30
rect 195 21 198 23
rect 200 21 203 23
rect 195 19 203 21
rect 205 28 213 30
rect 205 26 208 28
rect 210 26 213 28
rect 205 19 213 26
rect 215 23 222 30
rect 215 21 218 23
rect 220 21 222 23
rect 215 19 222 21
rect 181 16 189 18
rect 141 11 147 16
rect 141 9 143 11
rect 145 9 147 11
rect 141 7 147 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 42 19 59
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 42 39 59
rect 41 60 46 70
rect 64 60 69 68
rect 41 53 49 60
rect 41 51 44 53
rect 46 51 49 53
rect 41 46 49 51
rect 41 44 44 46
rect 46 44 49 46
rect 41 42 49 44
rect 51 53 59 60
rect 51 51 54 53
rect 56 51 59 53
rect 51 46 59 51
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 58 69 60
rect 61 56 64 58
rect 66 56 69 58
rect 61 51 69 56
rect 61 49 64 51
rect 66 49 69 51
rect 61 42 69 49
rect 71 53 79 68
rect 71 51 74 53
rect 76 51 79 53
rect 71 46 79 51
rect 71 44 74 46
rect 76 44 79 46
rect 71 42 79 44
rect 81 64 86 68
rect 81 62 89 64
rect 81 60 84 62
rect 86 60 89 62
rect 81 42 89 60
rect 91 46 99 64
rect 91 44 94 46
rect 96 44 99 46
rect 91 42 99 44
rect 101 54 109 64
rect 101 52 104 54
rect 106 52 109 54
rect 101 42 109 52
rect 111 46 119 64
rect 111 44 114 46
rect 116 44 119 46
rect 111 42 119 44
rect 121 54 129 64
rect 121 52 124 54
rect 126 52 129 54
rect 121 42 129 52
rect 131 46 139 64
rect 131 44 134 46
rect 136 44 139 46
rect 131 42 139 44
rect 141 53 149 64
rect 141 51 144 53
rect 146 51 149 53
rect 141 46 149 51
rect 141 44 144 46
rect 146 44 149 46
rect 141 42 149 44
rect 151 62 163 64
rect 151 60 158 62
rect 160 60 163 62
rect 151 42 163 60
rect 165 46 173 64
rect 165 44 168 46
rect 170 44 173 46
rect 165 42 173 44
rect 175 62 183 64
rect 175 60 178 62
rect 180 60 183 62
rect 175 42 183 60
rect 185 46 193 64
rect 185 44 188 46
rect 190 44 193 46
rect 185 42 193 44
rect 195 62 203 64
rect 195 60 198 62
rect 200 60 203 62
rect 195 42 203 60
rect 205 58 210 64
rect 205 53 213 58
rect 205 51 208 53
rect 210 51 213 53
rect 205 46 213 51
rect 205 44 208 46
rect 210 44 213 46
rect 205 42 213 44
rect 215 56 222 58
rect 215 54 218 56
rect 220 54 222 56
rect 215 48 222 54
rect 215 46 218 48
rect 220 46 222 48
rect 215 42 222 46
<< alu1 >>
rect -2 81 226 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 203 81
rect 205 79 211 81
rect 213 79 219 81
rect 221 79 226 81
rect -2 68 226 79
rect 2 37 22 39
rect 2 35 11 37
rect 13 35 19 37
rect 21 35 22 37
rect 2 33 22 35
rect 2 17 6 33
rect 53 53 57 55
rect 53 51 54 53
rect 56 51 57 53
rect 53 46 57 51
rect 73 53 78 56
rect 73 51 74 53
rect 76 51 78 53
rect 53 44 54 46
rect 56 44 57 46
rect 53 30 57 44
rect 73 46 78 51
rect 73 44 74 46
rect 76 44 78 46
rect 73 30 78 44
rect 92 46 98 47
rect 112 46 118 47
rect 132 46 138 47
rect 92 44 94 46
rect 96 44 114 46
rect 116 44 134 46
rect 136 44 138 46
rect 92 42 138 44
rect 98 30 102 42
rect 119 37 135 38
rect 119 35 121 37
rect 123 35 135 37
rect 119 34 135 35
rect 53 28 119 30
rect 53 26 54 28
rect 56 26 74 28
rect 76 26 94 28
rect 96 26 114 28
rect 116 26 119 28
rect 129 26 135 34
rect 146 37 166 39
rect 146 35 151 37
rect 153 35 159 37
rect 161 35 166 37
rect 146 33 166 35
rect 53 24 57 26
rect 73 21 78 26
rect 92 25 98 26
rect 112 25 119 26
rect 146 25 150 33
rect 73 19 74 21
rect 76 19 78 21
rect 73 17 78 19
rect -2 11 226 12
rect -2 9 143 11
rect 145 9 226 11
rect -2 1 226 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 203 1
rect 205 -1 211 1
rect 213 -1 219 1
rect 221 -1 226 1
rect -2 -2 226 -1
<< ptie >>
rect 0 1 224 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 203 1
rect 205 -1 211 1
rect 213 -1 219 1
rect 221 -1 224 1
rect 0 -3 224 -1
<< ntie >>
rect 0 81 224 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 203 81
rect 205 79 211 81
rect 213 79 219 81
rect 221 79 224 81
rect 0 77 224 79
<< nmos >>
rect 19 12 21 30
rect 29 12 31 30
rect 39 12 41 30
rect 49 12 51 30
rect 59 12 61 30
rect 69 12 71 30
rect 79 17 81 30
rect 89 17 91 30
rect 99 17 101 30
rect 109 17 111 30
rect 149 16 151 30
rect 159 16 161 30
rect 169 16 171 30
rect 179 16 181 30
rect 203 19 205 30
rect 213 19 215 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 60
rect 59 42 61 60
rect 69 42 71 68
rect 79 42 81 68
rect 89 42 91 64
rect 99 42 101 64
rect 109 42 111 64
rect 119 42 121 64
rect 129 42 131 64
rect 139 42 141 64
rect 149 42 151 64
rect 163 42 165 64
rect 173 42 175 64
rect 183 42 185 64
rect 193 42 195 64
rect 203 42 205 64
rect 213 42 215 58
<< polyct0 >>
rect 85 35 87 37
<< polyct1 >>
rect 11 35 13 37
rect 19 35 21 37
rect 121 35 123 37
rect 151 35 153 37
rect 159 35 161 37
<< ndifct0 >>
rect 14 22 16 24
rect 14 14 16 16
rect 24 26 26 28
rect 24 19 26 21
rect 34 14 36 16
rect 44 26 46 28
rect 44 19 46 21
rect 64 18 66 20
rect 84 19 86 21
rect 104 19 106 21
rect 154 26 156 28
rect 154 19 156 21
rect 164 18 166 20
rect 174 26 176 28
rect 174 19 176 21
rect 184 26 186 28
rect 184 18 186 20
rect 198 21 200 23
rect 208 26 210 28
rect 218 21 220 23
<< ndifct1 >>
rect 54 26 56 28
rect 74 26 76 28
rect 74 19 76 21
rect 94 26 96 28
rect 114 26 116 28
rect 143 9 145 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
rect 171 79 173 81
rect 179 79 181 81
rect 187 79 189 81
rect 195 79 197 81
rect 203 79 205 81
rect 211 79 213 81
rect 219 79 221 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
rect 171 -1 173 1
rect 179 -1 181 1
rect 187 -1 189 1
rect 195 -1 197 1
rect 203 -1 205 1
rect 211 -1 213 1
rect 219 -1 221 1
<< pdifct0 >>
rect 4 51 6 53
rect 4 44 6 46
rect 14 66 16 68
rect 14 59 16 61
rect 24 51 26 53
rect 24 44 26 46
rect 34 66 36 68
rect 34 59 36 61
rect 44 51 46 53
rect 44 44 46 46
rect 64 56 66 58
rect 64 49 66 51
rect 84 60 86 62
rect 104 52 106 54
rect 124 52 126 54
rect 144 51 146 53
rect 144 44 146 46
rect 158 60 160 62
rect 168 44 170 46
rect 178 60 180 62
rect 188 44 190 46
rect 198 60 200 62
rect 208 51 210 53
rect 208 44 210 46
rect 218 54 220 56
rect 218 46 220 48
<< pdifct1 >>
rect 54 51 56 53
rect 54 44 56 46
rect 74 51 76 53
rect 74 44 76 46
rect 94 44 96 46
rect 114 44 116 46
rect 134 44 136 46
<< alu0 >>
rect 13 66 14 68
rect 16 66 17 68
rect 13 61 17 66
rect 13 59 14 61
rect 16 59 17 61
rect 13 57 17 59
rect 33 66 34 68
rect 36 66 37 68
rect 33 61 37 66
rect 33 59 34 61
rect 36 59 37 61
rect 33 57 37 59
rect 43 62 88 63
rect 43 60 84 62
rect 86 60 88 62
rect 43 59 88 60
rect 93 59 154 63
rect 3 53 7 55
rect 3 51 4 53
rect 6 51 7 53
rect 3 46 7 51
rect 23 53 27 55
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 43 53 47 59
rect 63 58 67 59
rect 63 56 64 58
rect 66 56 67 58
rect 43 51 44 53
rect 46 51 47 53
rect 43 46 47 51
rect 3 44 4 46
rect 6 44 24 46
rect 26 44 44 46
rect 46 44 47 46
rect 3 42 47 44
rect 43 30 47 42
rect 23 28 47 30
rect 23 26 24 28
rect 26 26 44 28
rect 46 26 47 28
rect 13 24 17 26
rect 13 22 14 24
rect 16 22 17 24
rect 13 16 17 22
rect 23 21 27 26
rect 23 19 24 21
rect 26 19 27 21
rect 23 17 27 19
rect 43 21 47 26
rect 63 51 67 56
rect 63 49 64 51
rect 66 49 67 51
rect 63 47 67 49
rect 93 55 97 59
rect 150 55 154 59
rect 157 62 161 68
rect 157 60 158 62
rect 160 60 161 62
rect 157 58 161 60
rect 177 62 181 68
rect 177 60 178 62
rect 180 60 181 62
rect 177 58 181 60
rect 196 62 202 68
rect 196 60 198 62
rect 200 60 202 62
rect 196 59 202 60
rect 217 56 221 68
rect 84 51 97 55
rect 102 54 147 55
rect 102 52 104 54
rect 106 52 124 54
rect 126 53 147 54
rect 126 52 144 53
rect 102 51 144 52
rect 146 51 147 53
rect 150 53 211 55
rect 150 51 208 53
rect 210 51 211 53
rect 84 37 88 51
rect 142 47 147 51
rect 142 46 192 47
rect 142 44 144 46
rect 146 44 168 46
rect 170 44 188 46
rect 190 44 192 46
rect 142 43 192 44
rect 207 46 211 51
rect 207 44 208 46
rect 210 44 211 46
rect 217 54 218 56
rect 220 54 221 56
rect 217 48 221 54
rect 217 46 218 48
rect 220 46 221 48
rect 217 44 221 46
rect 84 35 85 37
rect 87 35 88 37
rect 84 33 88 35
rect 173 30 177 43
rect 153 28 177 30
rect 153 26 154 28
rect 156 26 174 28
rect 176 26 177 28
rect 153 22 158 26
rect 43 19 44 21
rect 46 20 68 21
rect 46 19 64 20
rect 43 18 64 19
rect 66 18 68 20
rect 13 14 14 16
rect 16 14 17 16
rect 13 12 17 14
rect 33 16 37 18
rect 43 17 68 18
rect 82 21 158 22
rect 82 19 84 21
rect 86 19 104 21
rect 106 19 154 21
rect 156 19 158 21
rect 82 18 158 19
rect 163 20 167 22
rect 163 18 164 20
rect 166 18 167 20
rect 33 14 34 16
rect 36 14 37 16
rect 33 12 37 14
rect 163 12 167 18
rect 173 21 177 26
rect 173 19 174 21
rect 176 19 177 21
rect 173 17 177 19
rect 183 28 187 30
rect 183 26 184 28
rect 186 26 187 28
rect 183 20 187 26
rect 207 28 211 44
rect 207 26 208 28
rect 210 26 211 28
rect 183 18 184 20
rect 186 18 187 20
rect 183 12 187 18
rect 197 23 201 25
rect 207 24 211 26
rect 197 21 198 23
rect 200 21 201 23
rect 197 12 201 21
rect 217 23 221 25
rect 217 21 218 23
rect 220 21 221 23
rect 217 12 221 21
<< labels >>
rlabel alu0 25 23 25 23 6 a1n
rlabel alu0 25 48 25 48 6 a1n
rlabel alu0 5 48 5 48 6 a1n
rlabel alu0 55 19 55 19 6 a1n
rlabel alu0 65 55 65 55 6 a1n
rlabel alu0 45 40 45 40 6 a1n
rlabel alu0 86 44 86 44 6 sn
rlabel alu0 65 61 65 61 6 a1n
rlabel alu0 120 20 120 20 6 a0n
rlabel alu0 155 24 155 24 6 a0n
rlabel alu0 175 32 175 32 6 a0n
rlabel alu0 144 49 144 49 6 a0n
rlabel alu0 124 53 124 53 6 a0n
rlabel alu0 167 45 167 45 6 a0n
rlabel alu0 209 39 209 39 6 sn
rlabel polyct1 12 36 12 36 6 a1
rlabel polyct1 20 36 20 36 6 a1
rlabel alu1 4 28 4 28 6 a1
rlabel alu1 100 36 100 36 6 z
rlabel alu1 108 28 108 28 6 z
rlabel alu1 92 28 92 28 6 z
rlabel alu1 76 36 76 36 6 z
rlabel alu1 60 28 60 28 6 z
rlabel alu1 68 28 68 28 6 z
rlabel alu1 84 28 84 28 6 z
rlabel alu1 108 44 108 44 6 z
rlabel alu1 112 6 112 6 6 vss
rlabel alu1 116 28 116 28 6 z
rlabel alu1 164 36 164 36 6 a0
rlabel alu1 156 36 156 36 6 a0
rlabel alu1 148 32 148 32 6 a0
rlabel alu1 124 36 124 36 6 s
rlabel alu1 132 32 132 32 6 s
rlabel alu1 132 44 132 44 6 z
rlabel alu1 124 44 124 44 6 z
rlabel alu1 116 44 116 44 6 z
rlabel alu1 112 74 112 74 6 vdd
<< end >>
