magic
tech scmos
timestamp 1199469431
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -2 48 82 104
<< pwell >>
rect -2 -4 82 48
<< poly >>
rect 11 93 13 98
rect 23 93 25 98
rect 31 93 33 98
rect 43 93 45 98
rect 55 93 57 98
rect 67 77 69 82
rect 11 53 13 67
rect 23 53 25 67
rect 31 53 33 67
rect 43 63 45 67
rect 43 61 51 63
rect 43 59 47 61
rect 49 59 51 61
rect 43 57 51 59
rect 11 51 25 53
rect 11 49 19 51
rect 21 49 25 51
rect 11 47 25 49
rect 29 51 39 53
rect 29 49 35 51
rect 37 49 39 51
rect 29 47 39 49
rect 11 31 13 47
rect 21 31 23 47
rect 29 31 31 47
rect 43 40 45 57
rect 55 53 57 67
rect 49 51 57 53
rect 49 49 51 51
rect 53 49 57 51
rect 49 47 57 49
rect 41 37 45 40
rect 41 31 43 37
rect 53 31 55 47
rect 67 43 69 57
rect 59 41 69 43
rect 59 39 61 41
rect 63 40 69 41
rect 63 39 67 40
rect 59 37 67 39
rect 65 33 67 37
rect 11 15 13 19
rect 21 14 23 19
rect 29 14 31 19
rect 41 14 43 19
rect 53 14 55 19
rect 65 18 67 23
<< ndif >>
rect 57 31 65 33
rect 6 25 11 31
rect 3 23 11 25
rect 3 21 5 23
rect 7 21 11 23
rect 3 19 11 21
rect 13 19 21 31
rect 23 19 29 31
rect 31 29 41 31
rect 31 27 35 29
rect 37 27 41 29
rect 31 19 41 27
rect 43 23 53 31
rect 43 21 47 23
rect 49 21 53 23
rect 43 19 53 21
rect 55 29 59 31
rect 61 29 65 31
rect 55 23 65 29
rect 67 31 75 33
rect 67 29 71 31
rect 73 29 75 31
rect 67 27 75 29
rect 67 23 72 27
rect 55 21 59 23
rect 61 21 63 23
rect 55 19 63 21
rect 15 13 19 19
rect 13 11 19 13
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 6 81 11 93
rect 3 79 11 81
rect 3 77 5 79
rect 7 77 11 79
rect 3 71 11 77
rect 3 69 5 71
rect 7 69 11 71
rect 3 67 11 69
rect 13 91 23 93
rect 13 89 17 91
rect 19 89 23 91
rect 13 67 23 89
rect 25 67 31 93
rect 33 71 43 93
rect 33 69 37 71
rect 39 69 43 71
rect 33 67 43 69
rect 45 81 55 93
rect 45 79 49 81
rect 51 79 55 81
rect 45 67 55 79
rect 57 91 65 93
rect 57 89 61 91
rect 63 89 65 91
rect 57 81 65 89
rect 57 79 61 81
rect 63 79 65 81
rect 57 77 65 79
rect 57 67 67 77
rect 59 57 67 67
rect 69 63 74 77
rect 69 61 77 63
rect 69 59 73 61
rect 75 59 77 61
rect 69 57 77 59
<< alu1 >>
rect -2 95 82 100
rect -2 93 73 95
rect 75 93 82 95
rect -2 91 82 93
rect -2 89 17 91
rect 19 89 61 91
rect 63 89 82 91
rect -2 88 82 89
rect 4 81 53 82
rect 4 79 49 81
rect 51 79 53 81
rect 4 77 5 79
rect 7 78 53 79
rect 60 81 64 88
rect 60 79 61 81
rect 63 79 64 81
rect 7 77 8 78
rect 60 77 64 79
rect 4 71 8 77
rect 68 72 73 83
rect 4 69 5 71
rect 7 69 8 71
rect 4 67 8 69
rect 26 71 41 72
rect 26 69 37 71
rect 39 69 41 71
rect 26 68 41 69
rect 46 68 73 72
rect 8 53 12 63
rect 8 51 22 53
rect 8 49 19 51
rect 21 49 22 51
rect 8 47 22 49
rect 8 37 12 47
rect 26 32 30 68
rect 38 53 42 63
rect 46 61 52 68
rect 46 59 47 61
rect 49 59 52 61
rect 46 57 52 59
rect 57 61 77 62
rect 57 59 73 61
rect 75 59 77 61
rect 57 58 77 59
rect 34 51 55 53
rect 34 49 35 51
rect 37 49 51 51
rect 53 49 55 51
rect 34 47 55 49
rect 38 37 42 47
rect 48 41 64 43
rect 48 39 61 41
rect 63 39 64 41
rect 48 37 64 39
rect 48 32 52 37
rect 68 33 72 58
rect 26 29 52 32
rect 26 28 35 29
rect 33 27 35 28
rect 37 28 52 29
rect 58 31 62 33
rect 58 29 59 31
rect 61 29 62 31
rect 37 27 39 28
rect 33 26 39 27
rect 3 23 9 24
rect 3 21 5 23
rect 7 21 9 23
rect 45 23 51 24
rect 45 21 47 23
rect 49 21 51 23
rect 3 17 51 21
rect 58 23 62 29
rect 68 31 74 33
rect 68 29 71 31
rect 73 29 74 31
rect 68 27 74 29
rect 58 21 59 23
rect 61 21 62 23
rect 58 12 62 21
rect -2 11 82 12
rect -2 9 15 11
rect 17 9 82 11
rect -2 7 82 9
rect -2 5 27 7
rect 29 5 37 7
rect 39 5 82 7
rect -2 0 82 5
<< ptie >>
rect 25 7 41 9
rect 25 5 27 7
rect 29 5 37 7
rect 39 5 41 7
rect 25 3 41 5
<< ntie >>
rect 71 95 77 97
rect 71 93 73 95
rect 75 93 77 95
rect 71 91 77 93
<< nmos >>
rect 11 19 13 31
rect 21 19 23 31
rect 29 19 31 31
rect 41 19 43 31
rect 53 19 55 31
rect 65 23 67 33
<< pmos >>
rect 11 67 13 93
rect 23 67 25 93
rect 31 67 33 93
rect 43 67 45 93
rect 55 67 57 93
rect 67 57 69 77
<< polyct1 >>
rect 47 59 49 61
rect 19 49 21 51
rect 35 49 37 51
rect 51 49 53 51
rect 61 39 63 41
<< ndifct1 >>
rect 5 21 7 23
rect 35 27 37 29
rect 47 21 49 23
rect 59 29 61 31
rect 71 29 73 31
rect 59 21 61 23
rect 15 9 17 11
<< ntiect1 >>
rect 73 93 75 95
<< ptiect1 >>
rect 27 5 29 7
rect 37 5 39 7
<< pdifct1 >>
rect 5 77 7 79
rect 5 69 7 71
rect 17 89 19 91
rect 37 69 39 71
rect 49 79 51 81
rect 61 89 63 91
rect 61 79 63 81
rect 73 59 75 61
<< labels >>
rlabel alu1 6 20 6 20 6 n4
rlabel alu1 10 50 10 50 6 a
rlabel alu1 6 74 6 74 6 n2
rlabel polyct1 20 50 20 50 6 a
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 40 50 40 50 6 b
rlabel alu1 33 70 33 70 6 zn
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 48 20 48 20 6 n4
rlabel alu1 39 30 39 30 6 zn
rlabel alu1 56 40 56 40 6 zn
rlabel alu1 50 50 50 50 6 b
rlabel alu1 60 60 60 60 6 z
rlabel alu1 50 65 50 65 6 c
rlabel alu1 60 70 60 70 6 c
rlabel alu1 28 80 28 80 6 n2
rlabel alu1 70 45 70 45 6 z
rlabel alu1 70 75 70 75 6 c
<< end >>
