magic
tech scmos
timestamp 1199469250
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -2 48 92 104
<< pwell >>
rect -2 -4 92 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 71 91 73 96
rect 47 83 49 88
rect 59 83 61 88
rect 11 52 13 55
rect 23 52 25 55
rect 35 52 37 55
rect 47 52 49 55
rect 11 50 49 52
rect 11 35 13 50
rect 23 48 29 50
rect 31 48 37 50
rect 23 46 37 48
rect 23 35 25 46
rect 35 35 37 46
rect 47 35 49 50
rect 59 43 61 55
rect 71 43 73 55
rect 59 41 73 43
rect 59 39 69 41
rect 71 39 73 41
rect 59 37 73 39
rect 59 33 61 37
rect 71 33 73 37
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 47 12 49 17
rect 59 12 61 17
rect 71 12 73 17
<< ndif >>
rect 3 31 11 35
rect 3 29 5 31
rect 7 29 11 31
rect 3 21 11 29
rect 3 19 5 21
rect 7 19 11 21
rect 3 17 11 19
rect 13 31 23 35
rect 13 29 17 31
rect 19 29 23 31
rect 13 21 23 29
rect 13 19 17 21
rect 19 19 23 21
rect 13 17 23 19
rect 25 31 35 35
rect 25 29 29 31
rect 31 29 35 31
rect 25 21 35 29
rect 25 19 29 21
rect 31 19 35 21
rect 25 17 35 19
rect 37 31 47 35
rect 37 29 41 31
rect 43 29 47 31
rect 37 21 47 29
rect 37 19 41 21
rect 43 19 47 21
rect 37 17 47 19
rect 49 33 57 35
rect 49 31 59 33
rect 49 29 53 31
rect 55 29 59 31
rect 49 21 59 29
rect 49 19 53 21
rect 55 19 59 21
rect 49 17 59 19
rect 61 31 71 33
rect 61 29 65 31
rect 67 29 71 31
rect 61 21 71 29
rect 61 19 65 21
rect 67 19 71 21
rect 61 17 71 19
rect 73 31 82 33
rect 73 29 77 31
rect 79 29 82 31
rect 73 23 82 29
rect 73 21 77 23
rect 79 21 82 23
rect 73 17 82 21
<< pdif >>
rect 3 91 11 94
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 55 11 69
rect 13 71 23 94
rect 13 69 17 71
rect 19 69 23 71
rect 13 63 23 69
rect 13 61 17 63
rect 19 61 23 63
rect 13 55 23 61
rect 25 91 35 94
rect 25 89 29 91
rect 31 89 35 91
rect 25 81 35 89
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 55 35 69
rect 37 83 42 94
rect 66 83 71 91
rect 37 71 47 83
rect 37 69 41 71
rect 43 69 47 71
rect 37 63 47 69
rect 37 61 41 63
rect 43 61 47 63
rect 37 55 47 61
rect 49 81 59 83
rect 49 79 53 81
rect 55 79 59 81
rect 49 71 59 79
rect 49 69 53 71
rect 55 69 59 71
rect 49 55 59 69
rect 61 71 71 83
rect 61 69 65 71
rect 67 69 71 71
rect 61 61 71 69
rect 61 59 65 61
rect 67 59 71 61
rect 61 55 71 59
rect 73 81 82 91
rect 73 79 77 81
rect 79 79 82 81
rect 73 71 82 79
rect 73 69 77 71
rect 79 69 82 71
rect 73 55 82 69
<< alu1 >>
rect -2 95 92 100
rect -2 93 53 95
rect 55 93 92 95
rect -2 91 92 93
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 92 91
rect -2 88 92 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 28 81 32 88
rect 28 79 29 81
rect 31 79 32 81
rect 4 69 5 71
rect 7 69 8 71
rect 4 67 8 69
rect 16 71 22 73
rect 16 69 17 71
rect 19 69 22 71
rect 16 63 22 69
rect 28 71 32 79
rect 52 81 56 88
rect 52 79 53 81
rect 55 79 56 81
rect 28 69 29 71
rect 31 69 32 71
rect 28 67 32 69
rect 38 71 44 73
rect 38 69 41 71
rect 43 69 44 71
rect 16 61 17 63
rect 19 62 22 63
rect 38 63 44 69
rect 52 71 56 79
rect 76 81 80 88
rect 76 79 77 81
rect 79 79 80 81
rect 52 69 53 71
rect 55 69 56 71
rect 52 67 56 69
rect 64 71 68 73
rect 64 69 65 71
rect 67 69 68 71
rect 38 62 41 63
rect 19 61 41 62
rect 43 61 44 63
rect 16 58 44 61
rect 64 61 68 69
rect 76 71 80 79
rect 76 69 77 71
rect 79 69 80 71
rect 76 67 80 69
rect 64 59 65 61
rect 67 59 68 61
rect 16 42 22 58
rect 64 51 68 59
rect 27 50 68 51
rect 27 48 29 50
rect 31 48 68 50
rect 27 47 68 48
rect 16 38 44 42
rect 4 31 8 33
rect 4 29 5 31
rect 7 29 8 31
rect 4 21 8 29
rect 4 19 5 21
rect 7 19 8 21
rect 4 12 8 19
rect 16 31 22 38
rect 16 29 17 31
rect 19 29 22 31
rect 16 21 22 29
rect 16 19 17 21
rect 19 19 22 21
rect 16 17 22 19
rect 28 31 32 33
rect 28 29 29 31
rect 31 29 32 31
rect 28 21 32 29
rect 28 19 29 21
rect 31 19 32 21
rect 28 12 32 19
rect 38 31 44 38
rect 60 33 64 47
rect 78 43 82 63
rect 68 41 82 43
rect 68 39 69 41
rect 71 39 82 41
rect 68 37 82 39
rect 38 29 41 31
rect 43 29 44 31
rect 38 21 44 29
rect 38 19 41 21
rect 43 19 44 21
rect 38 17 44 19
rect 52 31 56 33
rect 52 29 53 31
rect 55 29 56 31
rect 60 31 68 33
rect 60 29 65 31
rect 67 29 68 31
rect 52 21 56 29
rect 52 19 53 21
rect 55 19 56 21
rect 52 12 56 19
rect 64 21 68 29
rect 64 19 65 21
rect 67 19 68 21
rect 64 17 68 19
rect 76 31 80 33
rect 76 29 77 31
rect 79 29 80 31
rect 76 23 80 29
rect 76 21 77 23
rect 79 21 80 23
rect 76 12 80 21
rect -2 7 92 12
rect -2 5 22 7
rect 24 5 32 7
rect 34 5 92 7
rect -2 0 92 5
<< ptie >>
rect 20 7 36 9
rect 20 5 22 7
rect 24 5 32 7
rect 34 5 36 7
rect 20 3 36 5
<< ntie >>
rect 51 95 57 97
rect 51 93 53 95
rect 55 93 57 95
rect 51 91 57 93
<< nmos >>
rect 11 17 13 35
rect 23 17 25 35
rect 35 17 37 35
rect 47 17 49 35
rect 59 17 61 33
rect 71 17 73 33
<< pmos >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 55 37 94
rect 47 55 49 83
rect 59 55 61 83
rect 71 55 73 91
<< polyct1 >>
rect 29 48 31 50
rect 69 39 71 41
<< ndifct1 >>
rect 5 29 7 31
rect 5 19 7 21
rect 17 29 19 31
rect 17 19 19 21
rect 29 29 31 31
rect 29 19 31 21
rect 41 29 43 31
rect 41 19 43 21
rect 53 29 55 31
rect 53 19 55 21
rect 65 29 67 31
rect 65 19 67 21
rect 77 29 79 31
rect 77 21 79 23
<< ntiect1 >>
rect 53 93 55 95
<< ptiect1 >>
rect 22 5 24 7
rect 32 5 34 7
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 5 69 7 71
rect 17 69 19 71
rect 17 61 19 63
rect 29 89 31 91
rect 29 79 31 81
rect 29 69 31 71
rect 41 69 43 71
rect 41 61 43 63
rect 53 79 55 81
rect 53 69 55 71
rect 65 69 67 71
rect 65 59 67 61
rect 77 79 79 81
rect 77 69 79 71
<< labels >>
rlabel alu1 30 40 30 40 6 z
rlabel alu1 20 45 20 45 6 z
rlabel alu1 30 60 30 60 6 z
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 40 30 40 30 6 z
rlabel alu1 40 65 40 65 6 z
rlabel alu1 45 94 45 94 6 vdd
rlabel alu1 66 25 66 25 6 an
rlabel polyct1 70 40 70 40 6 a
rlabel pdifct1 66 60 66 60 6 an
rlabel alu1 80 50 80 50 6 a
<< end >>
