magic
tech scmos
timestamp 1199203711
<< ab >>
rect 0 0 168 72
<< nwell >>
rect -5 32 173 77
<< pwell >>
rect -5 -5 173 32
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 68 53 70
rect 29 65 31 68
rect 39 65 41 68
rect 51 51 53 68
rect 62 66 64 70
rect 72 66 74 70
rect 82 66 84 70
rect 92 66 94 70
rect 112 66 114 70
rect 122 66 124 70
rect 132 66 134 70
rect 48 49 54 51
rect 48 47 50 49
rect 52 47 54 49
rect 48 45 54 47
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 62 37 64 40
rect 72 37 74 40
rect 143 60 156 62
rect 143 57 145 60
rect 152 58 158 60
rect 152 56 154 58
rect 156 56 158 58
rect 152 54 158 56
rect 153 51 155 54
rect 143 38 145 42
rect 9 33 22 35
rect 29 33 41 35
rect 61 35 74 37
rect 82 35 84 38
rect 92 35 94 38
rect 112 35 114 38
rect 122 35 124 38
rect 61 33 67 35
rect 16 31 18 33
rect 20 31 22 33
rect 16 29 22 31
rect 9 24 11 29
rect 16 27 28 29
rect 16 24 18 27
rect 26 24 28 27
rect 33 24 35 33
rect 61 31 63 33
rect 65 31 67 33
rect 79 33 108 35
rect 79 31 81 33
rect 45 26 47 31
rect 55 29 67 31
rect 55 26 57 29
rect 65 26 67 29
rect 75 29 81 31
rect 102 31 104 33
rect 106 31 108 33
rect 102 29 108 31
rect 112 33 118 35
rect 112 31 114 33
rect 116 31 118 33
rect 112 29 118 31
rect 122 33 128 35
rect 122 31 124 33
rect 126 31 128 33
rect 132 34 134 38
rect 132 32 146 34
rect 122 29 128 31
rect 140 30 142 32
rect 144 30 146 32
rect 75 26 77 29
rect 85 27 91 29
rect 85 25 87 27
rect 89 25 91 27
rect 85 23 97 25
rect 85 20 87 23
rect 95 20 97 23
rect 113 20 115 29
rect 122 25 124 29
rect 140 28 146 30
rect 140 25 142 28
rect 153 26 155 38
rect 120 23 124 25
rect 120 20 122 23
rect 130 20 132 25
rect 9 4 11 12
rect 16 8 18 12
rect 26 8 28 12
rect 33 4 35 12
rect 9 2 35 4
rect 45 4 47 12
rect 55 8 57 12
rect 65 8 67 12
rect 75 4 77 12
rect 45 2 77 4
rect 85 3 87 8
rect 95 3 97 8
rect 140 8 142 12
rect 113 2 115 7
rect 120 2 122 7
rect 130 4 132 7
rect 153 4 155 15
rect 130 2 155 4
<< ndif >>
rect 37 24 45 26
rect 2 16 9 24
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 12 16 24
rect 18 22 26 24
rect 18 20 21 22
rect 23 20 26 22
rect 18 12 26 20
rect 28 12 33 24
rect 35 12 45 24
rect 47 24 55 26
rect 47 22 50 24
rect 52 22 55 24
rect 47 12 55 22
rect 57 17 65 26
rect 57 15 60 17
rect 62 15 65 17
rect 57 12 65 15
rect 67 24 75 26
rect 67 22 70 24
rect 72 22 75 24
rect 67 17 75 22
rect 67 15 70 17
rect 72 15 75 17
rect 67 12 75 15
rect 77 20 82 26
rect 148 25 153 26
rect 135 20 140 25
rect 77 16 85 20
rect 77 14 80 16
rect 82 14 85 16
rect 77 12 85 14
rect 37 7 43 12
rect 37 5 39 7
rect 41 5 43 7
rect 37 3 43 5
rect 80 8 85 12
rect 87 17 95 20
rect 87 15 90 17
rect 92 15 95 17
rect 87 8 95 15
rect 97 10 113 20
rect 97 8 104 10
rect 106 8 113 10
rect 99 7 113 8
rect 115 7 120 20
rect 122 17 130 20
rect 122 15 125 17
rect 127 15 130 17
rect 122 7 130 15
rect 132 18 140 20
rect 132 16 135 18
rect 137 16 140 18
rect 132 12 140 16
rect 142 17 153 25
rect 142 15 147 17
rect 149 15 153 17
rect 155 24 162 26
rect 155 22 158 24
rect 160 22 162 24
rect 155 20 162 22
rect 155 15 160 20
rect 142 12 151 15
rect 132 7 137 12
rect 99 5 111 7
<< pdif >>
rect 4 58 9 65
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 4 38 9 45
rect 11 49 19 65
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 57 29 65
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 42 39 65
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 59 46 65
rect 41 57 49 59
rect 41 55 45 57
rect 47 55 49 57
rect 41 53 49 55
rect 41 38 46 53
rect 55 64 62 66
rect 55 62 57 64
rect 59 62 62 64
rect 55 57 62 62
rect 55 55 57 57
rect 59 55 62 57
rect 55 53 62 55
rect 56 40 62 53
rect 64 56 72 66
rect 64 54 67 56
rect 69 54 72 56
rect 64 49 72 54
rect 64 47 67 49
rect 69 47 72 49
rect 64 40 72 47
rect 74 64 82 66
rect 74 62 77 64
rect 79 62 82 64
rect 74 57 82 62
rect 74 55 77 57
rect 79 55 82 57
rect 74 40 82 55
rect 77 38 82 40
rect 84 42 92 66
rect 84 40 87 42
rect 89 40 92 42
rect 84 38 92 40
rect 94 64 101 66
rect 94 62 97 64
rect 99 62 101 64
rect 94 57 101 62
rect 107 59 112 66
rect 94 55 97 57
rect 99 55 101 57
rect 94 38 101 55
rect 105 57 112 59
rect 105 55 107 57
rect 109 55 112 57
rect 105 53 112 55
rect 107 38 112 53
rect 114 50 122 66
rect 114 48 117 50
rect 119 48 122 50
rect 114 38 122 48
rect 124 49 132 66
rect 124 47 127 49
rect 129 47 132 49
rect 124 42 132 47
rect 124 40 127 42
rect 129 40 132 42
rect 124 38 132 40
rect 134 64 141 66
rect 134 62 137 64
rect 139 62 141 64
rect 134 57 141 62
rect 134 42 143 57
rect 145 51 150 57
rect 145 46 153 51
rect 145 44 148 46
rect 150 44 153 46
rect 145 42 153 44
rect 134 38 141 42
rect 148 38 153 42
rect 155 49 166 51
rect 155 47 162 49
rect 164 47 166 49
rect 155 38 166 47
<< alu1 >>
rect -2 67 170 72
rect -2 65 161 67
rect 163 65 170 67
rect -2 64 170 65
rect 2 57 49 58
rect 2 56 24 57
rect 2 54 4 56
rect 6 55 24 56
rect 26 55 45 57
rect 47 55 49 57
rect 6 54 49 55
rect 146 58 158 59
rect 2 49 6 54
rect 2 47 4 49
rect 2 26 6 47
rect 57 33 87 34
rect 57 31 63 33
rect 65 31 87 33
rect 57 30 87 31
rect 2 22 24 26
rect 20 20 21 22
rect 23 20 24 22
rect 81 22 87 30
rect 20 18 24 20
rect 20 17 64 18
rect 20 15 60 17
rect 62 15 64 17
rect 20 14 64 15
rect 146 56 154 58
rect 156 56 158 58
rect 146 53 158 56
rect 154 45 158 53
rect 145 29 158 35
rect 145 22 151 29
rect -2 7 170 8
rect -2 5 39 7
rect 41 5 160 7
rect 162 5 170 7
rect -2 0 170 5
<< ptie >>
rect 157 7 165 9
rect 157 5 160 7
rect 162 5 165 7
rect 157 3 165 5
<< ntie >>
rect 159 67 165 69
rect 159 65 161 67
rect 163 65 165 67
rect 159 63 165 65
<< nmos >>
rect 9 12 11 24
rect 16 12 18 24
rect 26 12 28 24
rect 33 12 35 24
rect 45 12 47 26
rect 55 12 57 26
rect 65 12 67 26
rect 75 12 77 26
rect 85 8 87 20
rect 95 8 97 20
rect 113 7 115 20
rect 120 7 122 20
rect 130 7 132 20
rect 140 12 142 25
rect 153 15 155 26
<< pmos >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 65
rect 62 40 64 66
rect 72 40 74 66
rect 82 38 84 66
rect 92 38 94 66
rect 112 38 114 66
rect 122 38 124 66
rect 132 38 134 66
rect 143 42 145 57
rect 153 38 155 51
<< polyct0 >>
rect 50 47 52 49
rect 18 31 20 33
rect 104 31 106 33
rect 114 31 116 33
rect 124 31 126 33
rect 142 30 144 32
rect 87 25 89 27
<< polyct1 >>
rect 154 56 156 58
rect 63 31 65 33
<< ndifct0 >>
rect 4 14 6 16
rect 50 22 52 24
rect 70 22 72 24
rect 70 15 72 17
rect 80 14 82 16
rect 90 15 92 17
rect 104 8 106 10
rect 125 15 127 17
rect 135 16 137 18
rect 147 15 149 17
rect 158 22 160 24
<< ndifct1 >>
rect 21 20 23 22
rect 60 15 62 17
rect 39 5 41 7
<< ntiect1 >>
rect 161 65 163 67
<< ptiect1 >>
rect 160 5 162 7
<< pdifct0 >>
rect 14 47 16 49
rect 14 40 16 42
rect 34 40 36 42
rect 57 62 59 64
rect 57 55 59 57
rect 67 54 69 56
rect 67 47 69 49
rect 77 62 79 64
rect 77 55 79 57
rect 87 40 89 42
rect 97 62 99 64
rect 97 55 99 57
rect 107 55 109 57
rect 117 48 119 50
rect 127 47 129 49
rect 127 40 129 42
rect 137 62 139 64
rect 148 44 150 46
rect 162 47 164 49
<< pdifct1 >>
rect 4 54 6 56
rect 4 47 6 49
rect 24 55 26 57
rect 45 55 47 57
<< alu0 >>
rect 55 62 57 64
rect 59 62 61 64
rect 55 57 61 62
rect 75 62 77 64
rect 79 62 81 64
rect 55 55 57 57
rect 59 55 61 57
rect 55 54 61 55
rect 66 56 70 58
rect 66 54 67 56
rect 69 54 70 56
rect 75 57 81 62
rect 75 55 77 57
rect 79 55 81 57
rect 75 54 81 55
rect 95 62 97 64
rect 99 62 101 64
rect 95 57 101 62
rect 135 62 137 64
rect 139 62 141 64
rect 135 61 141 62
rect 95 55 97 57
rect 99 55 101 57
rect 95 54 101 55
rect 105 57 138 58
rect 105 55 107 57
rect 109 55 138 57
rect 105 54 138 55
rect 6 45 7 54
rect 66 50 70 54
rect 115 50 121 51
rect 12 49 99 50
rect 12 47 14 49
rect 16 47 50 49
rect 52 47 67 49
rect 69 47 99 49
rect 12 46 99 47
rect 12 42 17 46
rect 12 40 14 42
rect 16 40 17 42
rect 12 38 17 40
rect 32 42 38 43
rect 85 42 91 43
rect 32 40 34 42
rect 36 40 38 42
rect 32 34 38 40
rect 48 40 87 42
rect 89 40 91 42
rect 48 38 91 40
rect 48 34 52 38
rect 16 33 52 34
rect 16 31 18 33
rect 20 31 52 33
rect 16 30 52 31
rect 48 26 52 30
rect 48 24 73 26
rect 48 22 50 24
rect 52 22 70 24
rect 72 22 73 24
rect 87 27 91 28
rect 89 25 91 27
rect 87 24 91 25
rect 48 21 54 22
rect 3 16 7 18
rect 3 14 4 16
rect 6 14 7 16
rect 69 17 73 22
rect 95 18 99 46
rect 69 15 70 17
rect 72 15 73 17
rect 3 8 7 14
rect 69 13 73 15
rect 79 16 83 18
rect 79 14 80 16
rect 82 14 83 16
rect 88 17 99 18
rect 88 15 90 17
rect 92 15 99 17
rect 88 14 99 15
rect 103 48 117 50
rect 119 48 121 50
rect 103 46 121 48
rect 126 49 130 51
rect 126 47 127 49
rect 129 47 130 49
rect 103 33 107 46
rect 126 42 130 47
rect 103 31 104 33
rect 106 31 107 33
rect 103 18 107 31
rect 113 40 127 42
rect 129 40 130 42
rect 113 38 130 40
rect 134 42 138 54
rect 147 46 151 48
rect 147 44 148 46
rect 150 44 151 46
rect 161 49 165 64
rect 161 47 162 49
rect 164 47 165 49
rect 161 45 165 47
rect 147 42 151 44
rect 134 38 166 42
rect 113 33 117 38
rect 134 34 138 38
rect 113 31 114 33
rect 116 31 117 33
rect 113 26 117 31
rect 122 33 138 34
rect 122 31 124 33
rect 126 31 138 33
rect 122 30 138 31
rect 141 32 145 34
rect 141 30 142 32
rect 144 30 145 32
rect 141 28 145 30
rect 113 22 138 26
rect 162 25 166 38
rect 156 24 166 25
rect 156 22 158 24
rect 160 22 166 24
rect 134 18 138 22
rect 156 21 166 22
rect 103 17 129 18
rect 103 15 125 17
rect 127 15 129 17
rect 103 14 129 15
rect 134 16 135 18
rect 137 16 138 18
rect 134 14 138 16
rect 145 17 151 18
rect 145 15 147 17
rect 149 15 151 17
rect 79 8 83 14
rect 102 10 108 11
rect 102 8 104 10
rect 106 8 108 10
rect 145 8 151 15
<< labels >>
rlabel alu0 35 36 35 36 6 zn
rlabel alu0 14 44 14 44 6 cn
rlabel alu0 71 19 71 19 6 zn
rlabel alu0 60 24 60 24 6 zn
rlabel alu0 68 52 68 52 6 cn
rlabel alu0 93 16 93 16 6 cn
rlabel polyct0 115 32 115 32 6 an
rlabel alu0 88 40 88 40 6 zn
rlabel polyct0 105 32 105 32 6 iz
rlabel alu0 55 48 55 48 6 cn
rlabel alu0 118 48 118 48 6 iz
rlabel alu0 116 16 116 16 6 iz
rlabel alu0 136 20 136 20 6 an
rlabel alu0 130 32 130 32 6 bn
rlabel alu0 161 23 161 23 6 bn
rlabel alu0 149 43 149 43 6 bn
rlabel alu0 128 44 128 44 6 an
rlabel alu0 121 56 121 56 6 bn
rlabel alu1 28 16 28 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 20 24 20 24 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 12 56 12 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 60 16 60 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 68 32 68 32 6 c
rlabel alu1 76 32 76 32 6 c
rlabel alu1 60 32 60 32 6 c
rlabel alu1 44 56 44 56 6 z
rlabel alu1 84 4 84 4 6 vss
rlabel alu1 84 28 84 28 6 c
rlabel alu1 84 68 84 68 6 vdd
rlabel alu1 148 28 148 28 6 a
rlabel alu1 156 32 156 32 6 a
rlabel alu1 156 52 156 52 6 b
rlabel alu1 148 56 148 56 6 b
<< end >>
