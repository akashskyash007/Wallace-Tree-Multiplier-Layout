magic
tech scmos
timestamp 1199469067
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 11 83 13 88
rect 23 83 25 88
rect 35 83 37 88
rect 47 83 49 88
rect 11 38 13 63
rect 23 48 25 63
rect 35 58 37 63
rect 35 56 43 58
rect 35 55 39 56
rect 37 54 39 55
rect 41 54 43 56
rect 37 52 43 54
rect 23 46 33 48
rect 23 45 29 46
rect 25 44 29 45
rect 31 44 33 46
rect 25 42 33 44
rect 11 36 21 38
rect 15 34 17 36
rect 19 34 21 36
rect 15 32 21 34
rect 17 26 19 32
rect 25 26 27 42
rect 37 26 39 52
rect 47 38 49 63
rect 47 36 53 38
rect 47 35 49 36
rect 45 34 49 35
rect 51 34 53 36
rect 45 32 53 34
rect 45 26 47 32
rect 17 12 19 17
rect 25 12 27 17
rect 37 12 39 17
rect 45 12 47 17
<< ndif >>
rect 9 17 17 26
rect 19 17 25 26
rect 27 21 37 26
rect 27 19 31 21
rect 33 19 37 21
rect 27 17 37 19
rect 39 17 45 26
rect 47 21 56 26
rect 47 19 51 21
rect 53 19 56 21
rect 47 17 56 19
rect 9 11 15 17
rect 9 9 11 11
rect 13 9 15 11
rect 9 7 15 9
<< pdif >>
rect 3 81 11 83
rect 3 79 5 81
rect 7 79 11 81
rect 3 77 11 79
rect 6 63 11 77
rect 13 71 23 83
rect 13 69 17 71
rect 19 69 23 71
rect 13 63 23 69
rect 25 81 35 83
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 63 35 69
rect 37 81 47 83
rect 37 79 41 81
rect 43 79 47 81
rect 37 63 47 79
rect 49 81 57 83
rect 49 79 53 81
rect 55 79 57 81
rect 49 73 57 79
rect 49 71 53 73
rect 55 71 57 73
rect 49 69 57 71
rect 49 63 54 69
<< alu1 >>
rect -2 95 62 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 62 95
rect -2 88 62 93
rect 3 81 33 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 79 33 81
rect 3 78 33 79
rect 8 71 23 73
rect 8 69 17 71
rect 19 69 23 71
rect 8 68 23 69
rect 27 72 33 78
rect 40 81 44 88
rect 40 79 41 81
rect 43 79 44 81
rect 40 77 44 79
rect 52 81 56 83
rect 52 79 53 81
rect 55 79 56 81
rect 52 73 56 79
rect 52 72 53 73
rect 27 71 53 72
rect 55 71 56 73
rect 27 69 29 71
rect 31 69 56 71
rect 27 68 56 69
rect 8 23 12 68
rect 17 58 32 63
rect 18 38 22 53
rect 16 36 22 38
rect 28 46 32 58
rect 28 44 29 46
rect 31 44 32 46
rect 28 37 32 44
rect 38 58 53 63
rect 38 56 42 58
rect 38 54 39 56
rect 41 54 42 56
rect 38 37 42 54
rect 16 34 17 36
rect 19 34 22 36
rect 16 32 22 34
rect 48 36 52 43
rect 48 34 49 36
rect 51 34 52 36
rect 48 33 52 34
rect 18 27 33 32
rect 38 27 52 33
rect 8 21 34 23
rect 8 19 31 21
rect 33 19 34 21
rect 8 17 34 19
rect 38 17 42 27
rect 50 21 54 23
rect 50 19 51 21
rect 53 19 54 21
rect 50 12 54 19
rect -2 11 62 12
rect -2 9 11 11
rect 13 9 62 11
rect -2 7 62 9
rect -2 5 39 7
rect 41 5 49 7
rect 51 5 62 7
rect -2 0 62 5
<< ptie >>
rect 37 7 53 9
rect 37 5 39 7
rect 41 5 49 7
rect 51 5 53 7
rect 37 3 53 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 17 17 19 26
rect 25 17 27 26
rect 37 17 39 26
rect 45 17 47 26
<< pmos >>
rect 11 63 13 83
rect 23 63 25 83
rect 35 63 37 83
rect 47 63 49 83
<< polyct1 >>
rect 39 54 41 56
rect 29 44 31 46
rect 17 34 19 36
rect 49 34 51 36
<< ndifct1 >>
rect 31 19 33 21
rect 51 19 53 21
rect 11 9 13 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 39 5 41 7
rect 49 5 51 7
<< pdifct1 >>
rect 5 79 7 81
rect 17 69 19 71
rect 29 79 31 81
rect 29 69 31 71
rect 41 79 43 81
rect 53 79 55 81
rect 53 71 55 73
<< labels >>
rlabel pdifct1 6 80 6 80 6 n3
rlabel pdifct1 30 80 30 80 6 n3
rlabel pdifct1 30 70 30 70 6 n3
rlabel pdifct1 54 72 54 72 6 n3
rlabel pdifct1 54 80 54 80 6 n3
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 40 20 40 6 b1
rlabel alu1 20 70 20 70 6 z
rlabel alu1 20 60 20 60 6 b2
rlabel alu1 30 20 30 20 6 z
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 40 25 40 25 6 a1
rlabel alu1 30 30 30 30 6 b1
rlabel alu1 40 50 40 50 6 a2
rlabel alu1 30 50 30 50 6 b2
rlabel alu1 30 94 30 94 6 vdd
rlabel polyct1 50 35 50 35 6 a1
rlabel alu1 50 60 50 60 6 a2
<< end >>
