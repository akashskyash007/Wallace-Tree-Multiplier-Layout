magic
tech scmos
timestamp 1199203597
<< ab >>
rect 0 0 160 72
<< nwell >>
rect -5 32 165 77
<< pwell >>
rect -5 -5 165 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 71 68
rect 49 63 51 66
rect 59 63 61 66
rect 69 63 71 66
rect 79 63 81 68
rect 89 63 91 68
rect 119 63 121 68
rect 129 63 131 68
rect 139 63 141 68
rect 149 63 151 68
rect 99 57 101 61
rect 109 57 111 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 33 41 35
rect 49 34 51 38
rect 59 34 61 38
rect 69 35 71 38
rect 79 35 81 38
rect 89 35 91 38
rect 99 35 101 38
rect 109 35 111 38
rect 119 35 121 38
rect 129 35 131 38
rect 139 35 141 38
rect 149 35 151 38
rect 66 33 72 35
rect 9 31 11 33
rect 13 31 32 33
rect 9 29 32 31
rect 66 31 68 33
rect 70 31 72 33
rect 20 26 22 29
rect 30 26 32 29
rect 50 26 52 30
rect 60 26 62 30
rect 66 29 72 31
rect 70 26 72 29
rect 77 33 94 35
rect 77 31 79 33
rect 81 31 86 33
rect 88 31 94 33
rect 77 29 94 31
rect 77 26 79 29
rect 92 26 94 29
rect 99 33 111 35
rect 99 31 101 33
rect 103 31 111 33
rect 99 29 111 31
rect 115 33 121 35
rect 115 31 117 33
rect 119 31 121 33
rect 115 29 121 31
rect 128 33 151 35
rect 128 31 147 33
rect 149 31 151 33
rect 128 29 151 31
rect 99 26 101 29
rect 109 26 111 29
rect 116 26 118 29
rect 128 26 130 29
rect 138 26 140 29
rect 20 2 22 7
rect 30 4 32 7
rect 50 4 52 7
rect 60 4 62 7
rect 30 2 62 4
rect 70 2 72 6
rect 77 2 79 6
rect 92 4 94 12
rect 99 8 101 12
rect 109 8 111 12
rect 116 4 118 12
rect 92 2 118 4
rect 128 2 130 7
rect 138 2 140 7
<< ndif >>
rect 13 19 20 26
rect 13 17 15 19
rect 17 17 20 19
rect 13 11 20 17
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
rect 22 24 30 26
rect 22 22 25 24
rect 27 22 30 24
rect 22 17 30 22
rect 22 15 25 17
rect 27 15 30 17
rect 22 7 30 15
rect 32 19 39 26
rect 45 19 50 26
rect 32 17 35 19
rect 37 17 39 19
rect 32 11 39 17
rect 43 17 50 19
rect 43 15 45 17
rect 47 15 50 17
rect 43 13 50 15
rect 32 9 35 11
rect 37 9 39 11
rect 32 7 39 9
rect 45 7 50 13
rect 52 24 60 26
rect 52 22 55 24
rect 57 22 60 24
rect 52 7 60 22
rect 62 17 70 26
rect 62 15 65 17
rect 67 15 70 17
rect 62 7 70 15
rect 65 6 70 7
rect 72 6 77 26
rect 79 12 92 26
rect 94 12 99 26
rect 101 17 109 26
rect 101 15 104 17
rect 106 15 109 17
rect 101 12 109 15
rect 111 12 116 26
rect 118 16 128 26
rect 118 14 121 16
rect 123 14 128 16
rect 118 12 128 14
rect 79 7 90 12
rect 79 6 84 7
rect 81 5 84 6
rect 86 5 90 7
rect 81 3 90 5
rect 120 7 128 12
rect 130 24 138 26
rect 130 22 133 24
rect 135 22 138 24
rect 130 17 138 22
rect 130 15 133 17
rect 135 15 138 17
rect 130 7 138 15
rect 140 19 147 26
rect 140 17 143 19
rect 145 17 147 19
rect 140 11 147 17
rect 140 9 143 11
rect 145 9 147 11
rect 140 7 147 9
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 19 66
rect 11 62 14 64
rect 16 62 19 64
rect 11 57 19 62
rect 11 55 14 57
rect 16 55 19 57
rect 11 38 19 55
rect 21 49 29 66
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 64 39 66
rect 31 62 34 64
rect 36 62 39 64
rect 31 57 39 62
rect 31 55 34 57
rect 36 55 39 57
rect 31 38 39 55
rect 41 63 46 66
rect 41 56 49 63
rect 41 54 44 56
rect 46 54 49 56
rect 41 49 49 54
rect 41 47 44 49
rect 46 47 49 49
rect 41 38 49 47
rect 51 58 59 63
rect 51 56 54 58
rect 56 56 59 58
rect 51 42 59 56
rect 51 40 54 42
rect 56 40 59 42
rect 51 38 59 40
rect 61 49 69 63
rect 61 47 64 49
rect 66 47 69 49
rect 61 42 69 47
rect 61 40 64 42
rect 66 40 69 42
rect 61 38 69 40
rect 71 58 79 63
rect 71 56 74 58
rect 76 56 79 58
rect 71 51 79 56
rect 71 49 74 51
rect 76 49 79 51
rect 71 38 79 49
rect 81 49 89 63
rect 81 47 84 49
rect 86 47 89 49
rect 81 42 89 47
rect 81 40 84 42
rect 86 40 89 42
rect 81 38 89 40
rect 91 57 96 63
rect 114 57 119 63
rect 91 51 99 57
rect 91 49 94 51
rect 96 49 99 51
rect 91 38 99 49
rect 101 42 109 57
rect 101 40 104 42
rect 106 40 109 42
rect 101 38 109 40
rect 111 50 119 57
rect 111 48 114 50
rect 116 48 119 50
rect 111 38 119 48
rect 121 49 129 63
rect 121 47 124 49
rect 126 47 129 49
rect 121 42 129 47
rect 121 40 124 42
rect 126 40 129 42
rect 121 38 129 40
rect 131 61 139 63
rect 131 59 134 61
rect 136 59 139 61
rect 131 53 139 59
rect 131 51 134 53
rect 136 51 139 53
rect 131 38 139 51
rect 141 49 149 63
rect 141 47 144 49
rect 146 47 149 49
rect 141 42 149 47
rect 141 40 144 42
rect 146 40 149 42
rect 141 38 149 40
rect 151 61 158 63
rect 151 59 154 61
rect 156 59 158 61
rect 151 53 158 59
rect 151 51 154 53
rect 156 51 158 53
rect 151 38 158 51
<< alu1 >>
rect -2 67 162 72
rect -2 65 104 67
rect 106 65 162 67
rect -2 64 162 65
rect 52 42 58 43
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 2 21 6 29
rect 42 40 54 42
rect 56 40 58 42
rect 42 38 58 40
rect 42 18 46 38
rect 154 34 158 43
rect 145 33 158 34
rect 145 31 147 33
rect 149 31 158 33
rect 145 29 158 31
rect 42 17 108 18
rect 42 15 45 17
rect 47 15 65 17
rect 67 15 104 17
rect 106 15 108 17
rect 42 14 108 15
rect -2 7 162 8
rect -2 5 5 7
rect 7 5 84 7
rect 86 5 153 7
rect 155 5 162 7
rect -2 0 162 5
<< ptie >>
rect 3 7 9 24
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 151 7 157 24
rect 151 5 153 7
rect 155 5 157 7
rect 151 3 157 5
<< ntie >>
rect 100 67 110 69
rect 100 65 104 67
rect 106 65 110 67
rect 100 63 110 65
<< nmos >>
rect 20 7 22 26
rect 30 7 32 26
rect 50 7 52 26
rect 60 7 62 26
rect 70 6 72 26
rect 77 6 79 26
rect 92 12 94 26
rect 99 12 101 26
rect 109 12 111 26
rect 116 12 118 26
rect 128 7 130 26
rect 138 7 140 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 63
rect 59 38 61 63
rect 69 38 71 63
rect 79 38 81 63
rect 89 38 91 63
rect 99 38 101 57
rect 109 38 111 57
rect 119 38 121 63
rect 129 38 131 63
rect 139 38 141 63
rect 149 38 151 63
<< polyct0 >>
rect 68 31 70 33
rect 79 31 81 33
rect 86 31 88 33
rect 101 31 103 33
rect 117 31 119 33
<< polyct1 >>
rect 11 31 13 33
rect 147 31 149 33
<< ndifct0 >>
rect 15 17 17 19
rect 15 9 17 11
rect 25 22 27 24
rect 25 15 27 17
rect 35 17 37 19
rect 35 9 37 11
rect 55 22 57 24
rect 121 14 123 16
rect 133 22 135 24
rect 133 15 135 17
rect 143 17 145 19
rect 143 9 145 11
<< ndifct1 >>
rect 45 15 47 17
rect 65 15 67 17
rect 104 15 106 17
rect 84 5 86 7
<< ntiect1 >>
rect 104 65 106 67
<< ptiect1 >>
rect 5 5 7 7
rect 153 5 155 7
<< pdifct0 >>
rect 4 47 6 49
rect 4 40 6 42
rect 14 62 16 64
rect 14 55 16 57
rect 24 47 26 49
rect 24 40 26 42
rect 34 62 36 64
rect 34 55 36 57
rect 44 54 46 56
rect 44 47 46 49
rect 54 56 56 58
rect 64 47 66 49
rect 64 40 66 42
rect 74 56 76 58
rect 74 49 76 51
rect 84 47 86 49
rect 84 40 86 42
rect 94 49 96 51
rect 104 40 106 42
rect 114 48 116 50
rect 124 47 126 49
rect 124 40 126 42
rect 134 59 136 61
rect 134 51 136 53
rect 144 47 146 49
rect 144 40 146 42
rect 154 59 156 61
rect 154 51 156 53
<< pdifct1 >>
rect 54 40 56 42
<< alu0 >>
rect 12 62 14 64
rect 16 62 18 64
rect 12 57 18 62
rect 12 55 14 57
rect 16 55 18 57
rect 12 54 18 55
rect 32 62 34 64
rect 36 62 38 64
rect 32 57 38 62
rect 133 61 137 64
rect 133 59 134 61
rect 136 59 137 61
rect 52 58 97 59
rect 32 55 34 57
rect 36 55 38 57
rect 32 54 38 55
rect 43 56 47 58
rect 43 54 44 56
rect 46 54 47 56
rect 52 56 54 58
rect 56 56 74 58
rect 76 56 97 58
rect 52 55 97 56
rect 43 50 47 54
rect 73 51 77 55
rect 93 51 97 55
rect 133 53 137 59
rect 133 51 134 53
rect 136 51 137 53
rect 153 61 157 64
rect 153 59 154 61
rect 156 59 157 61
rect 153 53 157 59
rect 153 51 154 53
rect 156 51 157 53
rect 2 49 68 50
rect 2 47 4 49
rect 6 47 24 49
rect 26 47 44 49
rect 46 47 64 49
rect 66 47 68 49
rect 73 49 74 51
rect 76 49 77 51
rect 73 47 77 49
rect 82 49 87 51
rect 82 47 84 49
rect 86 47 87 49
rect 93 49 94 51
rect 96 50 118 51
rect 96 49 114 50
rect 93 48 114 49
rect 116 48 118 50
rect 93 47 118 48
rect 123 49 127 51
rect 133 49 137 51
rect 143 49 147 51
rect 153 49 157 51
rect 123 47 124 49
rect 126 47 127 49
rect 2 46 68 47
rect 2 42 7 46
rect 2 40 4 42
rect 6 40 7 42
rect 2 38 7 40
rect 23 42 28 46
rect 62 43 68 46
rect 82 43 87 47
rect 23 40 24 42
rect 26 40 28 42
rect 23 38 28 40
rect 24 24 28 38
rect 24 22 25 24
rect 27 22 28 24
rect 14 19 18 21
rect 14 17 15 19
rect 17 17 18 19
rect 14 11 18 17
rect 24 17 28 22
rect 62 42 78 43
rect 62 40 64 42
rect 66 40 78 42
rect 62 39 78 40
rect 82 42 98 43
rect 82 40 84 42
rect 86 40 98 42
rect 82 39 98 40
rect 102 42 117 43
rect 102 40 104 42
rect 106 40 117 42
rect 102 39 117 40
rect 24 15 25 17
rect 27 15 28 17
rect 24 13 28 15
rect 34 19 38 21
rect 34 17 35 19
rect 37 17 38 19
rect 14 9 15 11
rect 17 9 18 11
rect 14 8 18 9
rect 34 11 38 17
rect 67 33 71 35
rect 67 31 68 33
rect 70 31 71 33
rect 67 26 71 31
rect 74 34 78 39
rect 94 34 98 39
rect 113 34 117 39
rect 123 42 127 47
rect 143 47 144 49
rect 146 47 147 49
rect 143 42 147 47
rect 123 40 124 42
rect 126 40 144 42
rect 146 40 147 42
rect 123 38 147 40
rect 74 33 90 34
rect 74 31 79 33
rect 81 31 86 33
rect 88 31 90 33
rect 74 30 90 31
rect 94 33 105 34
rect 94 31 101 33
rect 103 31 105 33
rect 94 30 105 31
rect 113 33 121 34
rect 113 31 117 33
rect 119 31 121 33
rect 113 30 121 31
rect 94 26 98 30
rect 132 26 136 38
rect 53 24 136 26
rect 53 22 55 24
rect 57 22 133 24
rect 135 22 136 24
rect 53 21 59 22
rect 120 16 124 18
rect 120 14 121 16
rect 123 14 124 16
rect 34 9 35 11
rect 37 9 38 11
rect 34 8 38 9
rect 120 8 124 14
rect 132 17 136 22
rect 132 15 133 17
rect 135 15 136 17
rect 132 13 136 15
rect 142 19 146 21
rect 142 17 143 19
rect 145 17 146 19
rect 142 11 146 17
rect 142 9 143 11
rect 145 9 146 11
rect 142 8 146 9
<< labels >>
rlabel alu0 4 44 4 44 6 bn
rlabel alu0 26 31 26 31 6 bn
rlabel alu0 69 28 69 28 6 an
rlabel alu0 35 48 35 48 6 bn
rlabel alu0 65 44 65 44 6 bn
rlabel alu0 70 41 70 41 6 bn
rlabel alu0 45 52 45 52 6 bn
rlabel alu0 82 32 82 32 6 bn
rlabel alu0 99 32 99 32 6 an
rlabel alu0 115 36 115 36 6 bn
rlabel alu0 84 45 84 45 6 an
rlabel alu0 109 41 109 41 6 bn
rlabel alu0 94 24 94 24 6 an
rlabel alu0 125 44 125 44 6 an
rlabel alu0 145 44 145 44 6 an
rlabel alu0 134 27 134 27 6 an
rlabel alu1 4 28 4 28 6 b
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 52 16 52 16 6 z
rlabel alu1 60 16 60 16 6 z
rlabel alu1 68 16 68 16 6 z
rlabel alu1 76 16 76 16 6 z
rlabel alu1 44 28 44 28 6 z
rlabel alu1 52 40 52 40 6 z
rlabel alu1 80 4 80 4 6 vss
rlabel alu1 100 16 100 16 6 z
rlabel alu1 92 16 92 16 6 z
rlabel alu1 84 16 84 16 6 z
rlabel alu1 80 68 80 68 6 vdd
rlabel polyct1 148 32 148 32 6 a
rlabel alu1 156 36 156 36 6 a
<< end >>
