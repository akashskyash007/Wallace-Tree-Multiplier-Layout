magic
tech scmos
timestamp 1199202294
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 21 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 9 30 11 33
rect 19 30 21 33
rect 9 6 11 11
rect 19 6 21 11
<< ndif >>
rect 2 22 9 30
rect 2 20 4 22
rect 6 20 9 22
rect 2 15 9 20
rect 2 13 4 15
rect 6 13 9 15
rect 2 11 9 13
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 11 19 19
rect 21 22 29 30
rect 21 20 24 22
rect 26 20 29 22
rect 21 15 29 20
rect 21 13 24 15
rect 26 13 29 15
rect 21 11 29 13
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 30 6 50
rect 26 38 30 47
rect 15 37 30 38
rect 15 35 17 37
rect 19 35 30 37
rect 15 34 30 35
rect 2 28 23 30
rect 2 26 14 28
rect 16 26 23 28
rect 13 21 17 26
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 11 11 30
rect 19 11 21 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
<< polyct1 >>
rect 17 35 19 37
<< ndifct0 >>
rect 4 20 6 22
rect 4 13 6 15
rect 24 20 26 22
rect 24 13 26 15
<< ndifct1 >>
rect 14 26 16 28
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 66 26 68
rect 24 59 26 61
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 61 28 66
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 2 22 8 23
rect 2 20 4 22
rect 6 20 8 22
rect 2 15 8 20
rect 22 22 28 23
rect 22 20 24 22
rect 26 20 28 22
rect 2 13 4 15
rect 6 13 8 15
rect 2 12 8 13
rect 22 15 28 20
rect 22 13 24 15
rect 26 13 28 15
rect 22 12 28 13
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 20 28 20 28 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 44 28 44 6 a
<< end >>
