magic
tech scmos
timestamp 1199202784
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 9 39 11 50
rect 19 47 21 50
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 19 41 25 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 36 15 37
rect 13 35 16 36
rect 9 33 16 35
rect 14 30 16 33
rect 21 30 23 41
rect 29 39 31 50
rect 39 39 41 50
rect 49 47 51 50
rect 29 37 41 39
rect 29 36 33 37
rect 28 35 33 36
rect 35 35 41 37
rect 28 33 41 35
rect 45 45 51 47
rect 45 43 47 45
rect 49 43 51 45
rect 45 41 51 43
rect 28 30 30 33
rect 38 30 40 33
rect 45 30 47 41
rect 59 39 61 50
rect 55 37 61 39
rect 55 36 57 37
rect 52 35 57 36
rect 59 35 61 37
rect 52 33 61 35
rect 52 30 54 33
rect 14 6 16 10
rect 21 6 23 10
rect 28 6 30 10
rect 38 6 40 10
rect 45 6 47 10
rect 52 6 54 10
<< ndif >>
rect 6 14 14 30
rect 6 12 9 14
rect 11 12 14 14
rect 6 10 14 12
rect 16 10 21 30
rect 23 10 28 30
rect 30 21 38 30
rect 30 19 33 21
rect 35 19 38 21
rect 30 10 38 19
rect 40 10 45 30
rect 47 10 52 30
rect 54 28 62 30
rect 54 26 57 28
rect 59 26 62 28
rect 54 21 62 26
rect 54 19 57 21
rect 59 19 62 21
rect 54 17 62 19
rect 54 10 59 17
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 50 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 50 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 50 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 50 39 52
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 50 49 66
rect 51 61 59 70
rect 51 59 54 61
rect 56 59 59 61
rect 51 54 59 59
rect 51 52 54 54
rect 56 52 59 54
rect 51 50 59 52
rect 61 68 68 70
rect 61 66 64 68
rect 66 66 68 68
rect 61 61 68 66
rect 61 59 64 61
rect 66 59 68 61
rect 61 50 68 59
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 32 61 58 62
rect 32 59 34 61
rect 36 59 54 61
rect 56 59 58 61
rect 32 58 58 59
rect 32 54 37 58
rect 53 54 58 58
rect 2 52 14 54
rect 16 52 34 54
rect 36 52 37 54
rect 2 50 37 52
rect 2 22 6 50
rect 41 46 47 54
rect 53 52 54 54
rect 56 52 63 54
rect 53 50 63 52
rect 19 45 55 46
rect 19 43 21 45
rect 23 43 47 45
rect 49 43 55 45
rect 19 42 55 43
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 25 37 39 38
rect 25 35 33 37
rect 35 35 39 37
rect 25 34 39 35
rect 44 37 63 38
rect 44 35 57 37
rect 59 35 63 37
rect 44 34 63 35
rect 44 30 48 34
rect 10 26 48 30
rect 2 21 37 22
rect 2 19 33 21
rect 35 19 37 21
rect 2 18 37 19
rect 42 17 46 26
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 14 10 16 30
rect 21 10 23 30
rect 28 10 30 30
rect 38 10 40 30
rect 45 10 47 30
rect 52 10 54 30
<< pmos >>
rect 9 50 11 70
rect 19 50 21 70
rect 29 50 31 70
rect 39 50 41 70
rect 49 50 51 70
rect 59 50 61 70
<< polyct1 >>
rect 21 43 23 45
rect 11 35 13 37
rect 33 35 35 37
rect 47 43 49 45
rect 57 35 59 37
<< ndifct0 >>
rect 9 12 11 14
rect 57 26 59 28
rect 57 19 59 21
<< ndifct1 >>
rect 33 19 35 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 59 16 61
rect 24 66 26 68
rect 24 59 26 61
rect 44 66 46 68
rect 64 66 66 68
rect 64 59 66 61
<< pdifct1 >>
rect 14 52 16 54
rect 34 59 36 61
rect 34 52 36 54
rect 54 59 56 61
rect 54 52 56 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 61 28 66
rect 42 66 44 68
rect 46 66 48 68
rect 42 65 48 66
rect 62 66 64 68
rect 66 66 68 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 62 61 68 66
rect 62 59 64 61
rect 66 59 68 61
rect 62 58 68 59
rect 55 28 61 29
rect 55 26 57 28
rect 59 26 61 28
rect 55 21 61 26
rect 55 19 57 21
rect 59 19 61 21
rect 7 14 13 15
rect 7 12 9 14
rect 11 12 13 14
rect 55 12 61 19
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 28 36 28 36 6 c
rlabel alu1 28 44 28 44 6 b
rlabel alu1 36 36 36 36 6 c
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 44 24 44 24 6 a
rlabel alu1 52 36 52 36 6 a
rlabel alu1 52 44 52 44 6 b
rlabel alu1 44 48 44 48 6 b
rlabel alu1 44 60 44 60 6 z
rlabel alu1 52 60 52 60 6 z
rlabel alu1 60 36 60 36 6 a
rlabel alu1 60 52 60 52 6 z
<< end >>
