magic
tech scmos
timestamp 1199202570
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 9 39 11 46
rect 19 39 21 46
rect 29 39 31 46
rect 39 39 41 46
rect 49 40 51 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 19 33 31 35
rect 35 37 41 39
rect 35 35 37 37
rect 39 35 41 37
rect 35 33 41 35
rect 45 38 51 40
rect 45 36 47 38
rect 49 36 51 38
rect 45 34 51 36
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 30 38 33
rect 47 30 49 34
rect 47 11 49 16
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
<< ndif >>
rect 4 14 12 30
rect 4 12 7 14
rect 9 12 12 14
rect 4 10 12 12
rect 14 10 19 30
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 10 29 19
rect 31 10 36 30
rect 38 21 47 30
rect 38 19 41 21
rect 43 19 47 21
rect 38 16 47 19
rect 49 28 56 30
rect 49 26 52 28
rect 54 26 56 28
rect 49 21 56 26
rect 49 19 52 21
rect 54 19 56 21
rect 49 16 56 19
rect 38 14 45 16
rect 38 12 41 14
rect 43 12 45 14
rect 38 10 45 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 46 9 59
rect 11 60 19 70
rect 11 58 14 60
rect 16 58 19 60
rect 11 53 19 58
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 46 29 59
rect 31 60 39 70
rect 31 58 34 60
rect 36 58 39 60
rect 31 53 39 58
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 61 49 66
rect 41 59 44 61
rect 46 59 49 61
rect 41 46 49 59
rect 43 43 49 46
rect 51 56 56 70
rect 51 54 58 56
rect 51 52 54 54
rect 56 52 58 54
rect 51 47 58 52
rect 51 45 54 47
rect 56 45 58 47
rect 51 43 58 45
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 33 60 38 63
rect 33 58 34 60
rect 36 58 38 60
rect 33 54 38 58
rect 2 53 38 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 51 38 53
rect 2 50 38 51
rect 2 22 6 50
rect 42 46 46 55
rect 17 38 23 46
rect 33 42 50 46
rect 46 38 50 42
rect 17 37 31 38
rect 17 35 27 37
rect 29 35 31 37
rect 17 34 31 35
rect 46 36 47 38
rect 49 36 50 38
rect 46 34 50 36
rect 2 21 31 22
rect 2 19 24 21
rect 26 19 31 21
rect 2 18 31 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 47 16 49 30
<< pmos >>
rect 9 46 11 70
rect 19 46 21 70
rect 29 46 31 70
rect 39 46 41 70
rect 49 43 51 70
<< polyct0 >>
rect 11 35 13 37
rect 37 35 39 37
<< polyct1 >>
rect 27 35 29 37
rect 47 36 49 38
<< ndifct0 >>
rect 7 12 9 14
rect 41 19 43 21
rect 52 26 54 28
rect 52 19 54 21
rect 41 12 43 14
<< ndifct1 >>
rect 24 19 26 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 58 16 60
rect 24 66 26 68
rect 24 59 26 61
rect 44 66 46 68
rect 44 59 46 61
rect 54 52 56 54
rect 54 45 56 47
<< pdifct1 >>
rect 14 51 16 53
rect 34 58 36 60
rect 34 51 36 53
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 60 17 62
rect 13 58 14 60
rect 16 58 17 60
rect 22 61 28 66
rect 42 66 44 68
rect 46 66 48 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 42 61 48 66
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 13 54 17 58
rect 53 54 57 56
rect 53 52 54 54
rect 56 52 57 54
rect 53 47 57 52
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 35 37 41 38
rect 35 35 37 37
rect 39 35 41 37
rect 35 30 41 35
rect 53 45 54 47
rect 56 45 57 47
rect 53 30 57 45
rect 10 28 57 30
rect 10 26 52 28
rect 54 26 57 28
rect 39 21 45 22
rect 39 19 41 21
rect 43 19 45 21
rect 5 14 11 15
rect 5 12 7 14
rect 9 12 11 14
rect 39 14 45 19
rect 51 21 55 26
rect 51 19 52 21
rect 54 19 55 21
rect 51 17 55 19
rect 39 12 41 14
rect 43 12 45 14
<< labels >>
rlabel alu0 12 32 12 32 6 an
rlabel alu0 38 32 38 32 6 an
rlabel alu0 53 23 53 23 6 an
rlabel alu0 55 41 55 41 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel polyct1 28 36 28 36 6 b
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 44 36 44 6 a
rlabel alu1 44 48 44 48 6 a
rlabel alu1 36 60 36 60 6 z
rlabel alu1 32 74 32 74 6 vdd
<< end >>
