magic
tech scmos
timestamp 1199973035
<< ab >>
rect 0 0 32 88
<< nwell >>
rect -5 40 37 97
<< pwell >>
rect -5 -9 37 40
<< poly >>
rect 2 81 11 83
rect 2 79 7 81
rect 9 79 11 81
rect 2 77 11 79
rect 9 74 11 77
rect 21 81 30 83
rect 21 79 24 81
rect 26 79 30 81
rect 21 77 30 79
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 37 14 43
rect 18 37 30 43
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndif >>
rect 2 14 9 34
rect 11 25 21 34
rect 11 23 15 25
rect 17 23 21 25
rect 11 18 21 23
rect 11 16 15 18
rect 17 16 21 18
rect 11 14 21 16
rect 23 29 30 34
rect 23 27 26 29
rect 28 27 30 29
rect 23 21 30 27
rect 23 19 26 21
rect 28 19 30 21
rect 23 14 30 19
rect 13 2 19 14
<< pdif >>
rect 13 81 19 86
rect 13 79 15 81
rect 17 79 19 81
rect 13 74 19 79
rect 2 46 9 74
rect 11 72 15 74
rect 17 72 21 74
rect 11 46 21 72
rect 23 53 30 74
rect 23 51 26 53
rect 28 51 30 53
rect 23 46 30 51
<< alu1 >>
rect -2 89 34 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 34 89
rect -2 86 34 87
rect 14 81 18 82
rect 14 79 15 81
rect 17 79 18 81
rect 14 78 18 79
rect 22 81 28 82
rect 22 79 24 81
rect 26 79 28 81
rect 22 66 28 79
rect 14 62 28 66
rect 14 41 18 62
rect 22 53 30 55
rect 22 51 26 53
rect 28 51 30 53
rect 22 50 30 51
rect 22 30 26 50
rect 22 29 29 30
rect 22 27 26 29
rect 28 27 29 29
rect 22 21 29 27
rect 22 19 26 21
rect 28 19 29 21
rect 22 17 29 19
rect 14 9 18 10
rect 14 7 15 9
rect 17 7 18 9
rect 14 6 18 7
rect -2 1 34 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< alu2 >>
rect -2 89 34 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 34 89
rect -2 81 34 87
rect -2 79 15 81
rect 17 79 34 81
rect -2 76 34 79
rect -2 9 34 12
rect -2 7 15 9
rect 17 7 34 9
rect -2 1 34 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 32 3
rect 25 -1 27 1
rect 29 -1 32 1
rect 25 -3 32 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 32 91
rect 25 87 27 89
rect 29 87 32 89
rect 25 85 32 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
<< polyct0 >>
rect 7 79 9 81
<< polyct1 >>
rect 24 79 26 81
<< ndifct0 >>
rect 15 23 17 25
rect 15 16 17 18
<< ndifct1 >>
rect 26 27 28 29
rect 26 19 28 21
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
<< pdifct0 >>
rect 15 72 17 74
<< pdifct1 >>
rect 15 79 17 81
rect 26 51 28 53
<< alu0 >>
rect 6 81 10 86
rect 6 79 7 81
rect 9 79 10 81
rect 6 77 10 79
rect 14 82 18 86
rect 14 74 18 78
rect 14 72 15 74
rect 17 72 18 74
rect 14 70 18 72
rect 14 25 18 27
rect 14 23 15 25
rect 17 23 18 25
rect 14 18 18 23
rect 14 16 15 18
rect 17 16 18 18
rect 14 10 18 16
rect 14 2 18 6
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 15 79 17 81
rect 15 7 17 9
rect 7 -1 9 1
rect 23 -1 25 1
<< labels >>
rlabel alu1 16 52 16 52 6 a
rlabel alu1 24 36 24 36 6 z
rlabel alu1 24 68 24 68 6 a
rlabel alu2 16 6 16 6 6 vss
rlabel alu2 16 6 16 6 6 vss
rlabel alu2 16 82 16 82 6 vdd
<< end >>
