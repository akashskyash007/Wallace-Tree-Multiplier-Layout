magic
tech scmos
timestamp 1199201708
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 62 11 67
rect 19 61 21 65
rect 29 61 31 65
rect 41 62 43 66
rect 9 40 11 50
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 19 39 21 50
rect 29 47 31 50
rect 29 45 37 47
rect 29 44 33 45
rect 31 43 33 44
rect 35 43 37 45
rect 31 41 37 43
rect 19 37 26 39
rect 19 35 21 37
rect 23 35 26 37
rect 9 30 11 34
rect 19 33 26 35
rect 24 30 26 33
rect 31 30 33 41
rect 41 39 43 51
rect 41 37 47 39
rect 41 35 43 37
rect 45 35 47 37
rect 38 33 47 35
rect 38 30 40 33
rect 9 19 11 24
rect 24 14 26 19
rect 31 14 33 19
rect 38 15 40 19
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 11 24 24 30
rect 13 19 24 24
rect 26 19 31 30
rect 33 19 38 30
rect 40 25 45 30
rect 40 23 47 25
rect 40 21 43 23
rect 45 21 47 23
rect 40 19 47 21
rect 13 11 22 19
rect 13 9 16 11
rect 18 9 22 11
rect 13 7 22 9
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 67 19 69
rect 33 71 39 73
rect 33 69 35 71
rect 37 69 39 71
rect 13 62 17 67
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 56 9 58
rect 4 50 9 56
rect 11 61 17 62
rect 33 62 39 69
rect 33 61 41 62
rect 11 50 19 61
rect 21 54 29 61
rect 21 52 24 54
rect 26 52 29 54
rect 21 50 29 52
rect 31 51 41 61
rect 43 60 50 62
rect 43 58 46 60
rect 48 58 50 60
rect 43 56 50 58
rect 43 51 48 56
rect 31 50 39 51
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 15 71
rect 17 69 35 71
rect 37 69 58 71
rect -2 68 58 69
rect 2 60 14 63
rect 2 58 4 60
rect 6 58 14 60
rect 2 57 14 58
rect 2 28 6 57
rect 33 50 47 54
rect 33 46 37 50
rect 25 45 37 46
rect 25 43 33 45
rect 35 43 37 45
rect 25 42 37 43
rect 41 38 47 46
rect 2 26 4 28
rect 2 17 6 26
rect 17 37 30 38
rect 17 35 21 37
rect 23 35 30 37
rect 17 34 30 35
rect 26 25 30 34
rect 34 37 47 38
rect 34 35 43 37
rect 45 35 47 37
rect 34 34 47 35
rect 34 25 38 34
rect -2 11 58 12
rect -2 9 16 11
rect 18 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 24 11 30
rect 24 19 26 30
rect 31 19 33 30
rect 38 19 40 30
<< pmos >>
rect 9 50 11 62
rect 19 50 21 61
rect 29 50 31 61
rect 41 51 43 62
<< polyct0 >>
rect 11 36 13 38
<< polyct1 >>
rect 33 43 35 45
rect 21 35 23 37
rect 43 35 45 37
<< ndifct0 >>
rect 43 21 45 23
<< ndifct1 >>
rect 4 26 6 28
rect 16 9 18 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 24 52 26 54
rect 46 58 48 60
<< pdifct1 >>
rect 15 69 17 71
rect 35 69 37 71
rect 4 58 6 60
<< alu0 >>
rect 23 60 50 61
rect 23 58 46 60
rect 48 58 50 60
rect 23 57 50 58
rect 23 54 27 57
rect 10 52 24 54
rect 26 52 27 54
rect 10 50 27 52
rect 10 38 14 50
rect 10 36 11 38
rect 13 36 14 38
rect 6 24 7 30
rect 10 29 14 36
rect 10 25 19 29
rect 15 21 19 25
rect 42 23 46 25
rect 42 21 43 23
rect 45 21 46 23
rect 15 17 46 21
<< labels >>
rlabel alu0 12 39 12 39 6 zn
rlabel alu0 25 55 25 55 6 zn
rlabel alu0 30 19 30 19 6 zn
rlabel alu0 36 59 36 59 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 36 20 36 6 a
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 28 28 28 6 a
rlabel alu1 36 28 36 28 6 c
rlabel alu1 28 44 28 44 6 b
rlabel alu1 36 52 36 52 6 b
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 40 44 40 6 c
rlabel alu1 44 52 44 52 6 b
<< end >>
