magic
tech scmos
timestamp 1199203007
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 11 66 13 70
rect 18 66 20 70
rect 25 66 27 70
rect 35 66 37 70
rect 42 66 44 70
rect 49 66 51 70
rect 11 27 13 38
rect 18 35 20 38
rect 25 35 27 38
rect 35 35 37 38
rect 18 32 21 35
rect 25 33 37 35
rect 19 27 21 32
rect 35 27 37 33
rect 9 25 15 27
rect 9 23 11 25
rect 13 23 15 25
rect 9 21 15 23
rect 19 25 25 27
rect 19 23 21 25
rect 23 23 25 25
rect 19 21 25 23
rect 31 25 37 27
rect 31 23 33 25
rect 35 23 37 25
rect 42 29 44 38
rect 49 35 51 38
rect 49 33 58 35
rect 52 31 54 33
rect 56 31 58 33
rect 52 29 58 31
rect 42 27 48 29
rect 42 25 44 27
rect 46 25 48 27
rect 42 23 48 25
rect 31 21 37 23
rect 9 18 11 21
rect 21 18 23 21
rect 31 18 33 21
rect 9 3 11 8
rect 21 3 23 8
rect 31 3 33 8
<< ndif >>
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 4 8 9 12
rect 11 8 21 18
rect 23 16 31 18
rect 23 14 26 16
rect 28 14 31 16
rect 23 8 31 14
rect 33 8 42 18
rect 13 7 19 8
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
rect 35 7 42 8
rect 35 5 37 7
rect 39 5 42 7
rect 35 3 42 5
<< pdif >>
rect 4 64 11 66
rect 4 62 6 64
rect 8 62 11 64
rect 4 57 11 62
rect 4 55 6 57
rect 8 55 11 57
rect 4 38 11 55
rect 13 38 18 66
rect 20 38 25 66
rect 27 57 35 66
rect 27 55 30 57
rect 32 55 35 57
rect 27 50 35 55
rect 27 48 30 50
rect 32 48 35 50
rect 27 38 35 48
rect 37 38 42 66
rect 44 38 49 66
rect 51 64 58 66
rect 51 62 54 64
rect 56 62 58 64
rect 51 57 58 62
rect 51 55 54 57
rect 56 55 58 57
rect 51 38 58 55
<< alu1 >>
rect -2 64 66 72
rect 2 48 30 50
rect 32 48 39 50
rect 2 46 39 48
rect 2 17 6 46
rect 10 38 55 42
rect 10 25 14 38
rect 51 34 55 38
rect 10 23 11 25
rect 13 23 14 25
rect 10 21 14 23
rect 18 30 47 34
rect 51 33 58 34
rect 51 31 54 33
rect 56 31 58 33
rect 51 30 58 31
rect 18 25 24 30
rect 43 27 47 30
rect 18 23 21 25
rect 23 23 24 25
rect 18 21 24 23
rect 31 25 39 26
rect 31 23 33 25
rect 35 23 39 25
rect 31 22 39 23
rect 43 25 44 27
rect 46 26 47 27
rect 46 25 55 26
rect 43 22 55 25
rect 34 18 39 22
rect 2 16 30 17
rect 2 14 4 16
rect 6 14 26 16
rect 28 14 30 16
rect 2 13 30 14
rect 34 13 47 18
rect -2 7 66 8
rect -2 5 15 7
rect 17 5 37 7
rect 39 5 53 7
rect 55 5 66 7
rect -2 0 66 5
<< ptie >>
rect 51 7 57 24
rect 51 5 53 7
rect 55 5 57 7
rect 51 3 57 5
<< nmos >>
rect 9 8 11 18
rect 21 8 23 18
rect 31 8 33 18
<< pmos >>
rect 11 38 13 66
rect 18 38 20 66
rect 25 38 27 66
rect 35 38 37 66
rect 42 38 44 66
rect 49 38 51 66
<< polyct1 >>
rect 11 23 13 25
rect 21 23 23 25
rect 33 23 35 25
rect 54 31 56 33
rect 44 25 46 27
<< ndifct1 >>
rect 4 14 6 16
rect 26 14 28 16
rect 15 5 17 7
rect 37 5 39 7
<< ptiect1 >>
rect 53 5 55 7
<< pdifct0 >>
rect 6 62 8 64
rect 6 55 8 57
rect 30 55 32 57
rect 54 62 56 64
rect 54 55 56 57
<< pdifct1 >>
rect 30 48 32 50
<< alu0 >>
rect 4 62 6 64
rect 8 62 10 64
rect 4 57 10 62
rect 52 62 54 64
rect 56 62 58 64
rect 4 55 6 57
rect 8 55 10 57
rect 4 54 10 55
rect 29 57 33 59
rect 29 55 30 57
rect 32 55 33 57
rect 29 50 33 55
rect 52 57 58 62
rect 52 55 54 57
rect 56 55 58 57
rect 52 54 58 55
<< labels >>
rlabel alu1 12 28 12 28 6 a
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 32 28 32 6 b
rlabel alu1 20 24 20 24 6 b
rlabel alu1 20 40 20 40 6 a
rlabel alu1 28 40 28 40 6 a
rlabel alu1 28 48 28 48 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 44 16 44 16 6 c
rlabel alu1 36 20 36 20 6 c
rlabel alu1 36 32 36 32 6 b
rlabel alu1 44 32 44 32 6 b
rlabel alu1 44 40 44 40 6 a
rlabel alu1 36 40 36 40 6 a
rlabel alu1 36 48 36 48 6 z
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 24 52 24 6 b
rlabel alu1 52 40 52 40 6 a
<< end >>
