magic
tech scmos
timestamp 1199203517
<< ab >>
rect 0 0 128 80
<< nwell >>
rect -5 36 133 88
<< pwell >>
rect -5 -8 133 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 72 70 74 74
rect 79 70 81 74
rect 89 70 91 74
rect 107 70 109 74
rect 117 70 119 74
rect 49 62 51 67
rect 39 49 41 52
rect 49 49 51 52
rect 39 47 51 49
rect 42 45 44 47
rect 46 45 48 47
rect 42 43 48 45
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 72 39 74 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 29 37 63 39
rect 69 37 75 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 10 24 12 33
rect 19 29 21 33
rect 37 29 39 37
rect 69 35 71 37
rect 73 35 75 37
rect 69 33 75 35
rect 49 31 55 33
rect 49 29 51 31
rect 53 29 55 31
rect 69 30 71 33
rect 79 30 81 42
rect 89 39 91 42
rect 89 37 95 39
rect 89 35 91 37
rect 93 35 95 37
rect 107 35 109 42
rect 117 39 119 42
rect 89 33 109 35
rect 113 37 119 39
rect 113 35 115 37
rect 117 35 119 37
rect 113 33 119 35
rect 101 30 103 33
rect 17 27 21 29
rect 17 24 19 27
rect 27 24 29 29
rect 49 27 55 29
rect 49 23 51 27
rect 37 12 39 16
rect 88 20 94 22
rect 88 18 90 20
rect 92 18 94 20
rect 117 27 119 33
rect 88 16 94 18
rect 10 6 12 11
rect 17 6 19 11
rect 27 8 29 11
rect 49 8 51 12
rect 69 11 71 16
rect 79 13 81 16
rect 88 13 90 16
rect 101 14 103 19
rect 79 11 90 13
rect 117 11 119 16
rect 27 6 51 8
<< ndif >>
rect 32 24 37 29
rect 2 11 10 24
rect 12 11 17 24
rect 19 21 27 24
rect 19 19 22 21
rect 24 19 27 21
rect 19 11 27 19
rect 29 22 37 24
rect 29 20 32 22
rect 34 20 37 22
rect 29 16 37 20
rect 39 23 47 29
rect 39 16 49 23
rect 29 11 34 16
rect 41 14 43 16
rect 45 14 49 16
rect 41 12 49 14
rect 51 21 58 23
rect 64 22 69 30
rect 51 19 54 21
rect 56 19 58 21
rect 51 17 58 19
rect 62 20 69 22
rect 62 18 64 20
rect 66 18 69 20
rect 51 12 56 17
rect 62 16 69 18
rect 71 28 79 30
rect 71 26 74 28
rect 76 26 79 28
rect 71 16 79 26
rect 81 28 88 30
rect 81 26 84 28
rect 86 26 88 28
rect 81 24 88 26
rect 94 28 101 30
rect 94 26 96 28
rect 98 26 101 28
rect 94 24 101 26
rect 81 16 86 24
rect 96 19 101 24
rect 103 27 115 30
rect 103 19 117 27
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
rect 105 16 117 19
rect 119 22 124 27
rect 119 20 126 22
rect 119 18 122 20
rect 124 18 126 20
rect 119 16 126 18
rect 105 11 115 16
rect 105 9 109 11
rect 111 9 115 11
rect 105 7 115 9
<< pdif >>
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 42 9 58
rect 11 54 19 70
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 46 29 70
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 52 39 59
rect 41 62 46 70
rect 67 63 72 70
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 52 49 55
rect 51 60 58 62
rect 51 58 54 60
rect 56 58 58 60
rect 51 52 58 58
rect 65 61 72 63
rect 65 59 67 61
rect 69 59 72 61
rect 65 54 72 59
rect 65 52 67 54
rect 69 52 72 54
rect 31 42 37 52
rect 65 42 72 52
rect 74 42 79 70
rect 81 61 89 70
rect 81 59 84 61
rect 86 59 89 61
rect 81 54 89 59
rect 81 52 84 54
rect 86 52 89 54
rect 81 42 89 52
rect 91 58 96 70
rect 91 56 98 58
rect 91 54 94 56
rect 96 54 98 56
rect 91 52 98 54
rect 91 42 96 52
rect 102 48 107 70
rect 100 46 107 48
rect 100 44 102 46
rect 104 44 107 46
rect 100 42 107 44
rect 109 68 117 70
rect 109 66 112 68
rect 114 66 117 68
rect 109 61 117 66
rect 109 59 112 61
rect 114 59 117 61
rect 109 42 117 59
rect 119 55 124 70
rect 119 53 126 55
rect 119 51 122 53
rect 124 51 126 53
rect 119 46 126 51
rect 119 44 122 46
rect 124 44 126 46
rect 119 42 126 44
<< alu1 >>
rect -2 81 130 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 130 81
rect -2 68 130 79
rect 2 54 18 55
rect 2 52 14 54
rect 16 52 18 54
rect 2 50 18 52
rect 2 22 6 50
rect 41 47 54 48
rect 41 45 44 47
rect 46 45 54 47
rect 41 42 54 45
rect 2 21 26 22
rect 2 19 22 21
rect 24 19 26 21
rect 2 18 26 19
rect 50 31 54 42
rect 82 41 94 47
rect 50 29 51 31
rect 53 29 54 31
rect 50 27 54 29
rect 90 37 94 41
rect 90 35 91 37
rect 93 35 94 37
rect 90 33 94 35
rect 114 37 118 47
rect 114 35 115 37
rect 117 35 118 37
rect 114 31 118 35
rect 106 25 118 31
rect -2 11 130 12
rect -2 9 4 11
rect 6 9 109 11
rect 111 9 130 11
rect -2 1 130 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 130 1
rect -2 -2 130 -1
<< ptie >>
rect 0 1 128 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 128 1
rect 0 -3 128 -1
<< ntie >>
rect 0 81 128 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 128 81
rect 0 77 128 79
<< nmos >>
rect 10 11 12 24
rect 17 11 19 24
rect 27 11 29 24
rect 37 16 39 29
rect 49 12 51 23
rect 69 16 71 30
rect 79 16 81 30
rect 101 19 103 30
rect 117 16 119 27
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 52 41 70
rect 49 52 51 62
rect 72 42 74 70
rect 79 42 81 70
rect 89 42 91 70
rect 107 42 109 70
rect 117 42 119 70
<< polyct0 >>
rect 59 39 61 41
rect 11 35 13 37
rect 21 35 23 37
rect 71 35 73 37
rect 90 18 92 20
<< polyct1 >>
rect 44 45 46 47
rect 51 29 53 31
rect 91 35 93 37
rect 115 35 117 37
<< ndifct0 >>
rect 32 20 34 22
rect 43 14 45 16
rect 54 19 56 21
rect 64 18 66 20
rect 74 26 76 28
rect 84 26 86 28
rect 96 26 98 28
rect 122 18 124 20
<< ndifct1 >>
rect 22 19 24 21
rect 4 9 6 11
rect 109 9 111 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
<< pdifct0 >>
rect 4 60 6 62
rect 24 44 26 46
rect 34 66 36 68
rect 34 59 36 61
rect 44 55 46 57
rect 54 58 56 60
rect 67 59 69 61
rect 67 52 69 54
rect 84 59 86 61
rect 84 52 86 54
rect 94 54 96 56
rect 102 44 104 46
rect 112 66 114 68
rect 112 59 114 61
rect 122 51 124 53
rect 122 44 124 46
<< pdifct1 >>
rect 14 52 16 54
<< alu0 >>
rect 32 66 34 68
rect 36 66 38 68
rect 2 62 27 63
rect 2 60 4 62
rect 6 60 27 62
rect 2 59 27 60
rect 23 55 27 59
rect 32 61 38 66
rect 32 59 34 61
rect 36 59 38 61
rect 53 60 57 68
rect 32 58 38 59
rect 43 57 47 59
rect 43 55 44 57
rect 46 55 47 57
rect 53 58 54 60
rect 56 58 57 60
rect 53 56 57 58
rect 66 61 70 68
rect 110 66 112 68
rect 114 66 116 68
rect 66 59 67 61
rect 69 59 70 61
rect 23 51 47 55
rect 66 54 70 59
rect 83 61 88 63
rect 83 59 84 61
rect 86 59 88 61
rect 83 55 88 59
rect 110 61 116 66
rect 110 59 112 61
rect 114 59 116 61
rect 110 58 116 59
rect 66 52 67 54
rect 69 52 70 54
rect 10 46 28 47
rect 10 44 24 46
rect 26 44 28 46
rect 10 43 28 44
rect 10 37 14 43
rect 32 38 36 51
rect 66 50 70 52
rect 74 54 88 55
rect 74 52 84 54
rect 86 52 88 54
rect 74 51 88 52
rect 93 56 97 58
rect 93 54 94 56
rect 96 55 97 56
rect 96 54 126 55
rect 93 53 126 54
rect 93 51 122 53
rect 124 51 126 53
rect 74 46 78 51
rect 61 43 78 46
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 19 37 44 38
rect 19 35 21 37
rect 23 35 44 37
rect 19 34 44 35
rect 10 26 35 30
rect 31 22 35 26
rect 31 20 32 22
rect 34 20 35 22
rect 40 24 44 34
rect 58 42 78 43
rect 58 41 65 42
rect 58 39 59 41
rect 61 39 65 41
rect 58 37 65 39
rect 61 29 65 37
rect 69 37 86 38
rect 69 35 71 37
rect 73 35 86 37
rect 69 34 86 35
rect 82 29 86 34
rect 98 46 106 47
rect 98 44 102 46
rect 104 44 106 46
rect 98 43 106 44
rect 98 29 102 43
rect 121 46 126 51
rect 121 44 122 46
rect 124 44 126 46
rect 121 42 126 44
rect 61 28 78 29
rect 61 26 74 28
rect 76 26 78 28
rect 61 25 78 26
rect 82 28 102 29
rect 82 26 84 28
rect 86 26 96 28
rect 98 26 102 28
rect 82 25 102 26
rect 40 21 57 24
rect 122 21 126 42
rect 40 20 54 21
rect 31 18 35 20
rect 53 19 54 20
rect 56 19 57 21
rect 53 17 57 19
rect 62 20 126 21
rect 62 18 64 20
rect 66 18 90 20
rect 92 18 122 20
rect 124 18 126 20
rect 62 17 126 18
rect 41 16 47 17
rect 41 14 43 16
rect 45 14 47 16
rect 41 12 47 14
<< labels >>
rlabel polyct0 12 36 12 36 6 zn
rlabel alu0 33 24 33 24 6 zn
rlabel alu0 31 36 31 36 6 cn
rlabel alu0 19 45 19 45 6 zn
rlabel alu0 14 61 14 61 6 cn
rlabel alu0 45 55 45 55 6 cn
rlabel ndifct0 55 20 55 20 6 cn
rlabel alu0 61 40 61 40 6 iz
rlabel alu0 69 27 69 27 6 iz
rlabel alu0 77 36 77 36 6 bn
rlabel alu0 81 53 81 53 6 iz
rlabel alu0 85 57 85 57 6 iz
rlabel alu0 92 27 92 27 6 bn
rlabel alu0 94 19 94 19 6 an
rlabel alu0 102 45 102 45 6 bn
rlabel alu0 124 36 124 36 6 an
rlabel alu0 109 53 109 53 6 an
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 52 40 52 40 6 c
rlabel alu1 44 44 44 44 6 c
rlabel alu1 64 6 64 6 6 vss
rlabel alu1 92 40 92 40 6 b
rlabel alu1 84 44 84 44 6 b
rlabel alu1 64 74 64 74 6 vdd
rlabel polyct1 116 36 116 36 6 a
rlabel alu1 108 28 108 28 6 a
<< end >>
