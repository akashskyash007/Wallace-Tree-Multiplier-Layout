magic
tech scmos
timestamp 1199544109
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -2 48 102 104
<< pwell >>
rect -2 -4 102 48
<< poly >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 63 85 65 88
rect 75 85 77 88
rect 87 85 89 88
rect 35 63 37 75
rect 45 65 51 67
rect 45 63 47 65
rect 49 63 51 65
rect 63 63 65 65
rect 35 61 41 63
rect 45 61 65 63
rect 35 59 37 61
rect 39 59 41 61
rect 35 57 41 59
rect 75 57 77 65
rect 87 63 89 65
rect 81 61 89 63
rect 81 59 83 61
rect 85 59 89 61
rect 81 57 89 59
rect 35 55 77 57
rect 11 47 13 55
rect 23 47 25 55
rect 65 53 67 55
rect 69 53 71 55
rect 65 51 71 53
rect 91 47 97 49
rect 11 45 93 47
rect 95 45 97 47
rect 91 43 97 45
rect 11 37 61 39
rect 11 25 13 37
rect 23 25 25 37
rect 55 35 57 37
rect 59 35 61 37
rect 55 33 61 35
rect 65 37 89 39
rect 65 35 67 37
rect 69 35 71 37
rect 65 33 71 35
rect 29 31 37 33
rect 29 29 31 31
rect 33 29 37 31
rect 29 27 37 29
rect 45 31 51 33
rect 45 29 47 31
rect 49 29 51 31
rect 75 31 83 33
rect 75 29 79 31
rect 81 29 83 31
rect 45 27 65 29
rect 35 25 37 27
rect 63 25 65 27
rect 75 27 83 29
rect 75 25 77 27
rect 87 25 89 37
rect 35 12 37 15
rect 63 12 65 15
rect 75 12 77 15
rect 87 12 89 15
rect 11 2 13 5
rect 23 2 25 5
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 11 11 19
rect 3 9 5 11
rect 7 9 11 11
rect 3 5 11 9
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 5 23 19
rect 25 15 35 25
rect 37 21 45 25
rect 37 19 41 21
rect 43 19 45 21
rect 37 15 45 19
rect 55 21 63 25
rect 55 19 57 21
rect 59 19 63 21
rect 55 15 63 19
rect 65 15 75 25
rect 77 21 87 25
rect 77 19 81 21
rect 83 19 87 21
rect 77 15 87 19
rect 89 21 97 25
rect 89 19 93 21
rect 95 19 97 21
rect 89 15 97 19
rect 25 11 33 15
rect 25 9 29 11
rect 31 9 33 11
rect 67 11 73 15
rect 67 9 69 11
rect 71 9 73 11
rect 25 5 33 9
rect 67 7 73 9
<< pdif >>
rect 3 91 11 95
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 81 23 95
rect 13 79 17 81
rect 19 79 23 81
rect 13 71 23 79
rect 13 69 17 71
rect 19 69 23 71
rect 13 61 23 69
rect 13 59 17 61
rect 19 59 23 61
rect 13 55 23 59
rect 25 91 35 95
rect 25 89 29 91
rect 31 89 35 91
rect 25 75 35 89
rect 37 81 45 95
rect 79 91 85 95
rect 79 89 81 91
rect 83 89 85 91
rect 79 85 85 89
rect 37 79 41 81
rect 43 79 45 81
rect 37 75 45 79
rect 55 81 63 85
rect 55 79 57 81
rect 59 79 63 81
rect 25 55 33 75
rect 55 71 63 79
rect 55 69 57 71
rect 59 69 63 71
rect 55 65 63 69
rect 65 81 75 85
rect 65 79 69 81
rect 71 79 75 81
rect 65 71 75 79
rect 65 69 69 71
rect 71 69 75 71
rect 65 65 75 69
rect 77 65 87 85
rect 89 81 97 85
rect 89 79 93 81
rect 95 79 97 81
rect 89 71 97 79
rect 89 69 93 71
rect 95 69 97 71
rect 89 65 97 69
<< alu1 >>
rect -2 95 102 100
rect -2 93 53 95
rect 55 93 69 95
rect 71 93 102 95
rect -2 91 102 93
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 81 91
rect 83 89 102 91
rect -2 88 102 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 16 81 22 82
rect 16 79 17 81
rect 19 79 22 81
rect 16 78 22 79
rect 18 72 22 78
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 16 71 22 72
rect 16 69 17 71
rect 19 69 22 71
rect 16 68 22 69
rect 18 62 22 68
rect 4 59 5 61
rect 7 59 8 61
rect 4 58 8 59
rect 16 61 22 62
rect 16 59 17 61
rect 19 59 22 61
rect 16 58 22 59
rect 18 22 22 58
rect 4 21 8 22
rect 4 19 5 21
rect 7 19 8 21
rect 4 12 8 19
rect 16 21 22 22
rect 16 19 17 21
rect 19 19 22 21
rect 16 18 22 19
rect 28 62 32 82
rect 40 81 49 82
rect 40 79 41 81
rect 43 79 49 81
rect 40 78 49 79
rect 56 81 60 82
rect 56 79 57 81
rect 59 79 60 81
rect 56 78 60 79
rect 68 81 72 82
rect 92 81 96 82
rect 68 79 69 81
rect 71 79 93 81
rect 95 79 96 81
rect 68 78 72 79
rect 92 78 96 79
rect 47 66 49 78
rect 57 72 59 78
rect 69 72 71 78
rect 93 72 95 78
rect 56 71 60 72
rect 56 69 57 71
rect 59 69 60 71
rect 56 68 60 69
rect 68 71 72 72
rect 68 69 69 71
rect 71 69 72 71
rect 68 68 72 69
rect 46 65 50 66
rect 46 63 47 65
rect 49 63 50 65
rect 46 62 50 63
rect 28 61 40 62
rect 28 59 37 61
rect 39 59 40 61
rect 28 58 40 59
rect 28 32 32 58
rect 47 32 49 62
rect 57 38 59 68
rect 78 62 82 72
rect 92 71 96 72
rect 92 69 93 71
rect 95 69 96 71
rect 92 68 96 69
rect 78 61 86 62
rect 78 59 83 61
rect 85 59 86 61
rect 78 58 86 59
rect 66 55 70 56
rect 66 53 67 55
rect 69 53 70 55
rect 66 52 70 53
rect 67 38 69 52
rect 56 37 60 38
rect 56 35 57 37
rect 59 35 60 37
rect 56 34 60 35
rect 66 37 70 38
rect 66 35 67 37
rect 69 35 70 37
rect 66 34 70 35
rect 28 31 34 32
rect 28 29 31 31
rect 33 29 34 31
rect 28 28 34 29
rect 46 31 50 32
rect 46 29 47 31
rect 49 29 50 31
rect 46 28 50 29
rect 28 18 32 28
rect 47 22 49 28
rect 57 22 59 34
rect 78 31 82 58
rect 93 48 95 68
rect 92 47 96 48
rect 92 45 93 47
rect 95 45 96 47
rect 92 44 96 45
rect 78 29 79 31
rect 81 29 82 31
rect 78 28 82 29
rect 93 22 95 44
rect 40 21 49 22
rect 40 19 41 21
rect 43 19 49 21
rect 40 18 49 19
rect 56 21 60 22
rect 80 21 84 22
rect 56 19 57 21
rect 59 19 81 21
rect 83 19 84 21
rect 56 18 60 19
rect 80 18 84 19
rect 92 21 96 22
rect 92 19 93 21
rect 95 19 96 21
rect 92 18 96 19
rect -2 11 102 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 69 11
rect 71 9 102 11
rect -2 7 102 9
rect -2 5 41 7
rect 43 5 57 7
rect 59 5 81 7
rect 83 5 93 7
rect 95 5 102 7
rect -2 0 102 5
<< ptie >>
rect 39 7 61 9
rect 79 7 97 9
rect 39 5 41 7
rect 43 5 57 7
rect 59 5 61 7
rect 39 3 61 5
rect 79 5 81 7
rect 83 5 93 7
rect 95 5 97 7
rect 79 3 97 5
<< ntie >>
rect 51 95 73 97
rect 51 93 53 95
rect 55 93 69 95
rect 71 93 73 95
rect 51 91 73 93
<< nmos >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 15 37 25
rect 63 15 65 25
rect 75 15 77 25
rect 87 15 89 25
<< pmos >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 75 37 95
rect 63 65 65 85
rect 75 65 77 85
rect 87 65 89 85
<< polyct1 >>
rect 47 63 49 65
rect 37 59 39 61
rect 83 59 85 61
rect 67 53 69 55
rect 93 45 95 47
rect 57 35 59 37
rect 67 35 69 37
rect 31 29 33 31
rect 47 29 49 31
rect 79 29 81 31
<< ndifct1 >>
rect 5 19 7 21
rect 5 9 7 11
rect 17 19 19 21
rect 41 19 43 21
rect 57 19 59 21
rect 81 19 83 21
rect 93 19 95 21
rect 29 9 31 11
rect 69 9 71 11
<< ntiect1 >>
rect 53 93 55 95
rect 69 93 71 95
<< ptiect1 >>
rect 41 5 43 7
rect 57 5 59 7
rect 81 5 83 7
rect 93 5 95 7
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 5 69 7 71
rect 5 59 7 61
rect 17 79 19 81
rect 17 69 19 71
rect 17 59 19 61
rect 29 89 31 91
rect 81 89 83 91
rect 41 79 43 81
rect 57 79 59 81
rect 57 69 59 71
rect 69 79 71 81
rect 69 69 71 71
rect 93 79 95 81
rect 93 69 95 71
<< labels >>
rlabel alu1 20 50 20 50 6 q
rlabel alu1 30 50 30 50 6 cmd
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 50 94 50 94 6 vdd
rlabel alu1 80 50 80 50 6 i
<< end >>
