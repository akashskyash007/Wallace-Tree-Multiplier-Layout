magic
tech scmos
timestamp 1199203091
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 12 70 14 74
rect 22 70 24 74
rect 29 70 31 74
rect 12 49 14 55
rect 9 47 15 49
rect 9 45 11 47
rect 13 45 15 47
rect 9 43 15 45
rect 9 23 11 43
rect 39 68 41 72
rect 39 47 41 50
rect 39 45 55 47
rect 49 43 51 45
rect 53 43 55 45
rect 22 39 24 42
rect 17 37 24 39
rect 17 35 19 37
rect 21 35 24 37
rect 17 33 24 35
rect 29 39 31 42
rect 49 41 55 43
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 19 23 21 33
rect 29 23 31 33
rect 49 30 51 41
rect 49 16 51 21
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
<< ndif >>
rect 42 28 49 30
rect 42 26 44 28
rect 46 26 49 28
rect 42 24 49 26
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 21 19 23
rect 11 19 14 21
rect 16 19 19 21
rect 11 10 19 19
rect 21 14 29 23
rect 21 12 24 14
rect 26 12 29 14
rect 21 10 29 12
rect 31 21 38 23
rect 44 21 49 24
rect 51 25 58 30
rect 51 23 54 25
rect 56 23 58 25
rect 51 21 58 23
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
rect 31 10 36 17
<< pdif >>
rect 4 68 12 70
rect 4 66 7 68
rect 9 66 12 68
rect 4 55 12 66
rect 14 61 22 70
rect 14 59 17 61
rect 19 59 22 61
rect 14 55 22 59
rect 17 42 22 55
rect 24 42 29 70
rect 31 68 37 70
rect 31 66 39 68
rect 31 64 34 66
rect 36 64 39 66
rect 31 59 39 64
rect 31 57 34 59
rect 36 57 39 59
rect 31 50 39 57
rect 41 63 46 68
rect 41 61 48 63
rect 41 59 44 61
rect 46 59 48 61
rect 41 54 48 59
rect 41 52 44 54
rect 46 52 48 54
rect 41 50 48 52
rect 31 42 37 50
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 61 23 62
rect 2 59 17 61
rect 19 59 23 61
rect 2 58 23 59
rect 2 22 6 58
rect 10 47 14 49
rect 10 45 11 47
rect 13 45 14 47
rect 58 47 62 55
rect 10 30 14 45
rect 25 37 39 38
rect 25 35 31 37
rect 33 35 39 37
rect 25 34 39 35
rect 10 26 23 30
rect 33 26 39 34
rect 50 45 62 47
rect 50 43 51 45
rect 53 43 62 45
rect 50 41 62 43
rect 2 21 8 22
rect 2 19 4 21
rect 6 19 8 21
rect 2 17 8 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 10 11 23
rect 19 10 21 23
rect 29 10 31 23
rect 49 21 51 30
<< pmos >>
rect 12 55 14 70
rect 22 42 24 70
rect 29 42 31 70
rect 39 50 41 68
<< polyct0 >>
rect 19 35 21 37
<< polyct1 >>
rect 11 45 13 47
rect 51 43 53 45
rect 31 35 33 37
<< ndifct0 >>
rect 44 26 46 28
rect 14 19 16 21
rect 24 12 26 14
rect 54 23 56 25
rect 34 19 36 21
<< ndifct1 >>
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 7 66 9 68
rect 34 64 36 66
rect 34 57 36 59
rect 44 59 46 61
rect 44 52 46 54
<< pdifct1 >>
rect 17 59 19 61
<< alu0 >>
rect 5 66 7 68
rect 9 66 11 68
rect 5 65 11 66
rect 33 66 37 68
rect 33 64 34 66
rect 36 64 37 66
rect 33 59 37 64
rect 33 57 34 59
rect 36 57 37 59
rect 33 55 37 57
rect 43 61 47 63
rect 43 59 44 61
rect 46 59 47 61
rect 43 54 47 59
rect 43 52 44 54
rect 46 52 47 54
rect 43 46 47 52
rect 18 42 47 46
rect 18 37 22 42
rect 18 35 19 37
rect 21 35 22 37
rect 18 33 22 35
rect 43 28 47 42
rect 43 26 44 28
rect 46 26 47 28
rect 43 24 47 26
rect 53 25 57 27
rect 53 23 54 25
rect 56 23 57 25
rect 12 21 38 22
rect 12 19 14 21
rect 16 19 34 21
rect 36 19 38 21
rect 12 18 38 19
rect 22 14 28 15
rect 22 12 24 14
rect 26 12 28 14
rect 53 12 57 23
<< labels >>
rlabel alu0 25 20 25 20 6 n1
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 36 28 36 6 a1
rlabel alu1 20 60 20 60 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 32 36 32 6 a1
rlabel alu1 32 74 32 74 6 vdd
rlabel polyct1 52 44 52 44 6 a2
rlabel alu1 60 48 60 48 6 a2
<< end >>
