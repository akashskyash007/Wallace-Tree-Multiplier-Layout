magic
tech scmos
timestamp 1199202724
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 30 66 32 70
rect 40 66 42 70
rect 9 35 11 38
rect 19 35 21 38
rect 30 35 32 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 32 35
rect 19 31 27 33
rect 29 31 32 33
rect 40 35 42 38
rect 40 33 47 35
rect 40 31 43 33
rect 45 31 47 33
rect 19 29 32 31
rect 13 25 15 29
rect 20 25 22 29
rect 30 25 32 29
rect 37 29 47 31
rect 37 25 39 29
rect 13 2 15 7
rect 20 2 22 7
rect 30 2 32 7
rect 37 2 39 7
<< ndif >>
rect 4 10 13 25
rect 4 8 7 10
rect 9 8 13 10
rect 4 7 13 8
rect 15 7 20 25
rect 22 17 30 25
rect 22 15 25 17
rect 27 15 30 17
rect 22 7 30 15
rect 32 7 37 25
rect 39 18 47 25
rect 39 16 42 18
rect 44 16 47 18
rect 39 11 47 16
rect 39 9 42 11
rect 44 9 47 11
rect 39 7 47 9
rect 4 5 11 7
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 56 9 62
rect 2 54 4 56
rect 6 54 9 56
rect 2 38 9 54
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 64 30 66
rect 21 62 24 64
rect 26 62 30 64
rect 21 57 30 62
rect 21 55 24 57
rect 26 55 30 57
rect 21 38 30 55
rect 32 56 40 66
rect 32 54 35 56
rect 37 54 40 56
rect 32 49 40 54
rect 32 47 35 49
rect 37 47 40 49
rect 32 38 40 47
rect 42 64 50 66
rect 42 62 45 64
rect 47 62 50 64
rect 42 57 50 62
rect 42 55 45 57
rect 47 55 50 57
rect 42 38 50 55
<< alu1 >>
rect -2 64 58 72
rect 34 56 39 59
rect 34 54 35 56
rect 37 54 39 56
rect 34 50 39 54
rect 12 49 39 50
rect 12 47 14 49
rect 16 47 35 49
rect 37 47 39 49
rect 12 46 39 47
rect 12 43 18 46
rect 2 42 18 43
rect 2 40 14 42
rect 16 40 18 42
rect 2 39 18 40
rect 2 18 6 39
rect 25 38 39 42
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 25 33 31 38
rect 25 31 27 33
rect 29 31 31 33
rect 25 30 31 31
rect 41 33 47 34
rect 41 31 43 33
rect 45 31 47 33
rect 41 26 47 31
rect 10 22 47 26
rect 2 17 31 18
rect 2 15 25 17
rect 27 15 31 17
rect 2 14 31 15
rect -2 0 58 8
<< nmos >>
rect 13 7 15 25
rect 20 7 22 25
rect 30 7 32 25
rect 37 7 39 25
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 30 38 32 66
rect 40 38 42 66
<< polyct1 >>
rect 11 31 13 33
rect 27 31 29 33
rect 43 31 45 33
<< ndifct0 >>
rect 7 8 9 10
rect 42 16 44 18
rect 42 9 44 11
<< ndifct1 >>
rect 25 15 27 17
<< pdifct0 >>
rect 4 62 6 64
rect 4 54 6 56
rect 24 62 26 64
rect 24 55 26 57
rect 45 62 47 64
rect 45 55 47 57
<< pdifct1 >>
rect 14 47 16 49
rect 14 40 16 42
rect 35 54 37 56
rect 35 47 37 49
<< alu0 >>
rect 3 62 4 64
rect 6 62 7 64
rect 3 56 7 62
rect 3 54 4 56
rect 6 54 7 56
rect 22 62 24 64
rect 26 62 28 64
rect 22 57 28 62
rect 43 62 45 64
rect 47 62 49 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 43 57 49 62
rect 43 55 45 57
rect 47 55 49 57
rect 43 54 49 55
rect 3 52 7 54
rect 40 18 46 19
rect 40 16 42 18
rect 44 16 46 18
rect 40 11 46 16
rect 5 10 11 11
rect 5 8 7 10
rect 9 8 11 10
rect 40 9 42 11
rect 44 9 46 11
rect 40 8 46 9
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 20 24 20 24 6 a
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 16 28 16 6 z
rlabel alu1 28 24 28 24 6 a
rlabel alu1 36 24 36 24 6 a
rlabel alu1 36 40 36 40 6 b
rlabel alu1 28 36 28 36 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 28 44 28 6 a
<< end >>
