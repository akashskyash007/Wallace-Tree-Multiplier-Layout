magic
tech scmos
timestamp 1199202552
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 57 11 62
rect 19 57 21 62
rect 29 57 31 62
rect 9 40 11 43
rect 2 38 11 40
rect 19 39 21 43
rect 2 36 4 38
rect 6 36 11 38
rect 2 34 11 36
rect 9 30 11 34
rect 16 37 23 39
rect 16 35 19 37
rect 21 35 23 37
rect 16 33 23 35
rect 16 30 18 33
rect 29 31 31 43
rect 28 29 34 31
rect 28 27 30 29
rect 32 27 34 29
rect 28 25 34 27
rect 28 22 30 25
rect 9 14 11 18
rect 16 14 18 18
rect 28 10 30 15
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 18 9 24
rect 11 18 16 30
rect 18 22 26 30
rect 18 18 28 22
rect 20 15 28 18
rect 30 20 38 22
rect 30 18 34 20
rect 36 18 38 20
rect 30 15 38 18
rect 20 11 26 15
rect 20 9 22 11
rect 24 9 26 11
rect 20 7 26 9
<< pdif >>
rect 2 71 8 73
rect 2 69 4 71
rect 6 69 8 71
rect 2 67 8 69
rect 2 57 7 67
rect 2 43 9 57
rect 11 54 19 57
rect 11 52 14 54
rect 16 52 19 54
rect 11 47 19 52
rect 11 45 14 47
rect 16 45 19 47
rect 11 43 19 45
rect 21 55 29 57
rect 21 53 24 55
rect 26 53 29 55
rect 21 43 29 53
rect 31 49 36 57
rect 31 47 38 49
rect 31 45 34 47
rect 36 45 38 47
rect 31 43 38 45
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 71 42 79
rect -2 69 4 71
rect 6 69 42 71
rect -2 68 42 69
rect 2 58 15 63
rect 2 38 6 58
rect 10 45 14 47
rect 16 45 23 47
rect 10 42 23 45
rect 2 36 4 38
rect 2 33 6 36
rect 10 29 14 42
rect 2 28 14 29
rect 2 26 4 28
rect 6 26 14 28
rect 2 25 14 26
rect 34 31 38 39
rect 26 29 38 31
rect 26 27 30 29
rect 32 27 38 29
rect 26 25 38 27
rect -2 11 42 12
rect -2 9 22 11
rect 24 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 18 11 30
rect 16 18 18 30
rect 28 15 30 22
<< pmos >>
rect 9 43 11 57
rect 19 43 21 57
rect 29 43 31 57
<< polyct0 >>
rect 19 35 21 37
<< polyct1 >>
rect 4 36 6 38
rect 30 27 32 29
<< ndifct0 >>
rect 34 18 36 20
<< ndifct1 >>
rect 4 26 6 28
rect 22 9 24 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 52 16 54
rect 24 53 26 55
rect 34 45 36 47
<< pdifct1 >>
rect 4 69 6 71
rect 14 45 16 47
<< alu0 >>
rect 23 55 27 68
rect 12 54 18 55
rect 12 52 14 54
rect 16 52 18 54
rect 12 47 18 52
rect 23 53 24 55
rect 26 53 27 55
rect 23 51 27 53
rect 32 47 38 48
rect 26 45 34 47
rect 36 45 38 47
rect 26 43 38 45
rect 6 34 7 40
rect 26 39 30 43
rect 18 37 30 39
rect 18 35 19 37
rect 21 35 30 37
rect 18 21 22 35
rect 18 20 38 21
rect 18 18 34 20
rect 36 18 38 20
rect 18 17 38 18
<< labels >>
rlabel alu0 20 28 20 28 6 an
rlabel alu0 28 19 28 19 6 an
rlabel alu0 35 45 35 45 6 an
rlabel alu1 4 48 4 48 6 b
rlabel alu1 12 36 12 36 6 z
rlabel alu1 12 60 12 60 6 b
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 28 28 28 6 a
rlabel alu1 20 44 20 44 6 z
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 32 36 32 6 a
<< end >>
