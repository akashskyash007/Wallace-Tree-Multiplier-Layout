magic
tech scmos
timestamp 1199203057
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 18 66 20 70
rect 25 66 27 70
rect 32 66 34 70
rect 39 66 41 70
rect 18 41 20 44
rect 9 39 20 41
rect 9 37 11 39
rect 13 37 15 39
rect 9 35 15 37
rect 25 35 27 44
rect 9 21 11 35
rect 19 33 27 35
rect 19 31 21 33
rect 23 32 27 33
rect 23 31 25 32
rect 19 29 25 31
rect 19 21 21 29
rect 32 28 34 44
rect 39 41 41 44
rect 39 39 47 41
rect 39 37 43 39
rect 45 37 47 39
rect 39 35 47 37
rect 29 26 35 28
rect 29 24 31 26
rect 33 24 35 26
rect 29 22 35 24
rect 29 19 31 22
rect 39 19 41 35
rect 9 11 11 15
rect 19 11 21 15
rect 29 8 31 13
rect 39 8 41 13
<< ndif >>
rect 2 19 9 21
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 19 19 21
rect 11 17 14 19
rect 16 17 19 19
rect 11 15 19 17
rect 21 19 27 21
rect 21 15 29 19
rect 23 13 29 15
rect 31 17 39 19
rect 31 15 34 17
rect 36 15 39 17
rect 31 13 39 15
rect 41 13 50 19
rect 23 9 27 13
rect 21 7 27 9
rect 21 5 23 7
rect 25 5 27 7
rect 21 3 27 5
rect 44 7 50 13
rect 44 5 46 7
rect 48 5 50 7
rect 44 3 50 5
<< pdif >>
rect 13 59 18 66
rect 11 57 18 59
rect 11 55 13 57
rect 15 55 18 57
rect 11 53 18 55
rect 13 44 18 53
rect 20 44 25 66
rect 27 44 32 66
rect 34 44 39 66
rect 41 64 48 66
rect 41 62 44 64
rect 46 62 48 64
rect 41 56 48 62
rect 41 54 44 56
rect 46 54 48 56
rect 41 44 48 54
<< alu1 >>
rect -2 67 58 72
rect -2 65 5 67
rect 7 65 58 67
rect -2 64 58 65
rect 2 57 17 59
rect 2 55 13 57
rect 15 55 17 57
rect 2 54 17 55
rect 2 30 6 54
rect 10 46 23 50
rect 10 39 14 46
rect 34 42 38 59
rect 10 37 11 39
rect 13 37 14 39
rect 10 35 14 37
rect 22 38 38 42
rect 42 39 46 43
rect 42 37 43 39
rect 45 37 46 39
rect 42 34 46 37
rect 2 26 17 30
rect 33 30 46 34
rect 13 19 17 26
rect 25 24 31 26
rect 33 24 47 26
rect 25 22 47 24
rect 13 17 14 19
rect 16 18 17 19
rect 16 17 38 18
rect 13 15 34 17
rect 36 15 38 17
rect 13 14 38 15
rect 42 13 47 22
rect -2 7 58 8
rect -2 5 5 7
rect 7 5 13 7
rect 15 5 23 7
rect 25 5 46 7
rect 48 5 58 7
rect -2 0 58 5
<< ptie >>
rect 3 7 17 9
rect 3 5 5 7
rect 7 5 13 7
rect 15 5 17 7
rect 3 3 17 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 15 11 21
rect 19 15 21 21
rect 29 13 31 19
rect 39 13 41 19
<< pmos >>
rect 18 44 20 66
rect 25 44 27 66
rect 32 44 34 66
rect 39 44 41 66
<< polyct0 >>
rect 21 31 23 33
<< polyct1 >>
rect 11 37 13 39
rect 43 37 45 39
rect 31 24 33 26
<< ndifct0 >>
rect 4 17 6 19
<< ndifct1 >>
rect 14 17 16 19
rect 34 15 36 17
rect 23 5 25 7
rect 46 5 48 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
rect 13 5 15 7
<< pdifct0 >>
rect 44 62 46 64
rect 44 54 46 56
<< pdifct1 >>
rect 13 55 15 57
<< alu0 >>
rect 43 62 44 64
rect 46 62 47 64
rect 43 56 47 62
rect 43 54 44 56
rect 46 54 47 56
rect 43 52 47 54
rect 20 38 22 42
rect 20 33 24 38
rect 20 31 21 33
rect 23 31 24 33
rect 20 29 24 31
rect 29 26 35 27
rect 3 19 7 21
rect 3 17 4 19
rect 6 17 7 19
rect 3 8 7 17
<< labels >>
rlabel alu1 4 44 4 44 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 40 12 40 6 d
rlabel alu1 20 48 20 48 6 d
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 16 28 16 6 z
rlabel alu1 28 24 28 24 6 b
rlabel alu1 36 32 36 32 6 a
rlabel alu1 36 24 36 24 6 b
rlabel alu1 28 40 28 40 6 c
rlabel alu1 36 52 36 52 6 c
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 20 44 20 6 b
rlabel alu1 44 40 44 40 6 a
<< end >>
