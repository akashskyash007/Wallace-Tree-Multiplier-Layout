magic
tech scmos
timestamp 1199472694
<< ab >>
rect 0 0 40 100
<< nwell >>
rect -5 48 45 105
<< pwell >>
rect -5 -5 45 48
<< alu1 >>
rect -2 95 42 100
rect -2 93 5 95
rect 7 93 14 95
rect 16 93 24 95
rect 26 93 33 95
rect 35 93 42 95
rect -2 88 42 93
rect -2 7 42 12
rect -2 5 5 7
rect 7 5 14 7
rect 16 5 24 7
rect 26 5 33 7
rect 35 5 42 7
rect -2 0 42 5
<< ptie >>
rect 3 7 37 39
rect 3 5 5 7
rect 7 5 14 7
rect 16 5 24 7
rect 26 5 33 7
rect 35 5 37 7
rect 3 3 37 5
<< ntie >>
rect 3 95 37 97
rect 3 93 5 95
rect 7 93 14 95
rect 16 93 24 95
rect 26 93 33 95
rect 35 93 37 95
rect 3 55 37 93
<< ntiect1 >>
rect 5 93 7 95
rect 14 93 16 95
rect 24 93 26 95
rect 33 93 35 95
<< ptiect1 >>
rect 5 5 7 7
rect 14 5 16 7
rect 24 5 26 7
rect 33 5 35 7
<< labels >>
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 94 20 94 6 vdd
<< end >>
