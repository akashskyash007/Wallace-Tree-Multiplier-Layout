magic
tech scmos
timestamp 1199202586
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 10 57 16 59
rect 10 55 12 57
rect 14 55 16 57
rect 10 53 16 55
rect 10 46 12 53
rect 20 46 22 51
rect 10 35 12 38
rect 20 35 22 38
rect 9 32 12 35
rect 16 33 23 35
rect 9 26 11 32
rect 16 31 19 33
rect 21 31 23 33
rect 16 29 23 31
rect 16 26 18 29
rect 9 14 11 19
rect 16 14 18 19
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 19 9 22
rect 11 19 16 26
rect 18 19 27 26
rect 20 16 27 19
rect 20 14 22 16
rect 24 14 27 16
rect 20 12 27 14
<< pdif >>
rect 2 67 8 69
rect 2 65 4 67
rect 6 65 8 67
rect 2 46 8 65
rect 2 38 10 46
rect 12 42 20 46
rect 12 40 15 42
rect 17 40 20 42
rect 12 38 20 40
rect 22 44 30 46
rect 22 42 26 44
rect 28 42 30 44
rect 22 38 30 42
<< alu1 >>
rect -2 67 34 72
rect -2 65 4 67
rect 6 65 17 67
rect 19 65 25 67
rect 27 65 34 67
rect -2 64 34 65
rect 2 57 16 59
rect 2 55 12 57
rect 14 55 16 57
rect 2 54 16 55
rect 2 45 6 54
rect 10 42 19 43
rect 10 40 15 42
rect 17 40 19 42
rect 2 39 19 40
rect 2 36 14 39
rect 2 26 6 36
rect 18 33 30 35
rect 18 31 19 33
rect 21 31 30 33
rect 18 29 30 31
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 20 7 22
rect 26 21 30 29
rect -2 7 34 8
rect -2 5 5 7
rect 7 5 12 7
rect 14 5 34 7
rect -2 0 34 5
<< ptie >>
rect 3 7 16 9
rect 3 5 5 7
rect 7 5 12 7
rect 14 5 16 7
rect 3 3 16 5
<< ntie >>
rect 15 67 29 69
rect 15 65 17 67
rect 19 65 25 67
rect 27 65 29 67
rect 15 63 29 65
<< nmos >>
rect 9 19 11 26
rect 16 19 18 26
<< pmos >>
rect 10 38 12 46
rect 20 38 22 46
<< polyct1 >>
rect 12 55 14 57
rect 19 31 21 33
<< ndifct0 >>
rect 22 14 24 16
<< ndifct1 >>
rect 4 22 6 24
<< ntiect1 >>
rect 17 65 19 67
rect 25 65 27 67
<< ptiect1 >>
rect 5 5 7 7
rect 12 5 14 7
<< pdifct0 >>
rect 26 42 28 44
<< pdifct1 >>
rect 4 65 6 67
rect 15 40 17 42
<< alu0 >>
rect 25 44 29 64
rect 25 42 26 44
rect 28 42 29 44
rect 25 40 29 42
rect 20 16 26 17
rect 20 14 22 16
rect 24 14 26 16
rect 20 8 26 14
<< labels >>
rlabel alu1 4 28 4 28 6 z
rlabel alu1 4 52 4 52 6 b
rlabel alu1 12 40 12 40 6 z
rlabel alu1 12 56 12 56 6 b
rlabel alu1 16 4 16 4 6 vss
rlabel polyct1 20 32 20 32 6 a
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 28 28 28 6 a
<< end >>
