magic
tech scmos
timestamp 1199202417
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 70 11 74
rect 9 39 11 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 30 11 33
rect 9 11 11 16
<< ndif >>
rect 2 27 9 30
rect 2 25 4 27
rect 6 25 9 27
rect 2 20 9 25
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 20 30
rect 13 11 20 16
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 13 71 20 73
rect 13 70 15 71
rect 4 57 9 70
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 48 9 53
rect 2 46 4 48
rect 6 46 9 48
rect 2 44 9 46
rect 4 42 9 44
rect 11 69 15 70
rect 17 69 20 71
rect 11 42 20 69
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 71 26 79
rect -2 69 15 71
rect 17 69 26 71
rect -2 68 26 69
rect 2 57 14 63
rect 2 55 6 57
rect 2 53 4 55
rect 2 48 6 53
rect 2 46 4 48
rect 2 27 6 46
rect 18 39 22 63
rect 10 37 22 39
rect 10 35 11 37
rect 13 35 22 37
rect 10 33 22 35
rect 2 25 4 27
rect 2 23 6 25
rect 2 20 14 23
rect 2 18 4 20
rect 6 18 14 20
rect 2 17 14 18
rect 18 17 22 33
rect -2 11 26 12
rect -2 9 15 11
rect 17 9 26 11
rect -2 1 26 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 16 11 30
<< pmos >>
rect 9 42 11 70
<< polyct1 >>
rect 11 35 13 37
<< ndifct1 >>
rect 4 25 6 27
rect 4 18 6 20
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct1 >>
rect 4 53 6 55
rect 4 46 6 48
rect 15 69 17 71
<< alu0 >>
rect 6 44 7 57
rect 6 23 7 29
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 12 60 12 60 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 40 20 40 6 a
<< end >>
