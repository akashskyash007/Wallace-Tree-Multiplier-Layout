magic
tech scmos
timestamp 1199202148
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 26 69 48 71
rect 56 69 58 74
rect 9 58 11 63
rect 19 58 21 63
rect 26 58 28 69
rect 46 66 48 69
rect 36 58 38 63
rect 9 37 11 42
rect 19 37 21 42
rect 26 39 28 42
rect 36 39 38 42
rect 9 35 21 37
rect 9 32 11 35
rect 5 30 11 32
rect 19 30 21 35
rect 25 37 31 39
rect 25 35 27 37
rect 29 35 31 37
rect 25 33 31 35
rect 36 37 42 39
rect 36 35 38 37
rect 40 35 42 37
rect 36 33 42 35
rect 26 30 28 33
rect 36 30 38 33
rect 46 30 48 50
rect 56 47 58 50
rect 56 45 63 47
rect 56 43 59 45
rect 61 43 63 45
rect 56 41 63 43
rect 56 30 58 41
rect 5 28 7 30
rect 9 28 11 30
rect 5 26 11 28
rect 9 23 11 26
rect 19 18 21 23
rect 26 18 28 23
rect 36 18 38 23
rect 46 18 48 23
rect 9 11 11 16
rect 56 15 58 20
<< ndif >>
rect 13 23 19 30
rect 21 23 26 30
rect 28 28 36 30
rect 28 26 31 28
rect 33 26 36 28
rect 28 23 36 26
rect 38 27 46 30
rect 38 25 41 27
rect 43 25 46 27
rect 38 23 46 25
rect 48 27 56 30
rect 48 25 51 27
rect 53 25 56 27
rect 48 23 56 25
rect 2 20 9 23
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 17 23
rect 50 20 56 23
rect 58 28 65 30
rect 58 26 61 28
rect 63 26 65 28
rect 58 24 65 26
rect 58 20 63 24
rect 13 11 19 16
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 65 19 69
rect 13 58 17 65
rect 50 66 56 69
rect 41 58 46 66
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 4 42 9 45
rect 11 42 19 58
rect 21 42 26 58
rect 28 54 36 58
rect 28 52 31 54
rect 33 52 36 54
rect 28 42 36 52
rect 38 56 46 58
rect 38 54 41 56
rect 43 54 46 56
rect 38 50 46 54
rect 48 64 56 66
rect 48 62 51 64
rect 53 62 56 64
rect 48 50 56 62
rect 58 63 63 69
rect 58 61 65 63
rect 58 59 61 61
rect 63 59 65 61
rect 58 54 65 59
rect 58 52 61 54
rect 63 52 65 54
rect 58 50 65 52
rect 38 42 43 50
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 71 74 79
rect -2 69 15 71
rect 17 69 74 71
rect -2 68 74 69
rect 10 54 35 55
rect 10 52 31 54
rect 33 52 35 54
rect 10 51 35 52
rect 10 49 22 51
rect 2 31 6 39
rect 2 30 14 31
rect 2 28 7 30
rect 9 28 14 30
rect 2 25 14 28
rect 18 29 22 49
rect 26 41 38 47
rect 26 37 30 41
rect 58 45 70 47
rect 58 43 59 45
rect 61 43 70 45
rect 58 41 70 43
rect 26 35 27 37
rect 29 35 30 37
rect 26 33 30 35
rect 66 33 70 41
rect 18 28 35 29
rect 18 26 31 28
rect 33 26 35 28
rect 18 25 35 26
rect -2 11 74 12
rect -2 9 15 11
rect 17 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 19 23 21 30
rect 26 23 28 30
rect 36 23 38 30
rect 46 23 48 30
rect 9 16 11 23
rect 56 20 58 30
<< pmos >>
rect 9 42 11 58
rect 19 42 21 58
rect 26 42 28 58
rect 36 42 38 58
rect 46 50 48 66
rect 56 50 58 69
<< polyct0 >>
rect 38 35 40 37
<< polyct1 >>
rect 27 35 29 37
rect 59 43 61 45
rect 7 28 9 30
<< ndifct0 >>
rect 41 25 43 27
rect 51 25 53 27
rect 4 18 6 20
rect 61 26 63 28
<< ndifct1 >>
rect 31 26 33 28
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 54 6 56
rect 4 47 6 49
rect 41 54 43 56
rect 51 62 53 64
rect 61 59 63 61
rect 61 52 63 54
<< pdifct1 >>
rect 15 69 17 71
rect 31 52 33 54
<< alu0 >>
rect 50 64 54 68
rect 3 59 44 63
rect 50 62 51 64
rect 53 62 54 64
rect 50 60 54 62
rect 60 61 64 63
rect 3 56 7 59
rect 3 54 4 56
rect 6 54 7 56
rect 40 56 44 59
rect 3 49 7 54
rect 40 54 41 56
rect 43 54 44 56
rect 60 59 61 61
rect 63 59 64 61
rect 60 54 64 59
rect 40 52 44 54
rect 50 52 61 54
rect 63 52 64 54
rect 3 47 4 49
rect 6 47 7 49
rect 3 45 7 47
rect 50 50 64 52
rect 50 38 54 50
rect 36 37 62 38
rect 36 35 38 37
rect 40 35 62 37
rect 36 34 62 35
rect 58 29 62 34
rect 40 27 44 29
rect 40 25 41 27
rect 43 25 44 27
rect 40 21 44 25
rect 2 20 44 21
rect 2 18 4 20
rect 6 18 44 20
rect 2 17 44 18
rect 50 27 54 29
rect 50 25 51 27
rect 53 25 54 27
rect 58 28 65 29
rect 58 26 61 28
rect 63 26 65 28
rect 58 25 65 26
rect 50 12 54 25
<< labels >>
rlabel alu0 5 54 5 54 6 n1
rlabel alu0 42 23 42 23 6 n3
rlabel alu0 23 19 23 19 6 n3
rlabel alu0 42 57 42 57 6 n1
rlabel alu0 49 36 49 36 6 cn
rlabel alu0 60 31 60 31 6 cn
rlabel alu0 62 56 62 56 6 cn
rlabel alu1 4 32 4 32 6 a
rlabel alu1 12 28 12 28 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 40 20 40 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 44 36 44 6 b
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 68 40 68 40 6 c
rlabel polyct1 60 44 60 44 6 c
<< end >>
