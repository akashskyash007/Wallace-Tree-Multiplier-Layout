magic
tech scmos
timestamp 1199470322
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -2 48 82 104
<< pwell >>
rect -2 -4 82 48
<< poly >>
rect 25 83 27 88
rect 37 83 39 88
rect 45 83 47 88
rect 57 83 59 88
rect 65 83 67 88
rect 25 52 27 63
rect 25 50 31 52
rect 25 48 27 50
rect 29 48 31 50
rect 12 46 31 48
rect 12 37 14 46
rect 37 43 39 57
rect 45 52 47 57
rect 45 50 53 52
rect 45 48 49 50
rect 51 48 53 50
rect 45 46 53 48
rect 35 41 41 43
rect 35 40 37 41
rect 33 39 37 40
rect 39 39 41 41
rect 33 37 41 39
rect 33 30 35 37
rect 45 30 47 46
rect 57 43 59 57
rect 65 52 67 57
rect 65 50 73 52
rect 65 49 69 50
rect 67 48 69 49
rect 71 48 73 50
rect 67 46 73 48
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 57 30 59 37
rect 67 30 69 46
rect 12 22 14 27
rect 33 13 35 18
rect 45 13 47 18
rect 57 13 59 18
rect 67 13 69 18
<< ndif >>
rect 3 31 12 37
rect 3 29 6 31
rect 8 29 12 31
rect 3 27 12 29
rect 14 35 22 37
rect 14 33 18 35
rect 20 33 22 35
rect 14 31 22 33
rect 14 27 19 31
rect 28 24 33 30
rect 25 22 33 24
rect 25 20 27 22
rect 29 20 33 22
rect 25 18 33 20
rect 35 28 45 30
rect 35 26 39 28
rect 41 26 45 28
rect 35 18 45 26
rect 47 22 57 30
rect 47 20 51 22
rect 53 20 57 22
rect 47 18 57 20
rect 59 18 67 30
rect 69 24 74 30
rect 69 22 77 24
rect 69 20 73 22
rect 75 20 77 22
rect 69 18 77 20
rect 61 11 65 18
rect 61 9 67 11
rect 61 7 63 9
rect 65 7 67 9
rect 61 5 67 7
<< pdif >>
rect 20 77 25 83
rect 17 75 25 77
rect 17 73 19 75
rect 21 73 25 75
rect 17 67 25 73
rect 17 65 19 67
rect 21 65 25 67
rect 17 63 25 65
rect 27 81 37 83
rect 27 79 31 81
rect 33 79 37 81
rect 27 63 37 79
rect 29 57 37 63
rect 39 57 45 83
rect 47 81 57 83
rect 47 79 51 81
rect 53 79 57 81
rect 47 73 57 79
rect 47 71 51 73
rect 53 71 57 73
rect 47 57 57 71
rect 59 57 65 83
rect 67 81 76 83
rect 67 79 71 81
rect 73 79 76 81
rect 67 57 76 79
<< alu1 >>
rect -2 95 82 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 82 95
rect -2 88 82 93
rect 18 75 22 83
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 77 34 79
rect 50 81 54 83
rect 50 79 51 81
rect 53 79 54 81
rect 18 73 19 75
rect 21 73 22 75
rect 18 67 22 73
rect 50 73 54 79
rect 70 81 74 88
rect 70 79 71 81
rect 73 79 74 81
rect 70 77 74 79
rect 50 72 51 73
rect 18 65 19 67
rect 21 65 22 67
rect 18 42 22 65
rect 28 71 51 72
rect 53 71 54 73
rect 28 68 54 71
rect 28 52 32 68
rect 58 67 72 73
rect 26 50 32 52
rect 26 48 27 50
rect 29 48 32 50
rect 26 46 32 48
rect 7 38 22 42
rect 17 35 22 38
rect 17 33 18 35
rect 20 33 22 35
rect 5 31 9 33
rect 5 29 6 31
rect 8 29 9 31
rect 5 12 9 29
rect 17 27 22 33
rect 28 32 32 46
rect 38 58 53 63
rect 38 43 42 58
rect 36 41 42 43
rect 36 39 37 41
rect 39 39 42 41
rect 36 37 42 39
rect 48 50 52 53
rect 48 48 49 50
rect 51 48 52 50
rect 48 32 52 48
rect 57 42 62 63
rect 68 50 72 67
rect 68 48 69 50
rect 71 48 72 50
rect 68 46 72 48
rect 57 41 73 42
rect 57 39 59 41
rect 61 39 73 41
rect 57 38 73 39
rect 28 28 43 32
rect 37 26 39 28
rect 41 26 43 28
rect 48 27 63 32
rect 37 25 43 26
rect 25 22 31 23
rect 25 20 27 22
rect 29 21 31 22
rect 49 22 55 23
rect 49 21 51 22
rect 29 20 51 21
rect 53 21 55 22
rect 71 22 77 23
rect 71 21 73 22
rect 53 20 73 21
rect 75 20 77 22
rect 25 17 77 20
rect -2 9 82 12
rect -2 7 63 9
rect 65 7 82 9
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 82 7
rect -2 0 82 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 12 27 14 37
rect 33 18 35 30
rect 45 18 47 30
rect 57 18 59 30
rect 67 18 69 30
<< pmos >>
rect 25 63 27 83
rect 37 57 39 83
rect 45 57 47 83
rect 57 57 59 83
rect 65 57 67 83
<< polyct1 >>
rect 27 48 29 50
rect 49 48 51 50
rect 37 39 39 41
rect 69 48 71 50
rect 59 39 61 41
<< ndifct1 >>
rect 6 29 8 31
rect 18 33 20 35
rect 27 20 29 22
rect 39 26 41 28
rect 51 20 53 22
rect 73 20 75 22
rect 63 7 65 9
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 19 73 21 75
rect 19 65 21 67
rect 31 79 33 81
rect 51 79 53 81
rect 51 71 53 73
rect 71 79 73 81
<< labels >>
rlabel alu1 10 40 10 40 6 z
rlabel alu1 20 55 20 55 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 40 28 40 28 6 zn
rlabel alu1 40 50 40 50 6 b1
rlabel alu1 30 50 30 50 6 zn
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 60 30 60 30 6 b2
rlabel alu1 50 40 50 40 6 b2
rlabel alu1 60 50 60 50 6 a2
rlabel alu1 50 60 50 60 6 b1
rlabel alu1 60 70 60 70 6 a1
rlabel alu1 52 75 52 75 6 zn
rlabel alu1 51 19 51 19 6 n3
rlabel alu1 70 40 70 40 6 a2
rlabel alu1 70 60 70 60 6 a1
<< end >>
