magic
tech scmos
timestamp 1199202964
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 70 48 74
rect 53 70 55 74
rect 12 39 14 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 15 39
rect 19 37 31 39
rect 36 39 38 42
rect 46 39 48 42
rect 53 39 55 42
rect 36 37 48 39
rect 52 37 58 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 22 35 24 37
rect 26 35 28 37
rect 22 33 28 35
rect 36 35 38 37
rect 40 35 44 37
rect 36 33 44 35
rect 13 30 15 33
rect 23 30 25 33
rect 42 30 44 33
rect 52 35 54 37
rect 56 35 58 37
rect 52 33 58 35
rect 52 30 54 33
rect 13 6 15 10
rect 23 6 25 10
rect 42 6 44 10
rect 52 6 54 10
<< ndif >>
rect 5 14 13 30
rect 5 12 8 14
rect 10 12 13 14
rect 5 10 13 12
rect 15 21 23 30
rect 15 19 18 21
rect 20 19 23 21
rect 15 10 23 19
rect 25 14 42 30
rect 25 12 33 14
rect 35 12 42 14
rect 25 10 42 12
rect 44 28 52 30
rect 44 26 47 28
rect 49 26 52 28
rect 44 21 52 26
rect 44 19 47 21
rect 49 19 52 21
rect 44 10 52 19
rect 54 21 62 30
rect 54 19 58 21
rect 60 19 62 21
rect 54 14 62 19
rect 54 12 58 14
rect 60 12 62 14
rect 54 10 62 12
<< pdif >>
rect 7 55 12 70
rect 5 53 12 55
rect 5 51 7 53
rect 9 51 12 53
rect 5 46 12 51
rect 5 44 7 46
rect 9 44 12 46
rect 5 42 12 44
rect 14 42 19 70
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 42 36 70
rect 38 61 46 70
rect 38 59 41 61
rect 43 59 46 61
rect 38 54 46 59
rect 38 52 41 54
rect 43 52 46 54
rect 38 42 46 52
rect 48 42 53 70
rect 55 68 62 70
rect 55 66 58 68
rect 60 66 62 68
rect 55 61 62 66
rect 55 59 58 61
rect 60 59 62 61
rect 55 42 62 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 40 61 46 63
rect 40 59 41 61
rect 43 59 46 61
rect 40 54 46 59
rect 5 53 41 54
rect 5 51 7 53
rect 9 52 41 53
rect 43 52 46 54
rect 9 51 46 52
rect 5 50 46 51
rect 5 47 11 50
rect 2 46 11 47
rect 2 44 7 46
rect 9 44 11 46
rect 2 43 11 44
rect 2 22 6 43
rect 22 42 55 46
rect 10 37 18 39
rect 10 35 11 37
rect 13 35 18 37
rect 10 33 18 35
rect 22 37 28 42
rect 49 38 55 42
rect 22 35 24 37
rect 26 35 28 37
rect 22 34 28 35
rect 33 37 42 38
rect 33 35 38 37
rect 40 35 42 37
rect 33 34 42 35
rect 49 37 58 38
rect 49 35 54 37
rect 56 35 58 37
rect 49 34 58 35
rect 14 30 18 33
rect 33 30 39 34
rect 14 26 39 30
rect 46 28 51 30
rect 46 26 47 28
rect 49 26 51 28
rect 46 22 51 26
rect 2 21 51 22
rect 2 19 18 21
rect 20 19 47 21
rect 49 19 51 21
rect 2 18 51 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 13 10 15 30
rect 23 10 25 30
rect 42 10 44 30
rect 52 10 54 30
<< pmos >>
rect 12 42 14 70
rect 19 42 21 70
rect 29 42 31 70
rect 36 42 38 70
rect 46 42 48 70
rect 53 42 55 70
<< polyct1 >>
rect 11 35 13 37
rect 24 35 26 37
rect 38 35 40 37
rect 54 35 56 37
<< ndifct0 >>
rect 8 12 10 14
rect 33 12 35 14
rect 58 19 60 21
rect 58 12 60 14
<< ndifct1 >>
rect 18 19 20 21
rect 47 26 49 28
rect 47 19 49 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 24 66 26 68
rect 24 59 26 61
rect 58 66 60 68
rect 58 59 60 61
<< pdifct1 >>
rect 7 51 9 53
rect 7 44 9 46
rect 41 59 43 61
rect 41 52 43 54
<< alu0 >>
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 56 66 58 68
rect 60 66 62 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 56 61 62 66
rect 56 59 58 61
rect 60 59 62 61
rect 56 58 62 59
rect 57 21 61 23
rect 57 19 58 21
rect 60 19 61 21
rect 6 14 12 15
rect 6 12 8 14
rect 10 12 12 14
rect 31 14 37 15
rect 31 12 33 14
rect 35 12 37 14
rect 57 14 61 19
rect 57 12 58 14
rect 60 12 61 14
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 b
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 44 28 44 6 a
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 32 36 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 40 52 40 6 a
<< end >>
