magic
tech scmos
timestamp 1199980682
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -8 40 72 97
<< pwell >>
rect -8 -9 72 40
<< poly >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 84 46 86
rect 37 82 42 84
rect 44 82 46 84
rect 37 80 46 82
rect 50 84 59 86
rect 50 82 52 84
rect 54 82 59 84
rect 50 80 59 82
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 42 43 48
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 2 32 17 38
rect 21 32 30 38
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 6 27 8
rect 18 4 23 6
rect 25 4 27 6
rect 18 2 27 4
rect 37 2 46 8
rect 50 2 59 8
<< ndif >>
rect 2 11 9 29
rect 11 15 21 29
rect 11 13 15 15
rect 17 13 21 15
rect 11 11 21 13
rect 23 11 30 29
rect 34 23 41 29
rect 34 21 36 23
rect 38 21 41 23
rect 34 16 41 21
rect 34 14 36 16
rect 38 14 41 16
rect 34 11 41 14
rect 43 25 53 29
rect 43 23 47 25
rect 49 23 53 25
rect 43 17 53 23
rect 43 15 47 17
rect 49 15 53 17
rect 43 11 53 15
rect 55 23 62 29
rect 55 21 58 23
rect 60 21 62 23
rect 55 16 62 21
rect 55 14 58 16
rect 60 14 62 16
rect 55 11 62 14
<< pdif >>
rect 2 74 9 77
rect 2 72 4 74
rect 6 72 9 74
rect 2 67 9 72
rect 2 65 4 67
rect 6 65 9 67
rect 2 51 9 65
rect 11 68 21 77
rect 11 66 15 68
rect 17 66 21 68
rect 11 61 21 66
rect 11 59 15 61
rect 17 59 21 61
rect 11 51 21 59
rect 23 75 30 77
rect 23 73 26 75
rect 28 73 30 75
rect 23 68 30 73
rect 23 66 26 68
rect 28 66 30 68
rect 23 51 30 66
rect 34 74 41 77
rect 34 72 36 74
rect 38 72 41 74
rect 34 61 41 72
rect 34 59 36 61
rect 38 59 41 61
rect 34 51 41 59
rect 43 65 53 77
rect 43 63 47 65
rect 49 63 53 65
rect 43 57 53 63
rect 43 55 47 57
rect 49 55 53 57
rect 43 51 53 55
rect 55 74 62 77
rect 55 72 58 74
rect 60 72 62 74
rect 55 67 62 72
rect 55 65 58 67
rect 60 65 62 67
rect 55 51 62 65
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect 62 85 66 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 81 34 83
rect 62 83 63 85
rect 65 83 66 85
rect 62 81 66 83
rect 3 74 7 81
rect 3 72 4 74
rect 6 72 7 74
rect 3 67 7 72
rect 25 75 29 81
rect 25 73 26 75
rect 28 73 29 75
rect 3 65 4 67
rect 6 65 7 67
rect 3 63 7 65
rect 25 68 29 73
rect 25 66 26 68
rect 28 66 29 68
rect 25 64 29 66
rect 46 65 50 67
rect 46 63 47 65
rect 49 63 50 65
rect 46 57 50 63
rect 46 55 47 57
rect 49 55 50 57
rect 5 46 26 50
rect 5 44 7 46
rect 9 44 11 46
rect 5 43 11 44
rect 22 44 23 46
rect 25 44 26 46
rect 22 34 26 44
rect 38 36 42 38
rect 38 34 39 36
rect 41 34 42 36
rect 22 30 42 34
rect 46 25 50 55
rect 54 46 58 59
rect 54 44 55 46
rect 57 44 58 46
rect 54 36 58 44
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 35 23 39 25
rect 35 21 36 23
rect 38 21 39 23
rect 14 15 18 17
rect 14 13 15 15
rect 17 13 18 15
rect 14 7 18 13
rect 35 16 39 21
rect 35 14 36 16
rect 38 14 39 16
rect 35 7 39 14
rect 46 23 47 25
rect 49 23 50 25
rect 46 17 50 23
rect 46 15 47 17
rect 49 15 50 17
rect 46 13 50 15
rect 57 23 61 25
rect 57 21 58 23
rect 60 21 61 23
rect 57 16 61 21
rect 57 14 58 16
rect 60 14 61 16
rect -2 6 39 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 4 23 6
rect 25 5 39 6
rect 25 4 31 5
rect 1 3 31 4
rect 33 3 39 5
rect 57 7 61 14
rect 57 5 66 7
rect 57 3 63 5
rect 65 3 66 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 -2 66 3
<< alu2 >>
rect -2 85 66 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 66 85
rect -2 80 66 83
rect -2 5 66 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 66 5
rect -2 -2 66 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polyct0 >>
rect 42 82 44 84
rect 52 82 54 84
<< polyct1 >>
rect 7 44 9 46
rect 23 44 25 46
rect 55 44 57 46
rect 39 34 41 36
rect 55 34 57 36
rect 7 4 9 6
rect 23 4 25 6
<< ndifct1 >>
rect 15 13 17 15
rect 36 21 38 23
rect 36 14 38 16
rect 47 23 49 25
rect 47 15 49 17
rect 58 21 60 23
rect 58 14 60 16
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< pdifct0 >>
rect 15 66 17 68
rect 15 59 17 61
rect 36 72 38 74
rect 36 59 38 61
rect 58 72 60 74
rect 58 65 60 67
<< pdifct1 >>
rect 4 72 6 74
rect 4 65 6 67
rect 26 73 28 75
rect 26 66 28 68
rect 47 63 49 65
rect 47 55 49 57
<< alu0 >>
rect 40 84 56 85
rect 40 82 42 84
rect 44 82 52 84
rect 54 82 56 84
rect 40 81 56 82
rect 14 68 18 70
rect 14 66 15 68
rect 17 66 18 68
rect 14 61 18 66
rect 35 74 61 76
rect 35 72 36 74
rect 38 72 58 74
rect 60 72 61 74
rect 35 61 39 72
rect 57 67 61 72
rect 14 59 15 61
rect 17 59 36 61
rect 38 59 39 61
rect 14 57 39 59
rect 57 65 58 67
rect 60 65 61 67
rect 57 63 61 65
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< labels >>
rlabel alu1 8 48 8 48 6 a
rlabel alu1 24 40 24 40 6 a
rlabel alu1 16 48 16 48 6 a
rlabel alu1 32 32 32 32 6 a
rlabel alu1 48 40 48 40 6 z
rlabel alu1 56 48 56 48 6 b
rlabel via1 32 4 32 4 6 vss
rlabel via1 32 84 32 84 6 vdd
<< end >>
