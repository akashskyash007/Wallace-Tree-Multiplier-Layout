magic
tech scmos
timestamp 1199201754
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 20 61 22 66
rect 30 61 32 66
rect 42 61 44 66
rect 52 61 54 66
rect 9 57 11 61
rect 9 35 11 39
rect 20 35 22 48
rect 30 45 32 48
rect 30 43 37 45
rect 30 41 33 43
rect 35 41 37 43
rect 30 39 37 41
rect 42 43 44 48
rect 42 41 48 43
rect 42 39 44 41
rect 46 39 48 41
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 20 33 26 35
rect 20 31 22 33
rect 24 31 26 33
rect 20 29 26 31
rect 9 24 11 29
rect 24 24 26 29
rect 31 24 33 39
rect 42 37 48 39
rect 42 35 44 37
rect 38 33 44 35
rect 52 35 54 48
rect 52 33 58 35
rect 38 24 40 33
rect 52 31 54 33
rect 56 31 58 33
rect 52 29 58 31
rect 45 27 58 29
rect 45 24 47 27
rect 9 11 11 15
rect 24 3 26 8
rect 31 3 33 8
rect 38 3 40 8
rect 45 3 47 8
<< ndif >>
rect 4 21 9 24
rect 2 19 9 21
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 15 24 24
rect 13 8 24 15
rect 26 8 31 24
rect 33 8 38 24
rect 40 8 45 24
rect 47 18 52 24
rect 47 16 54 18
rect 47 14 50 16
rect 52 14 54 16
rect 47 12 54 14
rect 47 8 52 12
rect 13 7 22 8
rect 13 5 16 7
rect 18 5 22 7
rect 13 3 22 5
<< pdif >>
rect 34 67 40 69
rect 34 65 36 67
rect 38 65 40 67
rect 34 61 40 65
rect 13 58 20 61
rect 13 57 15 58
rect 4 52 9 57
rect 2 50 9 52
rect 2 48 4 50
rect 6 48 9 50
rect 2 43 9 48
rect 2 41 4 43
rect 6 41 9 43
rect 2 39 9 41
rect 11 56 15 57
rect 17 56 20 58
rect 11 48 20 56
rect 22 58 30 61
rect 22 56 25 58
rect 27 56 30 58
rect 22 48 30 56
rect 32 48 42 61
rect 44 58 52 61
rect 44 56 47 58
rect 49 56 52 58
rect 44 48 52 56
rect 54 59 61 61
rect 54 57 57 59
rect 59 57 61 59
rect 54 52 61 57
rect 54 50 57 52
rect 59 50 61 52
rect 54 48 61 50
rect 11 39 18 48
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 36 67
rect 38 65 66 67
rect -2 64 66 65
rect 2 50 7 59
rect 2 48 4 50
rect 6 48 7 50
rect 2 43 7 48
rect 2 41 4 43
rect 6 41 7 43
rect 2 39 7 41
rect 2 19 6 39
rect 34 43 38 51
rect 25 41 33 42
rect 35 41 38 43
rect 25 38 38 41
rect 42 42 46 51
rect 42 41 55 42
rect 42 39 44 41
rect 46 39 55 41
rect 42 38 55 39
rect 20 33 31 34
rect 20 31 22 33
rect 24 31 31 33
rect 20 30 31 31
rect 41 33 62 34
rect 41 31 54 33
rect 56 31 62 33
rect 41 30 62 31
rect 27 26 31 30
rect 27 22 47 26
rect 2 17 4 19
rect 6 17 15 18
rect 2 13 15 17
rect 58 13 62 30
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 16 7
rect 18 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 15 11 24
rect 24 8 26 24
rect 31 8 33 24
rect 38 8 40 24
rect 45 8 47 24
<< pmos >>
rect 9 39 11 57
rect 20 48 22 61
rect 30 48 32 61
rect 42 48 44 61
rect 52 48 54 61
<< polyct0 >>
rect 33 42 34 43
rect 11 31 13 33
<< polyct1 >>
rect 34 42 35 43
rect 33 41 35 42
rect 44 39 46 41
rect 22 31 24 33
rect 54 31 56 33
<< ndifct0 >>
rect 50 14 52 16
<< ndifct1 >>
rect 4 17 6 19
rect 16 5 18 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 15 56 17 58
rect 25 56 27 58
rect 47 56 49 58
rect 57 57 59 59
rect 57 50 59 52
<< pdifct1 >>
rect 36 65 38 67
rect 4 48 6 50
rect 4 41 6 43
<< alu0 >>
rect 14 58 18 64
rect 56 59 60 64
rect 14 56 15 58
rect 17 56 18 58
rect 14 54 18 56
rect 22 58 51 59
rect 22 56 25 58
rect 27 56 47 58
rect 49 56 51 58
rect 22 55 51 56
rect 56 57 57 59
rect 59 57 60 59
rect 22 50 26 55
rect 56 52 60 57
rect 12 46 26 50
rect 12 35 16 46
rect 32 43 34 44
rect 32 42 33 43
rect 56 50 57 52
rect 59 50 60 52
rect 56 48 60 50
rect 10 33 16 35
rect 10 31 11 33
rect 13 31 16 33
rect 10 29 16 31
rect 12 26 16 29
rect 12 22 23 26
rect 6 18 7 21
rect 19 17 23 22
rect 19 16 54 17
rect 19 14 50 16
rect 52 14 54 16
rect 19 13 54 14
<< labels >>
rlabel alu0 14 36 14 36 6 zn
rlabel alu0 36 15 36 15 6 zn
rlabel alu0 36 57 36 57 6 zn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 44 32 44 32 6 d
rlabel alu1 36 48 36 48 6 b
rlabel alu1 44 48 44 48 6 c
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 60 20 60 20 6 d
rlabel alu1 52 32 52 32 6 d
rlabel alu1 52 40 52 40 6 c
<< end >>
