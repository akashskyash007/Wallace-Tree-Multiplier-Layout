magic
tech scmos
timestamp 1199980685
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -8 40 72 97
<< pwell >>
rect -8 -9 72 40
<< poly >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 2 32 17 38
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 32 62 38
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 2 27 8
rect 37 2 46 8
rect 50 6 59 8
rect 50 4 55 6
rect 57 4 59 6
rect 50 2 59 4
<< ndif >>
rect 2 11 9 29
rect 11 23 21 29
rect 11 21 15 23
rect 17 21 21 23
rect 11 15 21 21
rect 11 13 15 15
rect 17 13 21 15
rect 11 11 21 13
rect 23 25 30 29
rect 23 23 26 25
rect 28 23 30 25
rect 23 17 30 23
rect 23 15 26 17
rect 28 15 30 17
rect 23 11 30 15
rect 34 25 41 29
rect 34 23 36 25
rect 38 23 41 25
rect 34 17 41 23
rect 34 15 36 17
rect 38 15 41 17
rect 34 11 41 15
rect 43 23 53 29
rect 43 21 47 23
rect 49 21 53 23
rect 43 16 53 21
rect 43 14 47 16
rect 49 14 53 16
rect 43 11 53 14
rect 55 11 62 29
<< pdif >>
rect 2 74 9 77
rect 2 72 4 74
rect 6 72 9 74
rect 2 67 9 72
rect 2 65 4 67
rect 6 65 9 67
rect 2 51 9 65
rect 11 65 21 77
rect 11 63 15 65
rect 17 63 21 65
rect 11 58 21 63
rect 11 56 15 58
rect 17 56 21 58
rect 11 51 21 56
rect 23 74 30 77
rect 23 72 26 74
rect 28 72 30 74
rect 23 51 30 72
rect 34 74 41 77
rect 34 72 36 74
rect 38 72 41 74
rect 34 67 41 72
rect 34 65 36 67
rect 38 65 41 67
rect 34 51 41 65
rect 43 65 53 77
rect 43 63 47 65
rect 49 63 53 65
rect 43 57 53 63
rect 43 55 47 57
rect 49 55 53 57
rect 43 51 53 55
rect 55 74 62 77
rect 55 72 58 74
rect 60 72 62 74
rect 55 67 62 72
rect 55 65 58 67
rect 60 65 62 67
rect 55 51 62 65
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 81 34 83
rect 62 85 66 90
rect 62 83 63 85
rect 65 83 66 85
rect 62 81 66 83
rect 46 65 50 67
rect 46 63 47 65
rect 49 63 50 65
rect 46 59 50 63
rect 22 50 26 59
rect 5 46 26 50
rect 5 44 7 46
rect 9 44 11 46
rect 5 43 11 44
rect 22 44 23 46
rect 25 44 26 46
rect 22 36 26 44
rect 22 34 23 36
rect 25 34 26 36
rect 22 32 26 34
rect 30 57 50 59
rect 30 55 47 57
rect 49 55 50 57
rect 30 26 34 55
rect 46 53 50 55
rect 38 46 42 51
rect 38 44 39 46
rect 41 44 42 46
rect 38 42 42 44
rect 53 46 59 47
rect 53 44 55 46
rect 57 44 59 46
rect 53 42 59 44
rect 38 38 59 42
rect 38 36 42 38
rect 38 34 39 36
rect 41 34 42 36
rect 38 29 42 34
rect 24 25 34 26
rect 24 23 26 25
rect 28 23 34 25
rect 24 22 34 23
rect 30 18 34 22
rect 24 17 40 18
rect 24 15 26 17
rect 28 15 36 17
rect 38 15 40 17
rect 24 14 40 15
rect -2 6 66 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 5 55 6
rect 9 4 31 5
rect 1 3 31 4
rect 33 4 55 5
rect 57 5 66 6
rect 57 4 63 5
rect 33 3 63 4
rect 65 3 66 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 -2 66 3
<< alu2 >>
rect -2 85 66 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 66 85
rect -2 80 66 83
rect -2 5 66 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 66 5
rect -2 -2 66 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polyct1 >>
rect 7 44 9 46
rect 23 44 25 46
rect 39 44 41 46
rect 55 44 57 46
rect 23 34 25 36
rect 39 34 41 36
rect 7 4 9 6
rect 55 4 57 6
<< ndifct0 >>
rect 15 21 17 23
rect 15 13 17 15
rect 36 23 38 25
rect 47 21 49 23
rect 47 14 49 16
<< ndifct1 >>
rect 26 23 28 25
rect 26 15 28 17
rect 36 15 38 17
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< pdifct0 >>
rect 4 72 6 74
rect 4 65 6 67
rect 15 63 17 65
rect 15 56 17 58
rect 26 72 28 74
rect 36 72 38 74
rect 36 65 38 67
rect 58 72 60 74
rect 58 65 60 67
<< pdifct1 >>
rect 47 63 49 65
rect 47 55 49 57
<< alu0 >>
rect 3 74 7 81
rect 3 72 4 74
rect 6 72 7 74
rect 3 67 7 72
rect 25 74 29 81
rect 25 72 26 74
rect 28 72 29 74
rect 25 70 29 72
rect 35 74 61 76
rect 35 72 36 74
rect 38 72 58 74
rect 60 72 61 74
rect 35 67 39 72
rect 57 67 61 72
rect 3 65 4 67
rect 6 65 7 67
rect 3 63 7 65
rect 14 65 36 67
rect 38 65 39 67
rect 14 63 15 65
rect 17 63 39 65
rect 57 65 58 67
rect 60 65 61 67
rect 57 63 61 65
rect 14 58 18 63
rect 14 56 15 58
rect 17 56 18 58
rect 14 54 18 56
rect 34 25 40 26
rect 14 23 18 25
rect 14 21 15 23
rect 17 21 18 23
rect 34 23 36 25
rect 38 23 40 25
rect 34 22 40 23
rect 46 23 50 25
rect 14 15 18 21
rect 46 21 47 23
rect 49 21 50 23
rect 14 13 15 15
rect 17 13 18 15
rect 46 16 50 21
rect 46 14 47 16
rect 49 14 50 16
rect 14 7 18 13
rect 46 7 50 14
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< labels >>
rlabel alu1 8 48 8 48 6 a
rlabel alu1 24 48 24 48 6 a
rlabel alu1 16 48 16 48 6 a
rlabel alu1 32 36 32 36 6 z
rlabel alu1 40 40 40 40 6 b
rlabel alu1 48 40 48 40 6 b
rlabel alu1 56 40 56 40 6 b
rlabel alu1 48 60 48 60 6 z
rlabel via1 32 4 32 4 6 vss
rlabel via1 32 84 32 84 6 vdd
<< end >>
