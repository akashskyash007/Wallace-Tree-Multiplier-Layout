magic
tech scmos
timestamp 1199203330
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 28 62 30 67
rect 35 62 37 67
rect 42 62 44 67
rect 49 62 51 67
rect 9 55 11 60
rect 28 47 30 50
rect 19 45 30 47
rect 19 43 21 45
rect 23 43 25 45
rect 9 40 11 43
rect 19 41 25 43
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 9 30 11 34
rect 19 30 21 41
rect 35 39 37 50
rect 29 37 37 39
rect 29 35 31 37
rect 33 36 37 37
rect 33 35 35 36
rect 29 33 35 35
rect 29 30 31 33
rect 42 31 44 50
rect 49 47 51 50
rect 49 45 55 47
rect 49 43 51 45
rect 53 43 55 45
rect 49 41 55 43
rect 9 19 11 24
rect 19 19 21 24
rect 29 19 31 24
rect 39 29 45 31
rect 39 27 41 29
rect 43 27 45 29
rect 39 25 45 27
rect 39 22 41 25
rect 49 22 51 41
rect 39 11 41 16
rect 49 11 51 16
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 11 24 19 30
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 24 29 26
rect 31 24 37 30
rect 13 17 17 24
rect 33 22 37 24
rect 33 17 39 22
rect 13 15 19 17
rect 13 13 15 15
rect 17 13 19 15
rect 13 11 19 13
rect 31 16 39 17
rect 41 20 49 22
rect 41 18 44 20
rect 46 18 49 20
rect 41 16 49 18
rect 51 16 59 22
rect 31 11 37 16
rect 53 11 59 16
rect 31 9 33 11
rect 35 9 37 11
rect 31 7 37 9
rect 53 9 55 11
rect 57 9 59 11
rect 53 7 59 9
<< pdif >>
rect 53 71 59 73
rect 53 69 55 71
rect 57 69 59 71
rect 13 64 19 66
rect 13 62 15 64
rect 17 62 19 64
rect 53 62 59 69
rect 13 60 19 62
rect 13 55 17 60
rect 23 56 28 62
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 49 9 51
rect 4 43 9 49
rect 11 43 17 55
rect 21 54 28 56
rect 21 52 23 54
rect 25 52 28 54
rect 21 50 28 52
rect 30 50 35 62
rect 37 50 42 62
rect 44 50 49 62
rect 51 50 59 62
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 55 71
rect 57 69 66 71
rect -2 68 66 69
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 49 7 51
rect 2 30 6 49
rect 34 46 38 63
rect 42 57 54 63
rect 17 45 38 46
rect 17 43 21 45
rect 23 43 38 45
rect 17 42 38 43
rect 42 38 46 47
rect 50 45 54 57
rect 50 43 51 45
rect 53 43 54 45
rect 50 41 54 43
rect 29 37 46 38
rect 29 35 31 37
rect 33 35 46 37
rect 29 34 46 35
rect 2 28 16 30
rect 2 26 4 28
rect 6 26 16 28
rect 2 25 16 26
rect 39 29 62 30
rect 39 27 41 29
rect 43 27 62 29
rect 39 26 62 27
rect 58 17 62 26
rect -2 11 66 12
rect -2 9 33 11
rect 35 9 55 11
rect 57 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 24 11 30
rect 19 24 21 30
rect 29 24 31 30
rect 39 16 41 22
rect 49 16 51 22
<< pmos >>
rect 9 43 11 55
rect 28 50 30 62
rect 35 50 37 62
rect 42 50 44 62
rect 49 50 51 62
<< polyct0 >>
rect 11 36 13 38
<< polyct1 >>
rect 21 43 23 45
rect 31 35 33 37
rect 51 43 53 45
rect 41 27 43 29
<< ndifct0 >>
rect 24 26 26 28
rect 15 13 17 15
rect 44 18 46 20
<< ndifct1 >>
rect 4 26 6 28
rect 33 9 35 11
rect 55 9 57 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 15 62 17 64
rect 23 52 25 54
<< pdifct1 >>
rect 55 69 57 71
rect 4 51 6 53
<< alu0 >>
rect 14 64 18 68
rect 14 62 15 64
rect 17 62 18 64
rect 14 60 18 62
rect 10 54 27 55
rect 10 52 23 54
rect 25 52 27 54
rect 10 51 27 52
rect 10 38 14 51
rect 10 36 11 38
rect 13 36 25 38
rect 10 34 25 36
rect 21 29 25 34
rect 21 28 29 29
rect 21 26 24 28
rect 26 26 29 28
rect 21 25 29 26
rect 25 21 29 25
rect 25 20 48 21
rect 25 18 44 20
rect 46 18 48 20
rect 25 17 48 18
rect 14 15 18 17
rect 14 13 15 15
rect 17 13 18 15
rect 14 12 18 13
<< labels >>
rlabel alu0 12 44 12 44 6 zn
rlabel alu0 18 53 18 53 6 zn
rlabel alu0 36 19 36 19 6 zn
rlabel alu1 12 28 12 28 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 44 20 44 6 d
rlabel alu1 28 44 28 44 6 d
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 36 36 36 6 c
rlabel alu1 44 28 44 28 6 b
rlabel alu1 44 44 44 44 6 c
rlabel alu1 36 56 36 56 6 d
rlabel alu1 44 60 44 60 6 a
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 60 20 60 20 6 b
rlabel alu1 52 28 52 28 6 b
rlabel alu1 52 52 52 52 6 a
<< end >>
