magic
tech scmos
timestamp 1199203162
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 52 70 54 74
rect 59 70 61 74
rect 69 70 71 74
rect 76 70 78 74
rect 12 39 14 42
rect 19 39 21 42
rect 29 39 31 42
rect 36 39 38 42
rect 52 39 54 42
rect 59 39 61 42
rect 69 39 71 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 24 37
rect 26 35 31 37
rect 19 33 31 35
rect 35 37 41 39
rect 35 35 37 37
rect 39 35 41 37
rect 35 33 41 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 33
rect 49 37 55 39
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 59 37 71 39
rect 76 39 78 42
rect 76 37 87 39
rect 59 35 67 37
rect 69 35 71 37
rect 59 33 71 35
rect 49 30 51 33
rect 59 30 61 33
rect 69 30 71 33
rect 81 35 83 37
rect 85 35 87 37
rect 81 33 87 35
rect 81 30 83 33
rect 69 16 71 21
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 39 11 41 16
rect 49 11 51 16
rect 59 11 61 16
rect 81 16 83 21
<< ndif >>
rect 4 22 9 30
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 16 19 26
rect 21 20 29 30
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 16 39 26
rect 41 27 49 30
rect 41 25 44 27
rect 46 25 49 27
rect 41 20 49 25
rect 41 18 44 20
rect 46 18 49 20
rect 41 16 49 18
rect 51 20 59 30
rect 51 18 54 20
rect 56 18 59 20
rect 51 16 59 18
rect 61 28 69 30
rect 61 26 64 28
rect 66 26 69 28
rect 61 21 69 26
rect 71 21 81 30
rect 83 27 88 30
rect 83 25 90 27
rect 83 23 86 25
rect 88 23 90 25
rect 83 21 90 23
rect 61 16 66 21
rect 73 11 79 21
rect 73 9 75 11
rect 77 9 79 11
rect 73 7 79 9
<< pdif >>
rect 4 68 12 70
rect 4 66 7 68
rect 9 66 12 68
rect 4 61 12 66
rect 4 59 7 61
rect 9 59 12 61
rect 4 42 12 59
rect 14 42 19 70
rect 21 61 29 70
rect 21 59 24 61
rect 26 59 29 61
rect 21 54 29 59
rect 21 52 24 54
rect 26 52 29 54
rect 21 42 29 52
rect 31 42 36 70
rect 38 68 52 70
rect 38 66 45 68
rect 47 66 52 68
rect 38 61 52 66
rect 38 59 45 61
rect 47 59 52 61
rect 38 42 52 59
rect 54 42 59 70
rect 61 61 69 70
rect 61 59 64 61
rect 66 59 69 61
rect 61 54 69 59
rect 61 52 64 54
rect 66 52 69 54
rect 61 42 69 52
rect 71 42 76 70
rect 78 63 83 70
rect 78 61 88 63
rect 78 59 83 61
rect 85 59 88 61
rect 78 54 88 59
rect 78 52 83 54
rect 85 52 88 54
rect 78 42 88 52
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 63 61 70 63
rect 63 59 64 61
rect 66 59 70 61
rect 63 57 70 59
rect 63 54 67 57
rect 2 52 24 54
rect 26 52 64 54
rect 66 52 67 54
rect 2 50 67 52
rect 2 29 6 50
rect 74 46 78 55
rect 12 42 40 46
rect 36 39 40 42
rect 50 42 86 46
rect 17 37 31 38
rect 17 35 24 37
rect 26 35 31 37
rect 17 34 31 35
rect 36 37 46 39
rect 36 35 37 37
rect 39 35 46 37
rect 36 33 46 35
rect 50 37 54 42
rect 50 35 51 37
rect 53 35 54 37
rect 50 33 54 35
rect 65 37 78 38
rect 65 35 67 37
rect 69 35 78 37
rect 65 34 78 35
rect 2 28 38 29
rect 2 26 14 28
rect 16 26 34 28
rect 36 26 38 28
rect 2 25 38 26
rect 74 25 78 34
rect 82 37 86 42
rect 82 35 83 37
rect 85 35 86 37
rect 82 33 86 35
rect -2 11 98 12
rect -2 9 75 11
rect 77 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 30
rect 39 16 41 30
rect 49 16 51 30
rect 59 16 61 30
rect 69 21 71 30
rect 81 21 83 30
<< pmos >>
rect 12 42 14 70
rect 19 42 21 70
rect 29 42 31 70
rect 36 42 38 70
rect 52 42 54 70
rect 59 42 61 70
rect 69 42 71 70
rect 76 42 78 70
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 24 35 26 37
rect 37 35 39 37
rect 51 35 53 37
rect 67 35 69 37
rect 83 35 85 37
<< ndifct0 >>
rect 4 18 6 20
rect 24 18 26 20
rect 44 25 46 27
rect 44 18 46 20
rect 54 18 56 20
rect 64 26 66 28
rect 86 23 88 25
<< ndifct1 >>
rect 14 26 16 28
rect 34 26 36 28
rect 75 9 77 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 7 66 9 68
rect 7 59 9 61
rect 24 59 26 61
rect 45 66 47 68
rect 45 59 47 61
rect 83 59 85 61
rect 83 52 85 54
<< pdifct1 >>
rect 24 52 26 54
rect 64 59 66 61
rect 64 52 66 54
<< alu0 >>
rect 5 66 7 68
rect 9 66 11 68
rect 5 61 11 66
rect 43 66 45 68
rect 47 66 49 68
rect 5 59 7 61
rect 9 59 11 61
rect 5 58 11 59
rect 23 61 27 63
rect 23 59 24 61
rect 26 59 27 61
rect 23 54 27 59
rect 43 61 49 66
rect 43 59 45 61
rect 47 59 49 61
rect 43 58 49 59
rect 82 61 86 68
rect 82 59 83 61
rect 85 59 86 61
rect 82 54 86 59
rect 82 52 83 54
rect 85 52 86 54
rect 82 50 86 52
rect 10 42 12 46
rect 10 37 14 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 43 28 68 29
rect 43 27 64 28
rect 43 25 44 27
rect 46 26 64 27
rect 66 26 68 28
rect 46 25 68 26
rect 85 25 89 27
rect 43 21 48 25
rect 64 21 68 25
rect 85 23 86 25
rect 88 23 89 25
rect 85 21 89 23
rect 2 20 48 21
rect 2 18 4 20
rect 6 18 24 20
rect 26 18 44 20
rect 46 18 48 20
rect 2 17 48 18
rect 52 20 58 21
rect 52 18 54 20
rect 56 18 58 20
rect 52 12 58 18
rect 64 17 89 21
<< labels >>
rlabel alu0 45 23 45 23 6 n3
rlabel ndifct0 25 19 25 19 6 n3
rlabel alu0 55 27 55 27 6 n3
rlabel alu0 87 22 87 22 6 n3
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 36 20 36 6 b2
rlabel alu1 20 44 20 44 6 b1
rlabel alu1 28 36 28 36 6 b2
rlabel alu1 28 44 28 44 6 b1
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 36 44 36 44 6 b1
rlabel alu1 44 36 44 36 6 b1
rlabel polyct1 52 36 52 36 6 a1
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 76 28 76 28 6 a2
rlabel alu1 60 44 60 44 6 a1
rlabel polyct1 68 36 68 36 6 a2
rlabel alu1 68 44 68 44 6 a1
rlabel alu1 76 48 76 48 6 a1
rlabel alu1 60 52 60 52 6 z
rlabel alu1 68 60 68 60 6 z
rlabel polyct1 84 36 84 36 6 a1
<< end >>
