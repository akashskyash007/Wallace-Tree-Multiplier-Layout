magic
tech scmos
timestamp 1199202612
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 62 31 67
rect 39 62 41 67
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 19 33 31 35
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 37 42 39
rect 36 35 38 37
rect 40 35 42 37
rect 36 33 42 35
rect 36 30 38 33
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
<< ndif >>
rect 3 11 12 30
rect 3 9 6 11
rect 8 10 12 11
rect 14 10 19 30
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 10 29 19
rect 31 10 36 30
rect 38 21 46 30
rect 38 19 42 21
rect 44 19 46 21
rect 38 17 46 19
rect 38 10 43 17
rect 8 9 10 10
rect 3 7 10 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 62 27 70
rect 21 60 29 62
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 60 39 62
rect 31 58 34 60
rect 36 58 39 60
rect 31 53 39 58
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 60 49 62
rect 41 58 44 60
rect 46 58 49 60
rect 41 53 49 58
rect 41 51 44 53
rect 46 51 49 53
rect 41 42 49 51
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 33 60 38 63
rect 33 58 34 60
rect 36 58 38 60
rect 33 54 38 58
rect 12 53 38 54
rect 12 51 14 53
rect 16 51 34 53
rect 36 51 38 53
rect 12 50 38 51
rect 12 47 18 50
rect 2 46 18 47
rect 2 44 14 46
rect 16 44 18 46
rect 2 43 18 44
rect 2 22 6 43
rect 25 42 39 46
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 10 26 47 30
rect 2 21 31 22
rect 2 19 24 21
rect 26 19 31 21
rect 2 18 31 19
rect -2 11 58 12
rect -2 9 6 11
rect 8 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 62
rect 39 42 41 62
<< polyct0 >>
rect 38 35 40 37
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
<< ndifct0 >>
rect 42 19 44 21
<< ndifct1 >>
rect 6 9 8 11
rect 24 19 26 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 58 26 60
rect 44 58 46 60
rect 44 51 46 53
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
rect 34 58 36 60
rect 34 51 36 53
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 60 28 68
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 42 60 48 68
rect 42 58 44 60
rect 46 58 48 60
rect 42 53 48 58
rect 42 51 44 53
rect 46 51 48 53
rect 42 50 48 51
rect 36 37 42 38
rect 36 35 38 37
rect 40 35 42 37
rect 36 30 42 35
rect 40 21 46 22
rect 40 19 42 21
rect 44 19 46 21
rect 40 12 46 19
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a
<< end >>
