magic
tech scmos
timestamp 1199203479
<< ab >>
rect 0 0 104 80
<< nwell >>
rect -5 36 109 88
<< pwell >>
rect -5 -8 109 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 53 70 55 74
rect 63 68 65 73
rect 73 68 75 73
rect 83 61 85 66
rect 93 61 95 65
rect 9 23 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 37 28 39
rect 16 35 24 37
rect 26 35 28 37
rect 16 33 28 35
rect 23 30 25 33
rect 33 30 35 42
rect 43 39 45 50
rect 53 47 55 50
rect 63 47 65 50
rect 73 47 75 50
rect 53 45 65 47
rect 43 37 57 39
rect 43 35 51 37
rect 53 35 57 37
rect 43 33 57 35
rect 63 35 65 45
rect 69 45 75 47
rect 69 43 71 45
rect 73 43 75 45
rect 69 41 75 43
rect 83 35 85 42
rect 93 39 95 42
rect 93 37 102 39
rect 93 35 98 37
rect 100 35 102 37
rect 63 33 102 35
rect 43 30 45 33
rect 55 30 57 33
rect 78 30 80 33
rect 5 21 11 23
rect 5 19 7 21
rect 9 19 11 21
rect 5 17 11 19
rect 55 19 57 24
rect 63 20 69 22
rect 43 12 45 17
rect 23 6 25 11
rect 33 8 35 11
rect 63 18 65 20
rect 67 18 69 20
rect 63 16 69 18
rect 63 8 65 16
rect 33 6 65 8
rect 78 6 80 11
<< ndif >>
rect 18 23 23 30
rect 16 21 23 23
rect 16 19 18 21
rect 20 19 23 21
rect 16 17 23 19
rect 18 11 23 17
rect 25 28 33 30
rect 25 26 28 28
rect 30 26 33 28
rect 25 11 33 26
rect 35 28 43 30
rect 35 26 38 28
rect 40 26 43 28
rect 35 17 43 26
rect 45 24 55 30
rect 57 28 64 30
rect 57 26 60 28
rect 62 26 64 28
rect 57 24 64 26
rect 71 28 78 30
rect 71 26 73 28
rect 75 26 78 28
rect 45 17 53 24
rect 35 11 40 17
rect 47 14 53 17
rect 47 12 49 14
rect 51 12 53 14
rect 47 10 53 12
rect 71 21 78 26
rect 71 19 73 21
rect 75 19 78 21
rect 71 17 78 19
rect 73 11 78 17
rect 80 22 88 30
rect 80 20 83 22
rect 85 20 88 22
rect 80 15 88 20
rect 80 13 83 15
rect 85 13 88 15
rect 80 11 88 13
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 42 16 70
rect 18 61 26 70
rect 18 59 21 61
rect 23 59 26 61
rect 18 46 26 59
rect 18 44 21 46
rect 23 44 26 46
rect 18 42 26 44
rect 28 42 33 70
rect 35 68 43 70
rect 35 66 38 68
rect 40 66 43 68
rect 35 50 43 66
rect 45 54 53 70
rect 45 52 48 54
rect 50 52 53 54
rect 45 50 53 52
rect 55 68 60 70
rect 55 61 63 68
rect 55 59 58 61
rect 60 59 63 61
rect 55 50 63 59
rect 65 61 73 68
rect 65 59 68 61
rect 70 59 73 61
rect 65 54 73 59
rect 65 52 68 54
rect 70 52 73 54
rect 65 50 73 52
rect 75 61 81 68
rect 75 59 83 61
rect 75 57 78 59
rect 80 57 83 59
rect 75 50 83 57
rect 35 42 41 50
rect 77 42 83 50
rect 85 53 93 61
rect 85 51 88 53
rect 90 51 93 53
rect 85 46 93 51
rect 85 44 88 46
rect 90 44 93 46
rect 85 42 93 44
rect 95 59 102 61
rect 95 57 98 59
rect 100 57 102 59
rect 95 52 102 57
rect 95 50 98 52
rect 100 50 102 52
rect 95 42 102 50
<< alu1 >>
rect -2 81 106 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 106 81
rect -2 68 106 79
rect 18 61 63 62
rect 18 59 21 61
rect 23 59 58 61
rect 60 59 63 61
rect 18 58 63 59
rect 18 48 22 58
rect 18 47 24 48
rect 10 46 24 47
rect 10 44 21 46
rect 23 44 24 46
rect 10 42 24 44
rect 10 30 14 42
rect 49 45 75 46
rect 49 43 71 45
rect 73 43 75 45
rect 49 42 75 43
rect 49 37 55 42
rect 49 35 51 37
rect 53 35 55 37
rect 49 34 55 35
rect 97 37 102 39
rect 97 35 98 37
rect 100 35 102 37
rect 10 28 32 30
rect 10 26 28 28
rect 30 26 32 28
rect 26 25 32 26
rect 97 23 102 35
rect 90 17 102 23
rect -2 1 106 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 106 1
rect -2 -2 106 -1
<< ptie >>
rect 0 1 104 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 104 1
rect 0 -3 104 -1
<< ntie >>
rect 0 81 104 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 104 81
rect 0 77 104 79
<< nmos >>
rect 23 11 25 30
rect 33 11 35 30
rect 43 17 45 30
rect 55 24 57 30
rect 78 11 80 30
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 50 45 70
rect 53 50 55 70
rect 63 50 65 68
rect 73 50 75 68
rect 83 42 85 61
rect 93 42 95 61
<< polyct0 >>
rect 24 35 26 37
rect 7 19 9 21
rect 65 18 67 20
<< polyct1 >>
rect 51 35 53 37
rect 71 43 73 45
rect 98 35 100 37
<< ndifct0 >>
rect 18 19 20 21
rect 38 26 40 28
rect 60 26 62 28
rect 73 26 75 28
rect 49 12 51 14
rect 73 19 75 21
rect 83 20 85 22
rect 83 13 85 15
<< ndifct1 >>
rect 28 26 30 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 38 66 40 68
rect 48 52 50 54
rect 68 59 70 61
rect 68 52 70 54
rect 78 57 80 59
rect 88 51 90 53
rect 88 44 90 46
rect 98 57 100 59
rect 98 50 100 52
<< pdifct1 >>
rect 21 59 23 61
rect 21 44 23 46
rect 58 59 60 61
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 36 66 38 68
rect 40 66 42 68
rect 36 65 42 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 67 61 71 63
rect 67 59 68 61
rect 70 59 71 61
rect 46 54 52 55
rect 67 54 71 59
rect 77 59 81 68
rect 77 57 78 59
rect 80 57 81 59
rect 77 55 81 57
rect 97 59 101 68
rect 97 57 98 59
rect 100 57 101 59
rect 36 52 48 54
rect 50 52 68 54
rect 70 52 71 54
rect 36 50 71 52
rect 87 53 91 55
rect 87 51 88 53
rect 90 51 91 53
rect 36 38 40 50
rect 87 46 91 51
rect 97 52 101 57
rect 97 50 98 52
rect 100 50 101 52
rect 97 48 101 50
rect 22 37 40 38
rect 22 35 24 37
rect 26 35 40 37
rect 22 34 40 35
rect 87 44 88 46
rect 90 44 91 46
rect 87 38 91 44
rect 72 34 91 38
rect 36 30 40 34
rect 36 28 64 30
rect 36 26 38 28
rect 40 26 60 28
rect 62 26 64 28
rect 36 25 42 26
rect 58 25 64 26
rect 72 28 76 34
rect 72 26 73 28
rect 75 26 76 28
rect 72 22 76 26
rect 5 21 76 22
rect 5 19 7 21
rect 9 19 18 21
rect 20 20 73 21
rect 20 19 65 20
rect 5 18 65 19
rect 67 19 73 20
rect 75 19 76 21
rect 67 18 76 19
rect 63 17 76 18
rect 82 22 86 24
rect 82 20 83 22
rect 85 20 86 22
rect 82 15 86 20
rect 47 14 53 15
rect 47 12 49 14
rect 51 12 53 14
rect 82 13 83 15
rect 85 13 86 15
rect 82 12 86 13
<< labels >>
rlabel alu0 31 36 31 36 6 an
rlabel ndifct0 74 27 74 27 6 bn
rlabel alu0 40 20 40 20 6 bn
rlabel alu0 50 28 50 28 6 an
rlabel alu0 53 52 53 52 6 an
rlabel alu0 69 56 69 56 6 an
rlabel alu0 89 44 89 44 6 bn
rlabel alu1 20 28 20 28 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 28 28 28 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 52 6 52 6 6 vss
rlabel alu1 68 44 68 44 6 a
rlabel alu1 60 44 60 44 6 a
rlabel alu1 52 40 52 40 6 a
rlabel alu1 60 60 60 60 6 z
rlabel alu1 52 60 52 60 6 z
rlabel alu1 52 74 52 74 6 vdd
rlabel alu1 92 20 92 20 6 b
rlabel alu1 100 28 100 28 6 b
<< end >>
