magic
tech scmos
timestamp 1199468973
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 11 93 13 98
rect 23 83 25 88
rect 35 83 37 88
rect 47 83 49 88
rect 59 83 61 87
rect 11 47 13 55
rect 23 54 25 59
rect 35 54 37 59
rect 47 54 49 59
rect 23 52 31 54
rect 23 51 27 52
rect 25 50 27 51
rect 29 50 31 52
rect 25 48 31 50
rect 35 52 43 54
rect 35 50 39 52
rect 41 50 43 52
rect 35 48 43 50
rect 47 52 53 54
rect 59 53 61 59
rect 47 50 49 52
rect 51 50 53 52
rect 47 48 53 50
rect 57 51 63 53
rect 57 49 59 51
rect 61 49 63 51
rect 11 45 21 47
rect 15 43 17 45
rect 19 43 21 45
rect 15 41 21 43
rect 15 38 17 41
rect 29 38 31 48
rect 37 38 39 48
rect 47 44 49 48
rect 45 41 49 44
rect 57 47 63 49
rect 57 43 59 47
rect 53 41 59 43
rect 45 38 47 41
rect 53 38 55 41
rect 15 14 17 19
rect 29 5 31 10
rect 37 5 39 10
rect 45 5 47 10
rect 53 5 55 10
<< ndif >>
rect 7 36 15 38
rect 7 34 9 36
rect 11 34 15 36
rect 7 28 15 34
rect 7 26 9 28
rect 11 26 15 28
rect 7 24 15 26
rect 10 19 15 24
rect 17 22 29 38
rect 17 20 22 22
rect 24 20 29 22
rect 17 19 29 20
rect 19 14 29 19
rect 19 12 22 14
rect 24 12 29 14
rect 19 10 29 12
rect 31 10 37 38
rect 39 10 45 38
rect 47 10 53 38
rect 55 33 60 38
rect 55 31 63 33
rect 55 29 59 31
rect 61 29 63 31
rect 55 23 63 29
rect 55 21 59 23
rect 61 21 63 23
rect 55 19 63 21
rect 55 10 60 19
<< pdif >>
rect 61 93 67 95
rect 6 69 11 93
rect 3 67 11 69
rect 3 65 5 67
rect 7 65 11 67
rect 3 59 11 65
rect 3 57 5 59
rect 7 57 11 59
rect 3 55 11 57
rect 13 91 21 93
rect 39 91 45 93
rect 13 89 17 91
rect 19 89 21 91
rect 13 83 21 89
rect 39 89 41 91
rect 43 89 45 91
rect 61 91 63 93
rect 65 91 67 93
rect 61 89 67 91
rect 39 83 45 89
rect 63 83 67 89
rect 13 59 23 83
rect 25 81 35 83
rect 25 79 29 81
rect 31 79 35 81
rect 25 59 35 79
rect 37 59 47 83
rect 49 81 59 83
rect 49 79 53 81
rect 55 79 59 81
rect 49 59 59 79
rect 61 59 67 83
rect 13 55 21 59
<< alu1 >>
rect -2 95 72 100
rect -2 93 29 95
rect 31 93 72 95
rect -2 91 63 93
rect 65 91 72 93
rect -2 89 17 91
rect 19 89 41 91
rect 43 89 72 91
rect -2 88 72 89
rect 18 81 57 82
rect 18 79 29 81
rect 31 79 53 81
rect 55 79 57 81
rect 18 78 57 79
rect 8 68 12 73
rect 3 67 12 68
rect 3 65 5 67
rect 7 65 12 67
rect 3 64 12 65
rect 8 60 12 64
rect 3 59 12 60
rect 3 57 5 59
rect 7 57 12 59
rect 3 56 12 57
rect 8 36 12 56
rect 18 47 22 78
rect 28 68 43 73
rect 47 68 62 73
rect 28 54 32 68
rect 37 58 52 63
rect 26 52 32 54
rect 26 50 27 52
rect 29 50 32 52
rect 26 47 32 50
rect 38 52 42 54
rect 38 50 39 52
rect 41 50 42 52
rect 16 45 22 47
rect 16 43 17 45
rect 19 43 22 45
rect 16 42 22 43
rect 16 41 33 42
rect 18 38 33 41
rect 8 34 9 36
rect 11 34 12 36
rect 8 32 12 34
rect 8 28 23 32
rect 8 26 9 28
rect 11 26 12 28
rect 8 17 12 26
rect 21 22 25 24
rect 21 20 22 22
rect 24 20 25 22
rect 21 14 25 20
rect 29 22 33 38
rect 38 32 42 50
rect 48 52 52 58
rect 48 50 49 52
rect 51 50 52 52
rect 48 37 52 50
rect 58 51 62 68
rect 58 49 59 51
rect 61 49 62 51
rect 58 47 62 49
rect 38 27 53 32
rect 58 31 62 33
rect 58 29 59 31
rect 61 29 62 31
rect 58 23 62 29
rect 58 22 59 23
rect 29 21 59 22
rect 61 21 62 23
rect 29 18 62 21
rect 21 12 22 14
rect 24 12 25 14
rect -2 7 72 12
rect -2 5 9 7
rect 11 5 72 7
rect -2 0 72 5
<< ptie >>
rect 7 7 13 9
rect 7 5 9 7
rect 11 5 13 7
rect 7 3 13 5
<< ntie >>
rect 27 95 33 97
rect 27 93 29 95
rect 31 93 33 95
rect 27 91 33 93
<< nmos >>
rect 15 19 17 38
rect 29 10 31 38
rect 37 10 39 38
rect 45 10 47 38
rect 53 10 55 38
<< pmos >>
rect 11 55 13 93
rect 23 59 25 83
rect 35 59 37 83
rect 47 59 49 83
rect 59 59 61 83
<< polyct1 >>
rect 27 50 29 52
rect 39 50 41 52
rect 49 50 51 52
rect 59 49 61 51
rect 17 43 19 45
<< ndifct1 >>
rect 9 34 11 36
rect 9 26 11 28
rect 22 20 24 22
rect 22 12 24 14
rect 59 29 61 31
rect 59 21 61 23
<< ntiect1 >>
rect 29 93 31 95
<< ptiect1 >>
rect 9 5 11 7
<< pdifct1 >>
rect 5 65 7 67
rect 5 57 7 59
rect 17 89 19 91
rect 41 89 43 91
rect 63 91 65 93
rect 29 79 31 81
rect 53 79 55 81
<< labels >>
rlabel polyct1 18 44 18 44 6 zn
rlabel pdifct1 30 80 30 80 6 zn
rlabel ndifct1 60 22 60 22 6 zn
rlabel ndifct1 60 30 60 30 6 zn
rlabel pdifct1 54 80 54 80 6 zn
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 30 20 30 6 z
rlabel alu1 30 60 30 60 6 a
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 40 40 40 6 b
rlabel alu1 50 30 50 30 6 b
rlabel alu1 50 50 50 50 6 c
rlabel alu1 50 70 50 70 6 d
rlabel alu1 40 70 40 70 6 a
rlabel alu1 40 60 40 60 6 c
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 60 60 60 6 d
<< end >>
