magic
tech scmos
timestamp 1199202727
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 30 70 32 74
rect 40 70 42 74
rect 9 39 11 42
rect 19 39 21 42
rect 30 39 32 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 32 39
rect 19 35 27 37
rect 29 35 32 37
rect 40 39 42 42
rect 40 37 47 39
rect 40 35 43 37
rect 45 35 47 37
rect 19 33 32 35
rect 13 29 15 33
rect 20 29 22 33
rect 30 29 32 33
rect 37 33 47 35
rect 37 29 39 33
rect 13 6 15 11
rect 20 6 22 11
rect 30 6 32 11
rect 37 6 39 11
<< ndif >>
rect 4 14 13 29
rect 4 12 7 14
rect 9 12 13 14
rect 4 11 13 12
rect 15 11 20 29
rect 22 21 30 29
rect 22 19 25 21
rect 27 19 30 21
rect 22 11 30 19
rect 32 11 37 29
rect 39 22 47 29
rect 39 20 42 22
rect 44 20 47 22
rect 39 15 47 20
rect 39 13 42 15
rect 44 13 47 15
rect 39 11 47 13
rect 4 9 11 11
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 60 9 66
rect 2 58 4 60
rect 6 58 9 60
rect 2 42 9 58
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 30 70
rect 21 66 24 68
rect 26 66 30 68
rect 21 61 30 66
rect 21 59 24 61
rect 26 59 30 61
rect 21 42 30 59
rect 32 60 40 70
rect 32 58 35 60
rect 37 58 40 60
rect 32 53 40 58
rect 32 51 35 53
rect 37 51 40 53
rect 32 42 40 51
rect 42 68 50 70
rect 42 66 45 68
rect 47 66 50 68
rect 42 61 50 66
rect 42 59 45 61
rect 47 59 50 61
rect 42 42 50 59
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 34 60 39 63
rect 34 58 35 60
rect 37 58 39 60
rect 34 54 39 58
rect 12 53 39 54
rect 12 51 14 53
rect 16 51 35 53
rect 37 51 39 53
rect 12 50 39 51
rect 12 47 18 50
rect 2 46 18 47
rect 2 44 14 46
rect 16 44 18 46
rect 2 43 18 44
rect 2 22 6 43
rect 25 42 39 46
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 30 47 35
rect 10 26 47 30
rect 2 21 31 22
rect 2 19 25 21
rect 27 19 31 21
rect 2 18 31 19
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 13 11 15 29
rect 20 11 22 29
rect 30 11 32 29
rect 37 11 39 29
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 30 42 32 70
rect 40 42 42 70
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 43 35 45 37
<< ndifct0 >>
rect 7 12 9 14
rect 42 20 44 22
rect 42 13 44 15
<< ndifct1 >>
rect 25 19 27 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 58 6 60
rect 24 66 26 68
rect 24 59 26 61
rect 45 66 47 68
rect 45 59 47 61
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
rect 35 58 37 60
rect 35 51 37 53
<< alu0 >>
rect 3 66 4 68
rect 6 66 7 68
rect 3 60 7 66
rect 3 58 4 60
rect 6 58 7 60
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 43 66 45 68
rect 47 66 49 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 43 61 49 66
rect 43 59 45 61
rect 47 59 49 61
rect 43 58 49 59
rect 3 56 7 58
rect 40 22 46 23
rect 40 20 42 22
rect 44 20 46 22
rect 40 15 46 20
rect 5 14 11 15
rect 5 12 7 14
rect 9 12 11 14
rect 40 13 42 15
rect 44 13 46 15
rect 40 12 46 13
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 a
<< end >>
