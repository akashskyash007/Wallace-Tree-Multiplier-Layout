magic
tech scmos
timestamp 1199542547
<< ab >>
rect 0 0 120 100
<< nwell >>
rect -2 48 122 104
<< pwell >>
rect -2 -4 122 48
<< poly >>
rect 93 95 95 98
rect 105 95 107 98
rect 11 85 13 88
rect 23 85 25 88
rect 31 85 33 88
rect 47 85 49 88
rect 55 85 57 88
rect 67 85 69 88
rect 11 41 13 65
rect 23 63 25 65
rect 17 61 25 63
rect 17 59 19 61
rect 21 59 23 61
rect 17 57 23 59
rect 31 43 33 65
rect 47 57 49 65
rect 55 63 57 65
rect 55 61 63 63
rect 57 59 59 61
rect 61 59 63 61
rect 57 57 63 59
rect 47 55 53 57
rect 47 53 49 55
rect 51 53 53 55
rect 47 51 53 53
rect 37 49 43 51
rect 37 47 39 49
rect 41 47 43 49
rect 67 47 69 65
rect 73 51 79 53
rect 93 51 95 55
rect 105 51 107 55
rect 73 49 75 51
rect 77 49 107 51
rect 73 47 79 49
rect 37 45 69 47
rect 27 41 33 43
rect 11 39 29 41
rect 31 39 49 41
rect 11 15 13 39
rect 27 37 33 39
rect 17 31 23 33
rect 17 29 19 31
rect 21 29 23 31
rect 17 27 25 29
rect 23 15 25 27
rect 29 21 35 23
rect 29 19 31 21
rect 33 19 35 21
rect 29 17 35 19
rect 31 15 33 17
rect 47 15 49 39
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 55 27 63 29
rect 55 15 57 27
rect 67 15 69 45
rect 93 25 95 49
rect 105 25 107 49
rect 11 2 13 5
rect 23 2 25 5
rect 31 2 33 5
rect 47 2 49 5
rect 55 2 57 5
rect 67 2 69 5
rect 93 2 95 5
rect 105 2 107 5
<< ndif >>
rect 3 21 9 23
rect 3 19 5 21
rect 7 19 9 21
rect 3 15 9 19
rect 37 31 45 33
rect 37 29 39 31
rect 41 29 45 31
rect 37 15 45 29
rect 71 21 77 23
rect 71 19 73 21
rect 75 19 77 21
rect 71 15 77 19
rect 3 5 11 15
rect 13 11 23 15
rect 13 9 17 11
rect 19 9 23 11
rect 13 5 23 9
rect 25 5 31 15
rect 33 5 47 15
rect 49 5 55 15
rect 57 11 67 15
rect 57 9 61 11
rect 63 9 67 11
rect 57 5 67 9
rect 69 5 77 15
rect 85 21 93 25
rect 85 19 87 21
rect 89 19 93 21
rect 85 11 93 19
rect 85 9 87 11
rect 89 9 93 11
rect 85 5 93 9
rect 95 21 105 25
rect 95 19 99 21
rect 101 19 105 21
rect 95 5 105 19
rect 107 21 115 25
rect 107 19 111 21
rect 113 19 115 21
rect 107 11 115 19
rect 107 9 111 11
rect 113 9 115 11
rect 107 5 115 9
<< pdif >>
rect 15 91 21 93
rect 59 91 65 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 59 89 61 91
rect 63 89 65 91
rect 59 85 65 89
rect 85 91 93 95
rect 85 89 87 91
rect 89 89 93 91
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 65 23 85
rect 25 65 31 85
rect 33 81 47 85
rect 33 79 39 81
rect 41 79 47 81
rect 33 71 47 79
rect 33 69 39 71
rect 41 69 47 71
rect 33 65 47 69
rect 49 65 55 85
rect 57 65 67 85
rect 69 81 77 85
rect 69 79 73 81
rect 75 79 77 81
rect 69 69 77 79
rect 69 67 73 69
rect 75 67 77 69
rect 69 65 77 67
rect 85 81 93 89
rect 85 79 87 81
rect 89 79 93 81
rect 85 71 93 79
rect 85 69 87 71
rect 89 69 93 71
rect 85 61 93 69
rect 85 59 87 61
rect 89 59 93 61
rect 85 55 93 59
rect 95 81 105 95
rect 95 79 99 81
rect 101 79 105 81
rect 95 71 105 79
rect 95 69 99 71
rect 101 69 105 71
rect 95 61 105 69
rect 95 59 99 61
rect 101 59 105 61
rect 95 55 105 59
rect 107 91 115 95
rect 107 89 111 91
rect 113 89 115 91
rect 107 81 115 89
rect 107 79 111 81
rect 113 79 115 81
rect 107 71 115 79
rect 107 69 111 71
rect 113 69 115 71
rect 107 61 115 69
rect 107 59 111 61
rect 113 59 115 61
rect 107 55 115 59
<< alu1 >>
rect -2 95 122 100
rect -2 93 29 95
rect 31 93 39 95
rect 41 93 49 95
rect 51 93 122 95
rect -2 91 122 93
rect -2 89 17 91
rect 19 89 61 91
rect 63 89 87 91
rect 89 89 111 91
rect 113 89 122 91
rect -2 88 122 89
rect 4 81 8 82
rect 4 79 5 81
rect 7 79 8 81
rect 4 78 8 79
rect 5 72 7 78
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 22 7 68
rect 18 61 22 82
rect 18 59 19 61
rect 21 59 22 61
rect 18 31 22 59
rect 18 29 19 31
rect 21 29 22 31
rect 18 28 22 29
rect 28 41 32 82
rect 38 81 42 82
rect 38 79 39 81
rect 41 79 42 81
rect 38 78 42 79
rect 39 72 41 78
rect 38 71 42 72
rect 38 69 39 71
rect 41 69 42 71
rect 38 68 42 69
rect 39 50 41 68
rect 58 61 62 82
rect 72 81 76 82
rect 72 79 73 81
rect 75 79 76 81
rect 72 78 76 79
rect 86 81 90 88
rect 86 79 87 81
rect 89 79 90 81
rect 73 70 75 78
rect 86 71 90 79
rect 72 69 76 70
rect 72 67 73 69
rect 75 67 76 69
rect 72 66 76 67
rect 86 69 87 71
rect 89 69 90 71
rect 58 59 59 61
rect 61 59 62 61
rect 48 55 52 56
rect 48 53 49 55
rect 51 53 52 55
rect 48 52 52 53
rect 38 49 42 50
rect 38 47 39 49
rect 41 47 42 49
rect 38 46 42 47
rect 28 39 29 41
rect 31 39 32 41
rect 28 28 32 39
rect 39 32 41 46
rect 38 31 42 32
rect 38 29 39 31
rect 41 29 42 31
rect 38 28 42 29
rect 4 21 8 22
rect 30 21 34 22
rect 49 21 51 52
rect 4 19 5 21
rect 7 19 31 21
rect 33 19 51 21
rect 58 31 62 59
rect 58 29 59 31
rect 61 29 62 31
rect 4 18 8 19
rect 30 18 34 19
rect 58 18 62 29
rect 73 52 75 66
rect 86 61 90 69
rect 86 59 87 61
rect 89 59 90 61
rect 86 58 90 59
rect 98 81 102 82
rect 98 79 99 81
rect 101 79 102 81
rect 98 71 102 79
rect 98 69 99 71
rect 101 69 102 71
rect 98 61 102 69
rect 98 59 99 61
rect 101 59 102 61
rect 73 51 78 52
rect 73 49 75 51
rect 77 49 78 51
rect 73 48 78 49
rect 73 22 75 48
rect 72 21 76 22
rect 72 19 73 21
rect 75 19 76 21
rect 72 18 76 19
rect 86 21 90 22
rect 86 19 87 21
rect 89 19 90 21
rect 86 12 90 19
rect 98 21 102 59
rect 110 81 114 88
rect 110 79 111 81
rect 113 79 114 81
rect 110 71 114 79
rect 110 69 111 71
rect 113 69 114 71
rect 110 61 114 69
rect 110 59 111 61
rect 113 59 114 61
rect 110 58 114 59
rect 98 19 99 21
rect 101 19 102 21
rect 98 18 102 19
rect 110 21 114 22
rect 110 19 111 21
rect 113 19 114 21
rect 110 12 114 19
rect -2 11 122 12
rect -2 9 17 11
rect 19 9 61 11
rect 63 9 87 11
rect 89 9 111 11
rect 113 9 122 11
rect -2 0 122 9
<< ntie >>
rect 27 95 53 97
rect 27 93 29 95
rect 31 93 39 95
rect 41 93 49 95
rect 51 93 53 95
rect 27 91 53 93
<< nmos >>
rect 11 5 13 15
rect 23 5 25 15
rect 31 5 33 15
rect 47 5 49 15
rect 55 5 57 15
rect 67 5 69 15
rect 93 5 95 25
rect 105 5 107 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 31 65 33 85
rect 47 65 49 85
rect 55 65 57 85
rect 67 65 69 85
rect 93 55 95 95
rect 105 55 107 95
<< polyct1 >>
rect 19 59 21 61
rect 59 59 61 61
rect 49 53 51 55
rect 39 47 41 49
rect 75 49 77 51
rect 29 39 31 41
rect 19 29 21 31
rect 31 19 33 21
rect 59 29 61 31
<< ndifct1 >>
rect 5 19 7 21
rect 39 29 41 31
rect 73 19 75 21
rect 17 9 19 11
rect 61 9 63 11
rect 87 19 89 21
rect 87 9 89 11
rect 99 19 101 21
rect 111 19 113 21
rect 111 9 113 11
<< ntiect1 >>
rect 29 93 31 95
rect 39 93 41 95
rect 49 93 51 95
<< pdifct1 >>
rect 17 89 19 91
rect 61 89 63 91
rect 87 89 89 91
rect 5 79 7 81
rect 5 69 7 71
rect 39 79 41 81
rect 39 69 41 71
rect 73 79 75 81
rect 73 67 75 69
rect 87 79 89 81
rect 87 69 89 71
rect 87 59 89 61
rect 99 79 101 81
rect 99 69 101 71
rect 99 59 101 61
rect 111 89 113 91
rect 111 79 113 81
rect 111 69 113 71
rect 111 59 113 61
<< labels >>
rlabel alu1 20 55 20 55 6 i0
rlabel alu1 30 55 30 55 6 cmd
rlabel alu1 60 6 60 6 6 vss
rlabel alu1 60 50 60 50 6 i1
rlabel alu1 60 94 60 94 6 vdd
rlabel alu1 100 50 100 50 6 nq
<< end >>
