magic
tech scmos
timestamp 1199202376
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 62 11 66
rect 9 41 11 44
rect 9 39 22 41
rect 9 37 18 39
rect 20 37 22 39
rect 9 35 22 37
rect 9 30 11 35
rect 9 18 11 23
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 23 9 26
rect 11 23 20 30
rect 13 21 20 23
rect 13 19 15 21
rect 17 19 20 21
rect 13 17 20 19
<< pdif >>
rect 13 71 20 73
rect 13 69 15 71
rect 17 69 20 71
rect 13 62 20 69
rect 4 50 9 62
rect 2 48 9 50
rect 2 46 4 48
rect 6 46 9 48
rect 2 44 9 46
rect 11 44 20 62
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 71 26 79
rect -2 69 15 71
rect 17 69 26 71
rect -2 68 26 69
rect 2 57 22 63
rect 2 48 7 50
rect 2 46 4 48
rect 6 46 7 48
rect 2 31 7 46
rect 18 41 22 57
rect 16 39 22 41
rect 16 37 18 39
rect 20 37 22 39
rect 16 35 22 37
rect 2 28 22 31
rect 2 26 4 28
rect 6 26 22 28
rect 2 25 22 26
rect -2 1 26 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 23 11 30
<< pmos >>
rect 9 44 11 62
<< polyct1 >>
rect 18 37 20 39
<< ndifct0 >>
rect 15 19 17 21
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct1 >>
rect 15 69 17 71
rect 4 46 6 48
<< alu0 >>
rect 13 21 19 22
rect 13 19 15 21
rect 17 19 19 21
rect 13 12 19 19
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 4 60 4 60 6 a
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 60 12 60 6 a
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 28 20 28 6 z
rlabel alu1 20 52 20 52 6 a
<< end >>
