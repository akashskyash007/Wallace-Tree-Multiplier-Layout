magic
tech scmos
timestamp 1199202132
<< ab >>
rect 0 0 128 72
<< nwell >>
rect -5 32 133 77
<< pwell >>
rect -5 -5 133 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 51 66 53 70
rect 58 66 60 70
rect 68 66 70 70
rect 75 66 77 70
rect 87 66 89 70
rect 97 66 99 70
rect 107 66 109 70
rect 117 54 119 59
rect 9 35 11 38
rect 2 33 11 35
rect 2 31 4 33
rect 6 31 11 33
rect 2 29 11 31
rect 9 26 11 29
rect 19 35 21 38
rect 29 35 31 38
rect 19 33 31 35
rect 19 31 27 33
rect 29 31 31 33
rect 19 29 31 31
rect 19 26 21 29
rect 29 26 31 29
rect 39 35 41 38
rect 51 35 53 38
rect 39 33 53 35
rect 39 31 43 33
rect 45 31 53 33
rect 39 29 53 31
rect 39 26 41 29
rect 51 26 53 29
rect 58 35 60 38
rect 68 35 70 38
rect 58 33 70 35
rect 58 31 66 33
rect 68 31 70 33
rect 58 29 70 31
rect 58 26 60 29
rect 68 26 70 29
rect 75 35 77 38
rect 75 33 83 35
rect 75 31 79 33
rect 81 31 83 33
rect 75 29 83 31
rect 87 31 89 38
rect 97 31 99 38
rect 87 29 99 31
rect 75 26 77 29
rect 87 27 92 29
rect 94 27 99 29
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 39 7 41 12
rect 87 25 99 27
rect 87 22 89 25
rect 97 22 99 25
rect 107 35 109 38
rect 117 35 119 38
rect 107 33 119 35
rect 107 31 115 33
rect 117 31 119 33
rect 107 29 119 31
rect 107 22 109 29
rect 117 22 119 29
rect 68 11 70 15
rect 75 11 77 15
rect 51 4 53 9
rect 58 4 60 9
rect 87 3 89 8
rect 97 3 99 8
rect 107 6 109 11
rect 117 6 119 11
<< ndif >>
rect 2 23 9 26
rect 2 21 4 23
rect 6 21 9 23
rect 2 16 9 21
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 16 19 26
rect 11 14 14 16
rect 16 14 19 16
rect 11 12 19 14
rect 21 24 29 26
rect 21 22 24 24
rect 26 22 29 24
rect 21 12 29 22
rect 31 16 39 26
rect 31 14 34 16
rect 36 14 39 16
rect 31 12 39 14
rect 41 12 51 26
rect 43 9 51 12
rect 53 9 58 26
rect 60 24 68 26
rect 60 22 63 24
rect 65 22 68 24
rect 60 15 68 22
rect 70 15 75 26
rect 77 22 85 26
rect 77 15 87 22
rect 60 9 65 15
rect 43 7 49 9
rect 43 5 45 7
rect 47 5 49 7
rect 43 3 49 5
rect 79 8 87 15
rect 89 16 97 22
rect 89 14 92 16
rect 94 14 97 16
rect 89 8 97 14
rect 99 15 107 22
rect 99 13 102 15
rect 104 13 107 15
rect 99 11 107 13
rect 109 20 117 22
rect 109 18 112 20
rect 114 18 117 20
rect 109 11 117 18
rect 119 15 126 22
rect 119 13 122 15
rect 124 13 126 15
rect 119 11 126 13
rect 99 8 105 11
rect 79 7 85 8
rect 79 5 81 7
rect 83 5 85 7
rect 79 3 85 5
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 38 19 55
rect 21 42 29 66
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 38 39 55
rect 41 64 51 66
rect 41 62 45 64
rect 47 62 51 64
rect 41 38 51 62
rect 53 38 58 66
rect 60 42 68 66
rect 60 40 63 42
rect 65 40 68 42
rect 60 38 68 40
rect 70 38 75 66
rect 77 64 87 66
rect 77 62 81 64
rect 83 62 87 64
rect 77 38 87 62
rect 89 56 97 66
rect 89 54 92 56
rect 94 54 97 56
rect 89 49 97 54
rect 89 47 92 49
rect 94 47 97 49
rect 89 38 97 47
rect 99 64 107 66
rect 99 62 102 64
rect 104 62 107 64
rect 99 56 107 62
rect 99 54 102 56
rect 104 54 107 56
rect 99 38 107 54
rect 109 54 114 66
rect 109 49 117 54
rect 109 47 112 49
rect 114 47 117 49
rect 109 42 117 47
rect 109 40 112 42
rect 114 40 117 42
rect 109 38 117 40
rect 119 52 126 54
rect 119 50 122 52
rect 124 50 126 52
rect 119 44 126 50
rect 119 42 122 44
rect 124 42 126 44
rect 119 38 126 42
<< alu1 >>
rect -2 67 130 72
rect -2 65 121 67
rect 123 65 130 67
rect -2 64 130 65
rect 2 46 79 50
rect 2 33 7 46
rect 2 31 4 33
rect 6 31 7 33
rect 2 29 7 31
rect 17 40 24 42
rect 26 40 28 42
rect 17 38 28 40
rect 17 26 21 38
rect 33 34 39 42
rect 25 33 39 34
rect 25 31 27 33
rect 29 31 39 33
rect 25 30 39 31
rect 50 40 63 42
rect 65 40 67 42
rect 50 38 67 40
rect 73 42 79 46
rect 73 38 87 42
rect 50 26 54 38
rect 17 24 67 26
rect 17 22 24 24
rect 26 22 63 24
rect 65 22 67 24
rect 114 33 126 35
rect 114 31 115 33
rect 117 31 126 33
rect 114 29 126 31
rect 122 21 126 29
rect -2 7 130 8
rect -2 5 45 7
rect 47 5 71 7
rect 73 5 81 7
rect 83 5 130 7
rect -2 0 130 5
<< ptie >>
rect 69 7 75 9
rect 69 5 71 7
rect 73 5 75 7
rect 69 3 75 5
<< ntie >>
rect 119 67 125 69
rect 119 65 121 67
rect 123 65 125 67
rect 119 63 125 65
<< nmos >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 12 31 26
rect 39 12 41 26
rect 51 9 53 26
rect 58 9 60 26
rect 68 15 70 26
rect 75 15 77 26
rect 87 8 89 22
rect 97 8 99 22
rect 107 11 109 22
rect 117 11 119 22
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 51 38 53 66
rect 58 38 60 66
rect 68 38 70 66
rect 75 38 77 66
rect 87 38 89 66
rect 97 38 99 66
rect 107 38 109 66
rect 117 38 119 54
<< polyct0 >>
rect 43 31 45 33
rect 66 31 68 33
rect 79 31 81 33
rect 92 27 94 29
<< polyct1 >>
rect 4 31 6 33
rect 27 31 29 33
rect 115 31 117 33
<< ndifct0 >>
rect 4 21 6 23
rect 4 14 6 16
rect 14 14 16 16
rect 34 14 36 16
rect 92 14 94 16
rect 102 13 104 15
rect 112 18 114 20
rect 122 13 124 15
<< ndifct1 >>
rect 24 22 26 24
rect 63 22 65 24
rect 45 5 47 7
rect 81 5 83 7
<< ntiect1 >>
rect 121 65 123 67
<< ptiect1 >>
rect 71 5 73 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 55 16 57
rect 34 55 36 57
rect 45 62 47 64
rect 81 62 83 64
rect 92 54 94 56
rect 92 47 94 49
rect 102 62 104 64
rect 102 54 104 56
rect 112 47 114 49
rect 112 40 114 42
rect 122 50 124 52
rect 122 42 124 44
<< pdifct1 >>
rect 24 40 26 42
rect 63 40 65 42
<< alu0 >>
rect 3 62 4 64
rect 6 62 7 64
rect 3 57 7 62
rect 43 62 45 64
rect 47 62 49 64
rect 43 61 49 62
rect 79 62 81 64
rect 83 62 85 64
rect 79 61 85 62
rect 101 62 102 64
rect 104 62 105 64
rect 3 55 4 57
rect 6 55 7 57
rect 3 53 7 55
rect 12 57 95 58
rect 12 55 14 57
rect 16 55 34 57
rect 36 56 95 57
rect 36 55 92 56
rect 12 54 92 55
rect 94 54 95 56
rect 22 42 28 43
rect 42 33 46 46
rect 61 42 67 43
rect 42 31 43 33
rect 45 31 46 33
rect 42 29 46 31
rect 91 49 95 54
rect 101 56 105 62
rect 101 54 102 56
rect 104 54 105 56
rect 101 52 105 54
rect 121 52 125 64
rect 91 47 92 49
rect 94 47 95 49
rect 91 45 95 47
rect 111 49 115 52
rect 111 47 112 49
rect 114 47 115 49
rect 111 43 115 47
rect 106 42 115 43
rect 106 40 112 42
rect 114 40 115 42
rect 121 50 122 52
rect 124 50 125 52
rect 121 44 125 50
rect 121 42 122 44
rect 124 42 125 44
rect 121 40 125 42
rect 106 39 115 40
rect 64 33 75 34
rect 64 31 66 33
rect 68 31 75 33
rect 64 30 75 31
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 22 21 28 22
rect 61 21 67 22
rect 71 25 75 30
rect 78 33 82 38
rect 78 31 79 33
rect 81 31 82 33
rect 78 29 82 31
rect 91 29 95 31
rect 91 27 92 29
rect 94 27 95 29
rect 91 25 95 27
rect 106 25 110 39
rect 71 21 115 25
rect 3 16 7 21
rect 111 20 115 21
rect 111 18 112 20
rect 114 18 115 20
rect 3 14 4 16
rect 6 14 7 16
rect 3 8 7 14
rect 12 16 96 17
rect 12 14 14 16
rect 16 14 34 16
rect 36 14 92 16
rect 94 14 96 16
rect 12 13 96 14
rect 101 15 105 17
rect 111 16 115 18
rect 101 13 102 15
rect 104 13 105 15
rect 101 8 105 13
rect 121 15 125 17
rect 121 13 122 15
rect 124 13 125 15
rect 121 8 125 13
<< labels >>
rlabel alu0 69 32 69 32 6 bn
rlabel alu0 54 15 54 15 6 n3
rlabel alu0 113 20 113 20 6 bn
rlabel alu0 93 26 93 26 6 bn
rlabel alu0 113 45 113 45 6 bn
rlabel alu0 93 51 93 51 6 n1
rlabel alu0 53 56 53 56 6 n1
rlabel alu1 20 24 20 24 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 4 36 4 36 6 a
rlabel alu1 12 48 12 48 6 a
rlabel alu1 20 48 20 48 6 a
rlabel alu1 28 24 28 24 6 z
rlabel alu1 36 24 36 24 6 z
rlabel alu1 44 24 44 24 6 z
rlabel polyct1 28 32 28 32 6 c
rlabel alu1 36 36 36 36 6 c
rlabel alu1 28 48 28 48 6 a
rlabel alu1 36 48 36 48 6 a
rlabel alu1 44 48 44 48 6 a
rlabel alu1 64 4 64 4 6 vss
rlabel alu1 60 24 60 24 6 z
rlabel alu1 52 32 52 32 6 z
rlabel alu1 60 40 60 40 6 z
rlabel alu1 52 48 52 48 6 a
rlabel alu1 60 48 60 48 6 a
rlabel alu1 68 48 68 48 6 a
rlabel alu1 64 68 64 68 6 vdd
rlabel alu1 84 40 84 40 6 a
rlabel alu1 76 44 76 44 6 a
rlabel polyct1 116 32 116 32 6 b
rlabel alu1 124 28 124 28 6 b
<< end >>
