magic
tech scmos
timestamp 1199202967
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 50 66 52 70
rect 60 66 62 70
rect 67 66 69 70
rect 9 30 11 39
rect 16 36 18 39
rect 26 36 28 39
rect 33 36 35 39
rect 43 36 45 39
rect 16 34 29 36
rect 33 34 45 36
rect 50 35 52 39
rect 60 35 62 39
rect 23 33 29 34
rect 23 31 25 33
rect 27 31 29 33
rect 9 28 19 30
rect 13 26 15 28
rect 17 26 19 28
rect 13 24 19 26
rect 23 29 29 31
rect 36 32 42 34
rect 36 30 38 32
rect 40 30 42 32
rect 50 33 62 35
rect 67 34 69 39
rect 50 31 52 33
rect 54 31 62 33
rect 50 30 62 31
rect 13 21 15 24
rect 23 21 25 29
rect 36 28 42 30
rect 47 28 62 30
rect 66 32 72 34
rect 66 30 68 32
rect 70 30 72 32
rect 66 28 72 30
rect 37 25 39 28
rect 47 25 49 28
rect 59 25 61 28
rect 69 25 71 28
rect 13 2 15 6
rect 23 2 25 6
rect 37 2 39 6
rect 47 2 49 6
rect 59 2 61 6
rect 69 2 71 6
<< ndif >>
rect 27 21 37 25
rect 4 10 13 21
rect 4 8 8 10
rect 10 8 13 10
rect 4 6 13 8
rect 15 17 23 21
rect 15 15 18 17
rect 20 15 23 17
rect 15 6 23 15
rect 25 10 37 21
rect 25 8 30 10
rect 32 8 37 10
rect 25 6 37 8
rect 39 17 47 25
rect 39 15 42 17
rect 44 15 47 17
rect 39 6 47 15
rect 49 10 59 25
rect 49 8 53 10
rect 55 8 59 10
rect 49 6 59 8
rect 61 17 69 25
rect 61 15 64 17
rect 66 15 69 17
rect 61 6 69 15
rect 71 17 78 25
rect 71 15 74 17
rect 76 15 78 17
rect 71 10 78 15
rect 71 8 74 10
rect 76 8 78 10
rect 71 6 78 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 39 9 55
rect 11 39 16 66
rect 18 51 26 66
rect 18 49 21 51
rect 23 49 26 51
rect 18 43 26 49
rect 18 41 21 43
rect 23 41 26 43
rect 18 39 26 41
rect 28 39 33 66
rect 35 64 43 66
rect 35 62 38 64
rect 40 62 43 64
rect 35 57 43 62
rect 35 55 38 57
rect 40 55 43 57
rect 35 39 43 55
rect 45 39 50 66
rect 52 51 60 66
rect 52 49 55 51
rect 57 49 60 51
rect 52 43 60 49
rect 52 41 55 43
rect 57 41 60 43
rect 52 39 60 41
rect 62 39 67 66
rect 69 64 77 66
rect 69 62 72 64
rect 74 62 77 64
rect 69 57 77 62
rect 69 55 72 57
rect 74 55 77 57
rect 69 39 77 55
<< alu1 >>
rect -2 64 82 72
rect 18 51 24 53
rect 18 49 21 51
rect 23 50 24 51
rect 23 49 55 50
rect 57 49 63 50
rect 18 46 63 49
rect 18 43 24 46
rect 2 41 21 43
rect 23 41 24 43
rect 2 38 24 41
rect 29 38 49 42
rect 2 18 6 38
rect 29 34 33 38
rect 45 34 49 38
rect 23 33 33 34
rect 23 31 25 33
rect 27 31 33 33
rect 23 30 33 31
rect 45 33 56 34
rect 45 31 52 33
rect 54 31 56 33
rect 45 30 56 31
rect 65 32 71 34
rect 65 30 68 32
rect 70 30 71 32
rect 14 28 18 30
rect 14 26 15 28
rect 17 26 18 28
rect 65 26 71 30
rect 14 22 71 26
rect 2 17 68 18
rect 2 15 18 17
rect 20 15 42 17
rect 44 15 64 17
rect 66 15 68 17
rect 2 14 68 15
rect -2 0 82 8
<< nmos >>
rect 13 6 15 21
rect 23 6 25 21
rect 37 6 39 25
rect 47 6 49 25
rect 59 6 61 25
rect 69 6 71 25
<< pmos >>
rect 9 39 11 66
rect 16 39 18 66
rect 26 39 28 66
rect 33 39 35 66
rect 43 39 45 66
rect 50 39 52 66
rect 60 39 62 66
rect 67 39 69 66
<< polyct0 >>
rect 38 30 40 32
<< polyct1 >>
rect 25 31 27 33
rect 15 26 17 28
rect 52 31 54 33
rect 68 30 70 32
<< ndifct0 >>
rect 8 8 10 10
rect 30 8 32 10
rect 53 8 55 10
rect 74 15 76 17
rect 74 8 76 10
<< ndifct1 >>
rect 18 15 20 17
rect 42 15 44 17
rect 64 15 66 17
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 38 62 40 64
rect 38 55 40 57
rect 55 50 57 51
rect 55 41 57 43
rect 72 62 74 64
rect 72 55 74 57
<< pdifct1 >>
rect 21 49 23 51
rect 21 41 23 43
rect 55 49 57 50
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 36 62 38 64
rect 40 62 42 64
rect 36 57 42 62
rect 36 55 38 57
rect 40 55 42 57
rect 36 54 42 55
rect 70 62 72 64
rect 74 62 76 64
rect 70 57 76 62
rect 70 55 72 57
rect 74 55 76 57
rect 70 54 76 55
rect 54 51 58 53
rect 54 50 55 51
rect 57 50 58 51
rect 54 43 58 46
rect 54 41 55 43
rect 57 41 58 43
rect 54 39 58 41
rect 37 32 41 34
rect 37 30 38 32
rect 40 30 41 32
rect 37 26 41 30
rect 72 17 78 18
rect 72 15 74 17
rect 76 15 78 17
rect 6 10 12 11
rect 6 8 8 10
rect 10 8 12 10
rect 28 10 34 11
rect 28 8 30 10
rect 32 8 34 10
rect 51 10 57 11
rect 51 8 53 10
rect 55 8 57 10
rect 72 10 78 15
rect 72 8 74 10
rect 76 8 78 10
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 24 20 24 6 a
rlabel alu1 28 24 28 24 6 a
rlabel alu1 28 32 28 32 6 b
rlabel alu1 12 40 12 40 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 36 16 36 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 60 16 60 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 52 24 52 24 6 a
rlabel alu1 60 24 60 24 6 a
rlabel alu1 52 32 52 32 6 b
rlabel alu1 52 48 52 48 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 68 28 68 28 6 a
<< end >>
