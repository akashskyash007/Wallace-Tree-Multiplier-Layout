magic
tech scmos
timestamp 1199201658
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 67 31 72
rect 39 67 41 72
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 22 39
rect 9 35 16 37
rect 18 35 22 37
rect 9 33 22 35
rect 28 37 34 39
rect 28 35 30 37
rect 32 35 34 37
rect 28 33 34 35
rect 10 30 12 33
rect 20 30 22 33
rect 32 30 34 33
rect 39 37 47 39
rect 39 35 43 37
rect 45 35 47 37
rect 39 33 47 35
rect 39 30 41 33
rect 10 11 12 16
rect 20 11 22 16
rect 32 6 34 10
rect 39 6 41 10
<< ndif >>
rect 2 16 10 30
rect 12 21 20 30
rect 12 19 15 21
rect 17 19 20 21
rect 12 16 20 19
rect 22 16 32 30
rect 2 11 8 16
rect 24 14 32 16
rect 24 12 26 14
rect 28 12 32 14
rect 2 9 4 11
rect 6 9 8 11
rect 24 10 32 12
rect 34 10 39 30
rect 41 23 46 30
rect 41 21 48 23
rect 41 19 44 21
rect 46 19 48 21
rect 41 17 48 19
rect 41 10 46 17
rect 2 7 8 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 67 27 70
rect 21 65 29 67
rect 21 63 24 65
rect 26 63 29 65
rect 21 42 29 63
rect 31 61 39 67
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 42 39 52
rect 41 65 48 67
rect 41 63 44 65
rect 46 63 48 65
rect 41 57 48 63
rect 41 55 44 57
rect 46 55 48 57
rect 41 42 48 55
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 55 17 59
rect 2 54 17 55
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 22 6 50
rect 33 42 47 46
rect 25 37 37 38
rect 25 35 30 37
rect 32 35 37 37
rect 25 34 37 35
rect 41 37 47 42
rect 41 35 43 37
rect 45 35 47 37
rect 41 34 47 35
rect 33 30 37 34
rect 33 26 47 30
rect 2 21 19 22
rect 2 19 15 21
rect 17 19 19 21
rect 2 17 19 19
rect -2 11 58 12
rect -2 9 4 11
rect 6 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 10 16 12 30
rect 20 16 22 30
rect 32 10 34 30
rect 39 10 41 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 67
rect 39 42 41 67
<< polyct0 >>
rect 16 35 18 37
<< polyct1 >>
rect 30 35 32 37
rect 43 35 45 37
<< ndifct0 >>
rect 26 12 28 14
rect 44 19 46 21
<< ndifct1 >>
rect 15 19 17 21
rect 4 9 6 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 63 26 65
rect 34 59 36 61
rect 34 52 36 54
rect 44 63 46 65
rect 44 55 46 57
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 23 65 27 68
rect 23 63 24 65
rect 26 63 27 65
rect 43 65 47 68
rect 43 63 44 65
rect 46 63 47 65
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 23 61 27 63
rect 33 61 37 63
rect 33 59 34 61
rect 36 59 37 61
rect 33 54 37 59
rect 23 52 34 54
rect 36 52 37 54
rect 43 57 47 63
rect 43 55 44 57
rect 46 55 47 57
rect 43 53 47 55
rect 23 50 37 52
rect 23 46 27 50
rect 15 42 27 46
rect 15 37 19 42
rect 15 35 16 37
rect 18 35 19 37
rect 15 30 19 35
rect 15 26 28 30
rect 24 22 28 26
rect 24 21 48 22
rect 24 19 44 21
rect 46 19 48 21
rect 24 18 48 19
rect 24 14 30 15
rect 24 12 26 14
rect 28 12 30 14
<< labels >>
rlabel polyct0 17 36 17 36 6 zn
rlabel alu0 35 56 35 56 6 zn
rlabel alu0 36 20 36 20 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 36 28 36 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 40 44 40 6 b
<< end >>
