magic
tech scmos
timestamp 1199541795
<< ab >>
rect 0 0 40 100
<< nwell >>
rect -2 48 42 104
<< pwell >>
rect -2 -4 42 48
<< poly >>
rect 23 95 25 98
rect 11 67 13 70
rect 11 53 13 55
rect 11 51 19 53
rect 11 49 15 51
rect 17 49 19 51
rect 11 47 19 49
rect 3 42 9 43
rect 23 42 25 55
rect 3 41 25 42
rect 3 39 5 41
rect 7 39 25 41
rect 3 38 25 39
rect 3 37 9 38
rect 11 31 19 33
rect 11 29 15 31
rect 17 29 19 31
rect 11 27 19 29
rect 11 25 13 27
rect 23 25 25 38
rect 11 16 13 19
rect 23 2 25 5
<< ndif >>
rect 3 23 11 25
rect 3 21 5 23
rect 7 21 11 23
rect 3 19 11 21
rect 13 19 23 25
rect 15 11 23 19
rect 15 9 17 11
rect 19 9 23 11
rect 15 5 23 9
rect 25 21 33 25
rect 25 19 29 21
rect 31 19 33 21
rect 25 5 33 19
<< pdif >>
rect 15 91 23 95
rect 15 89 17 91
rect 19 89 23 91
rect 15 67 23 89
rect 3 61 11 67
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 55 23 67
rect 25 81 33 95
rect 25 79 29 81
rect 31 79 33 81
rect 25 71 33 79
rect 25 69 29 71
rect 31 69 33 71
rect 25 61 33 69
rect 25 59 29 61
rect 31 59 33 61
rect 25 55 33 59
<< alu1 >>
rect -2 95 42 100
rect -2 93 5 95
rect 7 93 42 95
rect -2 91 42 93
rect -2 89 17 91
rect 19 89 42 91
rect -2 88 42 89
rect 4 85 8 88
rect 4 83 5 85
rect 7 83 8 85
rect 4 82 8 83
rect 4 61 8 62
rect 4 59 5 61
rect 7 59 8 61
rect 4 58 8 59
rect 5 42 7 58
rect 18 52 22 82
rect 14 51 22 52
rect 14 49 15 51
rect 17 49 22 51
rect 14 48 22 49
rect 4 41 8 42
rect 4 39 5 41
rect 7 39 8 41
rect 4 38 8 39
rect 5 24 7 38
rect 18 32 22 48
rect 14 31 22 32
rect 14 29 15 31
rect 17 29 22 31
rect 14 28 22 29
rect 4 23 8 24
rect 4 21 5 23
rect 7 21 8 23
rect 4 20 8 21
rect 18 18 22 28
rect 28 81 32 82
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 28 21 32 59
rect 28 19 29 21
rect 31 19 32 21
rect 28 18 32 19
rect -2 11 42 12
rect -2 9 17 11
rect 19 9 42 11
rect -2 0 42 9
<< ntie >>
rect 3 95 9 97
rect 3 93 5 95
rect 7 93 9 95
rect 3 85 9 93
rect 3 83 5 85
rect 7 83 9 85
rect 3 81 9 83
<< nmos >>
rect 11 19 13 25
rect 23 5 25 25
<< pmos >>
rect 11 55 13 67
rect 23 55 25 95
<< polyct1 >>
rect 15 49 17 51
rect 5 39 7 41
rect 15 29 17 31
<< ndifct1 >>
rect 5 21 7 23
rect 17 9 19 11
rect 29 19 31 21
<< ntiect1 >>
rect 5 93 7 95
rect 5 83 7 85
<< pdifct1 >>
rect 17 89 19 91
rect 5 59 7 61
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
<< labels >>
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 50 20 50 6 i
rlabel alu1 20 94 20 94 6 vdd
rlabel alu1 30 50 30 50 6 q
<< end >>
