magic
tech scmos
timestamp 1199203501
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 9 50 11 55
rect 41 68 63 70
rect 21 57 27 59
rect 21 55 23 57
rect 25 55 27 57
rect 21 53 27 55
rect 31 57 37 59
rect 31 55 33 57
rect 35 55 37 57
rect 31 53 37 55
rect 21 50 23 53
rect 31 50 33 53
rect 41 50 43 68
rect 61 59 63 68
rect 51 50 53 55
rect 9 34 11 38
rect 9 32 15 34
rect 9 30 11 32
rect 13 30 15 32
rect 21 31 23 38
rect 31 35 33 38
rect 31 33 37 35
rect 41 34 43 38
rect 51 35 53 38
rect 61 35 63 47
rect 9 28 15 30
rect 19 28 23 31
rect 35 30 37 33
rect 48 33 54 35
rect 48 31 50 33
rect 52 31 54 33
rect 9 25 11 28
rect 19 25 21 28
rect 29 25 31 29
rect 35 28 41 30
rect 48 29 54 31
rect 58 33 64 35
rect 58 31 60 33
rect 62 31 64 33
rect 58 29 64 31
rect 39 25 41 28
rect 50 26 52 29
rect 9 14 11 19
rect 19 14 21 19
rect 29 4 31 19
rect 39 14 41 19
rect 50 15 52 20
rect 61 19 63 29
rect 61 4 63 13
rect 29 2 63 4
<< ndif >>
rect 43 25 50 26
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 19 19 25
rect 21 23 29 25
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 31 23 39 25
rect 31 21 34 23
rect 36 21 39 23
rect 31 19 39 21
rect 41 24 50 25
rect 41 22 45 24
rect 47 22 50 24
rect 41 20 50 22
rect 52 20 59 26
rect 41 19 46 20
rect 13 9 17 19
rect 11 7 17 9
rect 11 5 13 7
rect 15 5 17 7
rect 11 3 17 5
rect 54 19 59 20
rect 54 13 61 19
rect 63 17 70 19
rect 63 15 66 17
rect 68 15 70 17
rect 63 13 70 15
rect 54 12 59 13
rect 53 10 59 12
rect 53 8 55 10
rect 57 8 59 10
rect 53 6 59 8
<< pdif >>
rect 13 67 19 69
rect 13 65 15 67
rect 17 65 19 67
rect 13 50 19 65
rect 53 64 59 66
rect 53 62 55 64
rect 57 62 59 64
rect 53 59 59 62
rect 53 57 61 59
rect 55 50 61 57
rect 4 44 9 50
rect 2 42 9 44
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 38 21 50
rect 23 48 31 50
rect 23 46 26 48
rect 28 46 31 48
rect 23 38 31 46
rect 33 42 41 50
rect 33 40 36 42
rect 38 40 41 42
rect 33 38 41 40
rect 43 42 51 50
rect 43 40 46 42
rect 48 40 51 42
rect 43 38 51 40
rect 53 47 61 50
rect 63 57 70 59
rect 63 55 66 57
rect 68 55 70 57
rect 63 53 70 55
rect 63 47 68 53
rect 53 38 59 47
<< alu1 >>
rect -2 67 74 72
rect -2 65 5 67
rect 7 65 15 67
rect 17 65 30 67
rect 32 65 74 67
rect -2 64 74 65
rect 9 57 27 58
rect 9 55 23 57
rect 25 55 27 57
rect 9 54 27 55
rect 18 45 22 54
rect 2 42 14 43
rect 2 40 4 42
rect 6 40 14 42
rect 2 37 14 40
rect 2 25 6 37
rect 2 23 7 25
rect 2 21 4 23
rect 6 21 7 23
rect 2 19 7 21
rect 59 33 63 35
rect 59 31 60 33
rect 62 31 63 33
rect 59 26 63 31
rect 57 22 63 26
rect 57 18 61 22
rect 49 14 61 18
rect -2 7 74 8
rect -2 5 13 7
rect 15 5 23 7
rect 25 5 74 7
rect -2 0 74 5
<< ptie >>
rect 21 7 27 9
rect 21 5 23 7
rect 25 5 27 7
rect 21 3 27 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
rect 28 67 34 69
rect 28 65 30 67
rect 32 65 34 67
rect 28 63 34 65
<< nmos >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 19 31 25
rect 39 19 41 25
rect 50 20 52 26
rect 61 13 63 19
<< pmos >>
rect 9 38 11 50
rect 21 38 23 50
rect 31 38 33 50
rect 41 38 43 50
rect 51 38 53 50
rect 61 47 63 59
<< polyct0 >>
rect 33 55 35 57
rect 11 30 13 32
rect 50 31 52 33
<< polyct1 >>
rect 23 55 25 57
rect 60 31 62 33
<< ndifct0 >>
rect 24 21 26 23
rect 34 21 36 23
rect 45 22 47 24
rect 66 15 68 17
rect 55 8 57 10
<< ndifct1 >>
rect 4 21 6 23
rect 13 5 15 7
<< ntiect1 >>
rect 5 65 7 67
rect 30 65 32 67
<< ptiect1 >>
rect 23 5 25 7
<< pdifct0 >>
rect 55 62 57 64
rect 26 46 28 48
rect 36 40 38 42
rect 46 40 48 42
rect 66 55 68 57
<< pdifct1 >>
rect 15 65 17 67
rect 4 40 6 42
<< alu0 >>
rect 53 62 55 64
rect 57 62 59 64
rect 53 61 59 62
rect 31 57 70 58
rect 31 55 33 57
rect 35 55 66 57
rect 68 55 70 57
rect 31 54 70 55
rect 25 48 56 51
rect 25 46 26 48
rect 28 47 56 48
rect 28 46 29 47
rect 9 32 16 33
rect 9 30 11 32
rect 13 30 16 32
rect 9 29 16 30
rect 12 17 16 29
rect 25 24 29 46
rect 22 23 29 24
rect 22 21 24 23
rect 26 21 29 23
rect 22 20 29 21
rect 33 42 39 44
rect 33 40 36 42
rect 38 40 39 42
rect 33 38 39 40
rect 42 42 49 44
rect 42 40 46 42
rect 48 40 49 42
rect 42 38 49 40
rect 33 23 37 38
rect 33 21 34 23
rect 36 21 37 23
rect 42 25 46 38
rect 52 35 56 47
rect 49 33 56 35
rect 49 31 50 33
rect 52 31 56 33
rect 49 29 56 31
rect 42 24 49 25
rect 42 22 45 24
rect 47 22 49 24
rect 42 21 49 22
rect 33 17 37 21
rect 66 19 70 54
rect 12 13 37 17
rect 65 17 70 19
rect 65 15 66 17
rect 68 15 70 17
rect 65 13 70 15
rect 53 10 59 11
rect 53 8 55 10
rect 57 8 59 10
<< labels >>
rlabel polyct0 12 31 12 31 6 zn
rlabel alu0 27 35 27 35 6 an
rlabel alu0 45 41 45 41 6 ai
rlabel alu0 44 32 44 32 6 ai
rlabel alu0 35 28 35 28 6 zn
rlabel alu0 54 40 54 40 6 an
rlabel alu0 50 56 50 56 6 bn
rlabel alu0 68 35 68 35 6 bn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 12 56 12 56 6 a
rlabel alu1 20 52 20 52 6 a
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 52 16 52 16 6 b
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 24 60 24 6 b
<< end >>
