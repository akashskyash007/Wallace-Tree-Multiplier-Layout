magic
tech scmos
timestamp 1199201912
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 21 39
rect 9 35 11 37
rect 13 35 21 37
rect 9 33 21 35
rect 25 37 31 39
rect 25 35 27 37
rect 29 35 31 37
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 39 37 45 39
rect 39 35 41 37
rect 43 35 45 37
rect 25 33 35 35
rect 39 33 45 35
rect 49 37 63 39
rect 49 35 51 37
rect 53 35 59 37
rect 61 35 63 37
rect 49 33 63 35
rect 67 37 73 39
rect 67 35 69 37
rect 71 35 73 37
rect 67 33 73 35
rect 77 37 88 39
rect 77 35 84 37
rect 86 35 88 37
rect 77 33 88 35
rect 9 30 11 33
rect 19 30 21 33
rect 33 30 35 33
rect 41 30 43 33
rect 49 30 51 33
rect 61 30 63 33
rect 69 30 71 33
rect 77 30 79 33
rect 9 17 11 22
rect 19 17 21 22
rect 33 7 35 12
rect 41 7 43 12
rect 49 7 51 12
rect 61 7 63 12
rect 69 7 71 12
rect 77 7 79 12
<< ndif >>
rect 2 26 9 30
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 22 19 26
rect 21 22 33 30
rect 23 12 33 22
rect 35 12 41 30
rect 43 12 49 30
rect 51 21 61 30
rect 51 19 55 21
rect 57 19 61 21
rect 51 12 61 19
rect 63 12 69 30
rect 71 12 77 30
rect 79 16 87 30
rect 79 14 82 16
rect 84 14 87 16
rect 79 12 87 14
rect 23 11 31 12
rect 23 9 26 11
rect 28 9 31 11
rect 23 7 31 9
<< pdif >>
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 42 9 58
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 61 29 70
rect 21 59 24 61
rect 26 59 29 61
rect 21 54 29 59
rect 21 52 24 54
rect 26 52 29 54
rect 21 42 29 52
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 42 39 66
rect 41 61 49 70
rect 41 59 44 61
rect 46 59 49 61
rect 41 54 49 59
rect 41 52 44 54
rect 46 52 49 54
rect 41 42 49 52
rect 51 68 59 70
rect 51 66 54 68
rect 56 66 59 68
rect 51 61 59 66
rect 51 59 54 61
rect 56 59 59 61
rect 51 42 59 59
rect 61 60 69 70
rect 61 58 64 60
rect 66 58 69 60
rect 61 53 69 58
rect 61 51 64 53
rect 66 51 69 53
rect 61 42 69 51
rect 71 68 79 70
rect 71 66 74 68
rect 76 66 79 68
rect 71 61 79 66
rect 71 59 74 61
rect 76 59 79 61
rect 71 42 79 59
rect 81 55 86 70
rect 81 53 88 55
rect 81 51 84 53
rect 86 51 88 53
rect 81 46 88 51
rect 81 44 84 46
rect 86 44 88 46
rect 81 42 88 44
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 2 39 6 55
rect 12 53 18 54
rect 12 51 14 53
rect 16 51 18 53
rect 12 47 18 51
rect 12 46 22 47
rect 12 44 14 46
rect 16 44 22 46
rect 12 43 22 44
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 18 22 22 43
rect 39 42 73 46
rect 26 37 30 39
rect 26 35 27 37
rect 29 35 30 37
rect 26 30 30 35
rect 39 37 45 42
rect 67 38 73 42
rect 39 35 41 37
rect 43 35 45 37
rect 39 34 45 35
rect 49 37 63 38
rect 49 35 51 37
rect 53 35 59 37
rect 61 35 63 37
rect 49 34 63 35
rect 67 37 79 38
rect 67 35 69 37
rect 71 35 79 37
rect 67 34 79 35
rect 83 37 87 39
rect 83 35 84 37
rect 86 35 87 37
rect 83 30 87 35
rect 26 26 87 30
rect 18 21 59 22
rect 18 19 55 21
rect 57 19 59 21
rect 18 18 59 19
rect 66 17 70 26
rect -2 11 98 12
rect -2 9 26 11
rect 28 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 9 22 11 30
rect 19 22 21 30
rect 33 12 35 30
rect 41 12 43 30
rect 49 12 51 30
rect 61 12 63 30
rect 69 12 71 30
rect 77 12 79 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 42 81 70
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 41 35 43 37
rect 51 35 53 37
rect 59 35 61 37
rect 69 35 71 37
rect 84 35 86 37
<< ndifct0 >>
rect 4 24 6 26
rect 14 26 16 28
rect 82 14 84 16
<< ndifct1 >>
rect 55 19 57 21
rect 26 9 28 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 60 6 62
rect 24 59 26 61
rect 24 52 26 54
rect 34 66 36 68
rect 44 59 46 61
rect 44 52 46 54
rect 54 66 56 68
rect 54 59 56 61
rect 64 58 66 60
rect 64 51 66 53
rect 74 66 76 68
rect 74 59 76 61
rect 84 51 86 53
rect 84 44 86 46
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
<< alu0 >>
rect 33 66 34 68
rect 36 66 37 68
rect 33 64 37 66
rect 52 66 54 68
rect 56 66 58 68
rect 2 62 27 63
rect 2 60 4 62
rect 6 61 27 62
rect 6 60 24 61
rect 2 59 24 60
rect 26 59 27 61
rect 23 54 27 59
rect 43 61 47 63
rect 43 59 44 61
rect 46 59 47 61
rect 43 54 47 59
rect 52 61 58 66
rect 72 66 74 68
rect 76 66 78 68
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
rect 63 60 67 62
rect 63 58 64 60
rect 66 58 67 60
rect 72 61 78 66
rect 72 59 74 61
rect 76 59 78 61
rect 72 58 78 59
rect 63 54 67 58
rect 23 52 24 54
rect 26 52 44 54
rect 46 53 88 54
rect 46 52 64 53
rect 23 51 64 52
rect 66 51 84 53
rect 86 51 88 53
rect 23 50 88 51
rect 82 46 88 50
rect 12 28 18 29
rect 3 26 7 28
rect 3 24 4 26
rect 6 24 7 26
rect 12 26 14 28
rect 16 26 18 28
rect 12 25 18 26
rect 3 12 7 24
rect 82 44 84 46
rect 86 44 88 46
rect 82 43 88 44
rect 81 16 85 18
rect 81 14 82 16
rect 84 14 85 16
rect 81 12 85 14
<< labels >>
rlabel alu0 45 56 45 56 6 n3
rlabel alu0 14 61 14 61 6 n3
rlabel alu0 25 56 25 56 6 n3
rlabel alu0 65 56 65 56 6 n3
rlabel alu0 55 52 55 52 6 n3
rlabel alu0 85 48 85 48 6 n3
rlabel alu1 4 44 4 44 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 36 20 36 6 z
rlabel polyct1 28 36 28 36 6 a1
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 44 20 44 20 6 z
rlabel alu1 44 28 44 28 6 a1
rlabel alu1 52 20 52 20 6 z
rlabel alu1 52 28 52 28 6 a1
rlabel alu1 44 44 44 44 6 a2
rlabel polyct1 52 36 52 36 6 a3
rlabel alu1 52 44 52 44 6 a2
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 60 28 60 28 6 a1
rlabel alu1 68 24 68 24 6 a1
rlabel alu1 76 28 76 28 6 a1
rlabel polyct1 60 36 60 36 6 a3
rlabel alu1 60 44 60 44 6 a2
rlabel alu1 68 44 68 44 6 a2
rlabel alu1 76 36 76 36 6 a2
rlabel alu1 84 28 84 28 6 a1
<< end >>
