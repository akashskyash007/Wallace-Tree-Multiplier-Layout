magic
tech scmos
timestamp 1199201777
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 61 11 65
rect 20 64 22 69
rect 30 64 32 69
rect 42 64 44 69
rect 52 64 54 69
rect 9 39 11 43
rect 20 39 22 58
rect 30 47 32 58
rect 42 47 44 58
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 42 45 48 47
rect 42 43 44 45
rect 46 43 48 45
rect 42 41 48 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 25 11 33
rect 22 25 24 33
rect 29 25 31 41
rect 42 36 44 41
rect 36 34 44 36
rect 52 39 54 58
rect 52 37 58 39
rect 52 35 54 37
rect 56 35 58 37
rect 36 25 38 34
rect 52 33 58 35
rect 52 30 54 33
rect 43 28 54 30
rect 43 25 45 28
rect 9 11 11 16
rect 22 12 24 17
rect 29 12 31 17
rect 36 12 38 17
rect 43 12 45 17
<< ndif >>
rect 4 22 9 25
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 17 22 25
rect 24 17 29 25
rect 31 17 36 25
rect 38 17 43 25
rect 45 23 50 25
rect 45 21 52 23
rect 45 19 48 21
rect 50 19 52 21
rect 45 17 52 19
rect 11 16 20 17
rect 13 11 20 16
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 34 71 40 73
rect 34 69 36 71
rect 38 69 40 71
rect 34 64 40 69
rect 13 62 20 64
rect 13 61 15 62
rect 4 56 9 61
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 60 15 61
rect 17 60 20 62
rect 11 58 20 60
rect 22 62 30 64
rect 22 60 25 62
rect 27 60 30 62
rect 22 58 30 60
rect 32 58 42 64
rect 44 62 52 64
rect 44 60 47 62
rect 49 60 52 62
rect 44 58 52 60
rect 54 62 61 64
rect 54 60 57 62
rect 59 60 61 62
rect 54 58 61 60
rect 11 43 18 58
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 36 71
rect 38 69 66 71
rect -2 68 66 69
rect 2 54 7 63
rect 2 52 4 54
rect 6 52 7 54
rect 2 47 7 52
rect 2 45 4 47
rect 6 45 7 47
rect 2 43 7 45
rect 33 50 47 54
rect 2 22 6 43
rect 33 46 37 50
rect 58 46 62 55
rect 25 45 37 46
rect 25 43 31 45
rect 33 43 37 45
rect 25 42 37 43
rect 41 45 62 46
rect 41 43 44 45
rect 46 43 62 45
rect 41 42 62 43
rect 19 37 31 38
rect 19 35 21 37
rect 23 35 31 37
rect 19 34 31 35
rect 41 37 62 38
rect 41 35 54 37
rect 56 35 62 37
rect 41 34 62 35
rect 27 30 31 34
rect 27 26 47 30
rect 2 20 15 22
rect 2 18 4 20
rect 6 18 15 20
rect 2 17 15 18
rect 58 17 62 34
rect -2 11 66 12
rect -2 9 15 11
rect 17 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 16 11 25
rect 22 17 24 25
rect 29 17 31 25
rect 36 17 38 25
rect 43 17 45 25
<< pmos >>
rect 9 43 11 61
rect 20 58 22 64
rect 30 58 32 64
rect 42 58 44 64
rect 52 58 54 64
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 44 43 46 45
rect 21 35 23 37
rect 54 35 56 37
<< ndifct0 >>
rect 48 19 50 21
<< ndifct1 >>
rect 4 18 6 20
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 15 60 17 62
rect 25 60 27 62
rect 47 60 49 62
rect 57 60 59 62
<< pdifct1 >>
rect 36 69 38 71
rect 4 52 6 54
rect 4 45 6 47
<< alu0 >>
rect 14 62 18 68
rect 14 60 15 62
rect 17 60 18 62
rect 14 58 18 60
rect 23 62 51 63
rect 23 60 25 62
rect 27 60 47 62
rect 49 60 51 62
rect 23 59 51 60
rect 55 62 61 68
rect 55 60 57 62
rect 59 60 61 62
rect 55 59 61 60
rect 23 54 27 59
rect 11 50 27 54
rect 11 39 15 50
rect 10 37 15 39
rect 10 35 11 37
rect 13 35 15 37
rect 10 33 15 35
rect 11 30 15 33
rect 11 26 23 30
rect 19 22 23 26
rect 19 21 52 22
rect 19 19 48 21
rect 50 19 52 21
rect 19 18 52 19
<< labels >>
rlabel alu0 13 40 13 40 6 zn
rlabel alu0 35 20 35 20 6 zn
rlabel alu0 37 61 37 61 6 zn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 36 28 36 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 36 44 36 6 d
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 44 44 44 6 c
rlabel alu1 36 52 36 52 6 b
rlabel alu1 44 52 44 52 6 b
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 36 52 36 6 d
rlabel alu1 60 24 60 24 6 d
rlabel alu1 52 44 52 44 6 c
rlabel alu1 60 52 60 52 6 c
<< end >>
