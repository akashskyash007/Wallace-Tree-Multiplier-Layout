magic
tech scmos
timestamp 1199201931
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 31 66 33 71
rect 41 66 43 71
rect 9 57 11 62
rect 19 57 21 62
rect 31 48 33 51
rect 31 46 37 48
rect 31 44 33 46
rect 35 44 37 46
rect 9 38 11 43
rect 19 40 21 43
rect 31 42 37 44
rect 19 38 27 40
rect 9 36 15 38
rect 9 34 11 36
rect 13 34 15 36
rect 21 36 23 38
rect 25 36 27 38
rect 21 34 27 36
rect 9 32 17 34
rect 15 29 17 32
rect 22 29 24 34
rect 34 30 36 42
rect 41 39 43 51
rect 41 37 47 39
rect 41 35 43 37
rect 45 35 47 37
rect 41 33 47 35
rect 41 30 43 33
rect 15 12 17 17
rect 22 12 24 17
rect 34 12 36 17
rect 41 12 43 17
<< ndif >>
rect 26 29 34 30
rect 10 23 15 29
rect 8 21 15 23
rect 8 19 10 21
rect 12 19 15 21
rect 8 17 15 19
rect 17 17 22 29
rect 24 17 34 29
rect 36 17 41 30
rect 43 23 48 30
rect 43 21 50 23
rect 43 19 46 21
rect 48 19 50 21
rect 43 17 50 19
rect 26 11 32 17
rect 26 9 28 11
rect 30 9 32 11
rect 26 7 32 9
<< pdif >>
rect 23 71 29 73
rect 23 69 25 71
rect 27 69 29 71
rect 23 66 29 69
rect 23 57 31 66
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 43 9 53
rect 11 54 19 57
rect 11 52 14 54
rect 16 52 19 54
rect 11 47 19 52
rect 11 45 14 47
rect 16 45 19 47
rect 11 43 19 45
rect 21 51 31 57
rect 33 61 41 66
rect 33 59 36 61
rect 38 59 41 61
rect 33 51 41 59
rect 43 64 50 66
rect 43 62 46 64
rect 48 62 50 64
rect 43 56 50 62
rect 43 54 46 56
rect 48 54 50 56
rect 43 51 50 54
rect 21 43 29 51
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 25 71
rect 27 69 58 71
rect -2 68 58 69
rect 13 54 17 56
rect 13 52 14 54
rect 16 52 17 54
rect 13 47 17 52
rect 2 45 14 47
rect 16 45 17 47
rect 2 43 17 45
rect 2 23 6 43
rect 33 48 39 54
rect 32 46 39 48
rect 32 44 33 46
rect 35 44 47 46
rect 32 42 47 44
rect 10 36 14 39
rect 10 34 11 36
rect 13 34 14 36
rect 10 31 14 34
rect 10 27 22 31
rect 2 21 14 23
rect 2 19 10 21
rect 12 19 14 21
rect 2 17 14 19
rect 18 17 22 27
rect 34 37 47 38
rect 34 35 43 37
rect 45 35 47 37
rect 34 34 47 35
rect 34 25 38 34
rect -2 11 58 12
rect -2 9 28 11
rect 30 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 15 17 17 29
rect 22 17 24 29
rect 34 17 36 30
rect 41 17 43 30
<< pmos >>
rect 9 43 11 57
rect 19 43 21 57
rect 31 51 33 66
rect 41 51 43 66
<< polyct0 >>
rect 23 36 25 38
<< polyct1 >>
rect 33 44 35 46
rect 11 34 13 36
rect 43 35 45 37
<< ndifct0 >>
rect 46 19 48 21
<< ndifct1 >>
rect 10 19 12 21
rect 28 9 30 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 53 6 55
rect 36 59 38 61
rect 46 62 48 64
rect 46 54 48 56
<< pdifct1 >>
rect 25 69 27 71
rect 14 52 16 54
rect 14 45 16 47
<< alu0 >>
rect 3 55 7 68
rect 45 64 49 68
rect 45 62 46 64
rect 48 62 49 64
rect 23 61 40 62
rect 23 59 36 61
rect 38 59 40 61
rect 23 58 40 59
rect 3 53 4 55
rect 6 53 7 55
rect 3 51 7 53
rect 23 39 27 58
rect 45 56 49 62
rect 45 54 46 56
rect 48 54 49 56
rect 45 52 49 54
rect 19 38 30 39
rect 19 36 23 38
rect 25 36 30 38
rect 19 35 30 36
rect 26 22 30 35
rect 26 21 50 22
rect 26 19 46 21
rect 48 19 50 21
rect 26 18 50 19
<< labels >>
rlabel polyct0 24 37 24 37 6 an
rlabel alu0 31 60 31 60 6 an
rlabel alu0 38 20 38 20 6 an
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 36 12 36 6 b
rlabel alu1 20 24 20 24 6 b
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 36 48 36 48 6 a2
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 36 44 36 6 a1
rlabel alu1 44 44 44 44 6 a2
<< end >>
