magic
tech scmos
timestamp 1199471927
<< ab >>
rect 0 0 30 100
<< nwell >>
rect -5 48 35 105
<< pwell >>
rect -5 -5 35 48
<< poly >>
rect 19 85 21 89
rect 19 73 21 76
rect 9 71 15 73
rect 9 69 11 71
rect 13 69 15 71
rect 9 67 15 69
rect 19 71 26 73
rect 19 69 21 71
rect 23 69 26 71
rect 19 67 26 69
rect 11 64 13 67
rect 11 39 13 55
rect 11 30 13 33
rect 9 28 15 30
rect 9 26 11 28
rect 13 26 15 28
rect 24 27 26 67
rect 9 24 15 26
rect 19 25 26 27
rect 19 22 21 25
rect 19 11 21 16
<< ndif >>
rect 3 37 11 39
rect 3 35 5 37
rect 7 35 11 37
rect 3 33 11 35
rect 13 37 22 39
rect 13 35 18 37
rect 20 35 22 37
rect 13 33 22 35
rect 10 20 19 22
rect 10 18 12 20
rect 14 18 19 20
rect 10 16 19 18
rect 21 16 27 22
rect 23 9 27 16
rect 21 7 27 9
rect 21 5 23 7
rect 25 5 27 7
rect 21 3 27 5
<< pdif >>
rect 21 95 27 97
rect 21 93 23 95
rect 25 93 27 95
rect 21 91 27 93
rect 23 85 27 91
rect 14 82 19 85
rect 9 80 19 82
rect 9 78 11 80
rect 13 78 19 80
rect 9 76 19 78
rect 21 76 27 85
rect 3 62 11 64
rect 3 60 5 62
rect 7 60 11 62
rect 3 58 11 60
rect 6 55 11 58
rect 13 61 18 64
rect 13 59 21 61
rect 13 57 17 59
rect 19 57 21 59
rect 13 55 21 57
<< alu1 >>
rect -2 95 32 100
rect -2 93 9 95
rect 11 93 23 95
rect 25 93 32 95
rect -2 88 32 93
rect 2 63 6 88
rect 10 80 14 82
rect 10 78 11 80
rect 13 78 14 80
rect 10 71 14 78
rect 10 69 11 71
rect 13 69 14 71
rect 10 67 14 69
rect 18 73 22 83
rect 18 71 25 73
rect 18 69 21 71
rect 23 69 25 71
rect 18 67 25 69
rect 2 62 9 63
rect 2 60 5 62
rect 7 60 9 62
rect 2 58 9 60
rect 16 59 22 63
rect 16 57 17 59
rect 19 57 22 59
rect 16 52 22 57
rect 7 48 22 52
rect 2 37 9 39
rect 2 35 5 37
rect 7 35 9 37
rect 2 34 9 35
rect 16 37 22 48
rect 16 35 18 37
rect 20 35 22 37
rect 16 34 22 35
rect 2 12 6 34
rect 10 28 16 30
rect 10 26 11 28
rect 13 26 16 28
rect 10 20 16 26
rect 10 18 12 20
rect 14 18 16 20
rect 10 17 16 18
rect -2 7 32 12
rect -2 5 9 7
rect 11 5 23 7
rect 25 5 32 7
rect -2 0 32 5
<< ptie >>
rect 7 7 13 9
rect 7 5 9 7
rect 11 5 13 7
rect 7 3 13 5
<< ntie >>
rect 7 95 13 97
rect 7 93 9 95
rect 11 93 13 95
rect 7 91 13 93
<< nmos >>
rect 11 33 13 39
rect 19 16 21 22
<< pmos >>
rect 19 76 21 85
rect 11 55 13 64
<< polyct1 >>
rect 11 69 13 71
rect 21 69 23 71
rect 11 26 13 28
<< ndifct1 >>
rect 5 35 7 37
rect 18 35 20 37
rect 12 18 14 20
rect 23 5 25 7
<< ntiect1 >>
rect 9 93 11 95
<< ptiect1 >>
rect 9 5 11 7
<< pdifct1 >>
rect 23 93 25 95
rect 11 78 13 80
rect 5 60 7 62
rect 17 57 19 59
<< labels >>
rlabel polyct1 12 27 12 27 6 an
rlabel ndifct1 13 19 13 19 6 an
rlabel pdifct1 12 79 12 79 6 an
rlabel polyct1 12 70 12 70 6 an
rlabel alu1 10 50 10 50 6 z
rlabel alu1 15 6 15 6 6 vss
rlabel alu1 20 50 20 50 6 z
rlabel alu1 20 75 20 75 6 a
rlabel alu1 15 94 15 94 6 vdd
<< end >>
