magic
tech scmos
timestamp 1199203229
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 60 48 65
rect 53 60 55 65
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 21 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 35 31 44
rect 36 41 38 44
rect 46 41 48 44
rect 36 39 48 41
rect 53 41 55 44
rect 53 39 62 41
rect 41 37 48 39
rect 41 35 43 37
rect 45 35 48 37
rect 56 37 58 39
rect 60 37 62 39
rect 56 35 62 37
rect 29 33 37 35
rect 29 32 33 33
rect 31 31 33 32
rect 35 31 37 33
rect 31 29 37 31
rect 41 33 48 35
rect 31 26 33 29
rect 41 26 43 33
rect 9 11 11 16
rect 19 11 21 16
rect 31 9 33 14
rect 41 9 43 14
<< ndif >>
rect 2 20 9 30
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 16 19 19
rect 21 26 28 30
rect 21 16 31 26
rect 23 14 31 16
rect 33 21 41 26
rect 33 19 36 21
rect 38 19 41 21
rect 33 14 41 19
rect 43 18 51 26
rect 43 16 46 18
rect 48 16 51 18
rect 43 14 51 16
rect 23 11 29 14
rect 23 9 25 11
rect 27 9 29 11
rect 23 7 29 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 54 19 70
rect 11 52 14 54
rect 16 52 19 54
rect 11 46 19 52
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 44 29 59
rect 31 44 36 70
rect 38 60 43 70
rect 38 53 46 60
rect 38 51 41 53
rect 43 51 46 53
rect 38 44 46 51
rect 48 44 53 60
rect 55 58 62 60
rect 55 56 58 58
rect 60 56 62 58
rect 55 44 62 56
rect 21 42 27 44
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 13 54 17 56
rect 13 52 14 54
rect 16 52 17 54
rect 13 47 17 52
rect 2 46 17 47
rect 2 44 14 46
rect 16 44 17 46
rect 2 42 17 44
rect 2 30 6 42
rect 58 46 62 47
rect 2 28 17 30
rect 2 26 14 28
rect 16 26 17 28
rect 2 25 17 26
rect 13 21 17 25
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect 32 42 62 46
rect 32 33 36 42
rect 32 31 33 33
rect 35 31 36 33
rect 32 29 36 31
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 31 47 35
rect 58 39 62 42
rect 60 37 62 39
rect 58 33 62 37
rect 41 25 54 31
rect -2 11 66 12
rect -2 9 25 11
rect 27 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 31 14 33 26
rect 41 14 43 26
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 44 31 70
rect 36 44 38 70
rect 46 44 48 60
rect 53 44 55 60
<< polyct0 >>
rect 17 35 19 37
<< polyct1 >>
rect 43 35 45 37
rect 58 37 60 39
rect 33 31 35 33
<< ndifct0 >>
rect 4 18 6 20
rect 36 19 38 21
rect 46 16 48 18
<< ndifct1 >>
rect 14 26 16 28
rect 14 19 16 21
rect 25 9 27 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 66 26 68
rect 24 59 26 61
rect 41 51 43 53
rect 58 56 60 58
<< pdifct1 >>
rect 14 52 16 54
rect 14 44 16 46
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 57 58 61 68
rect 57 56 58 58
rect 60 56 61 58
rect 57 54 61 56
rect 23 53 45 54
rect 23 51 41 53
rect 43 51 45 53
rect 23 50 45 51
rect 23 38 27 50
rect 15 37 27 38
rect 15 35 17 37
rect 19 35 27 37
rect 15 34 27 35
rect 2 20 8 21
rect 2 18 4 20
rect 6 18 8 20
rect 2 12 8 18
rect 23 22 27 34
rect 57 33 58 42
rect 23 21 40 22
rect 23 19 36 21
rect 38 19 40 21
rect 23 18 40 19
rect 45 18 49 20
rect 45 16 46 18
rect 48 16 49 18
rect 45 12 49 16
<< labels >>
rlabel alu0 21 36 21 36 6 zn
rlabel alu0 31 20 31 20 6 zn
rlabel alu0 34 52 34 52 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 32 44 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 b
rlabel alu1 60 40 60 40 6 a
rlabel alu1 52 44 52 44 6 a
<< end >>
