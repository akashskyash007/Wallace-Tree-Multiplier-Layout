magic
tech scmos
timestamp 1199202591
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 10 57 12 62
rect 20 57 22 61
rect 10 35 12 43
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 9 19 11 29
rect 20 28 22 43
rect 20 26 26 28
rect 20 24 22 26
rect 24 24 26 26
rect 16 22 26 24
rect 16 19 18 22
rect 9 2 11 7
rect 16 2 18 7
<< ndif >>
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 7 9 13
rect 11 7 16 19
rect 18 11 30 19
rect 18 9 26 11
rect 28 9 30 11
rect 18 7 30 9
<< pdif >>
rect 2 57 8 59
rect 2 55 4 57
rect 6 55 10 57
rect 2 43 10 55
rect 12 55 20 57
rect 12 53 15 55
rect 17 53 20 55
rect 12 48 20 53
rect 12 46 15 48
rect 17 46 20 48
rect 12 43 20 46
rect 22 55 30 57
rect 22 53 26 55
rect 28 53 30 55
rect 22 48 30 53
rect 22 46 26 48
rect 28 46 30 48
rect 22 43 30 46
<< alu1 >>
rect -2 67 34 72
rect -2 65 17 67
rect 19 65 25 67
rect 27 65 34 67
rect -2 64 34 65
rect 2 46 15 50
rect 2 19 6 46
rect 17 38 23 42
rect 10 34 23 38
rect 10 33 14 34
rect 10 31 11 33
rect 13 31 14 33
rect 10 29 14 31
rect 18 26 30 27
rect 18 24 22 26
rect 24 24 30 26
rect 18 21 30 24
rect 2 17 7 19
rect 2 15 4 17
rect 6 15 7 17
rect 2 13 7 15
rect 18 13 22 21
rect -2 0 34 8
<< ntie >>
rect 15 67 29 69
rect 15 65 17 67
rect 19 65 25 67
rect 27 65 29 67
rect 15 63 29 65
<< nmos >>
rect 9 7 11 19
rect 16 7 18 19
<< pmos >>
rect 10 43 12 57
rect 20 43 22 57
<< polyct1 >>
rect 11 31 13 33
rect 22 24 24 26
<< ndifct0 >>
rect 26 9 28 11
<< ndifct1 >>
rect 4 15 6 17
<< ntiect1 >>
rect 17 65 19 67
rect 25 65 27 67
<< pdifct0 >>
rect 4 55 6 57
rect 15 53 17 55
rect 15 46 17 48
rect 26 53 28 55
rect 26 46 28 48
<< alu0 >>
rect 2 57 8 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 55 19 56
rect 13 53 15 55
rect 17 53 19 55
rect 13 50 19 53
rect 15 48 19 50
rect 17 46 19 48
rect 6 45 19 46
rect 24 55 30 64
rect 24 53 26 55
rect 28 53 30 55
rect 24 48 30 53
rect 24 46 26 48
rect 28 46 30 48
rect 24 45 30 46
rect 25 11 29 13
rect 25 9 26 11
rect 28 9 29 11
rect 25 8 29 9
<< labels >>
rlabel alu1 4 28 4 28 6 z
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 12 48 12 48 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 20 20 20 6 a
rlabel alu1 20 40 20 40 6 b
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 24 28 24 6 a
<< end >>
