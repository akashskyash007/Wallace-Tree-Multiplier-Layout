magic
tech scmos
timestamp 1199201684
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 60 11 65
rect 19 56 21 61
rect 29 56 31 61
rect 9 39 11 42
rect 19 39 21 50
rect 29 47 31 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 28 11 33
rect 22 23 24 33
rect 29 23 31 41
rect 9 15 11 19
rect 22 12 24 17
rect 29 12 31 17
<< ndif >>
rect 4 25 9 28
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 23 20 28
rect 11 19 22 23
rect 13 17 22 19
rect 24 17 29 23
rect 31 21 38 23
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
rect 13 11 20 17
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 13 67 19 69
rect 13 65 15 67
rect 17 65 19 67
rect 13 63 19 65
rect 32 67 38 69
rect 32 65 34 67
rect 36 65 38 67
rect 32 63 38 65
rect 13 60 17 63
rect 4 55 9 60
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 56 17 60
rect 33 56 38 63
rect 11 50 19 56
rect 21 54 29 56
rect 21 52 24 54
rect 26 52 29 54
rect 21 50 29 52
rect 31 50 38 56
rect 11 42 17 50
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 2 23 6 42
rect 34 46 38 55
rect 25 45 38 46
rect 25 43 31 45
rect 33 43 38 45
rect 25 42 38 43
rect 17 37 31 38
rect 17 35 21 37
rect 23 35 31 37
rect 17 34 31 35
rect 25 26 31 34
rect 2 21 4 23
rect 6 21 14 23
rect 2 17 14 21
rect -2 11 42 12
rect -2 9 15 11
rect 17 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 19 11 28
rect 22 17 24 23
rect 29 17 31 23
<< pmos >>
rect 9 42 11 60
rect 19 50 21 56
rect 29 50 31 56
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 21 35 23 37
<< ndifct0 >>
rect 34 19 36 21
<< ndifct1 >>
rect 4 21 6 23
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 15 65 17 67
rect 34 65 36 67
rect 24 52 26 54
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 14 67 18 68
rect 14 65 15 67
rect 17 65 18 67
rect 14 63 18 65
rect 33 67 37 68
rect 33 65 34 67
rect 36 65 37 67
rect 33 63 37 65
rect 10 54 28 55
rect 10 52 24 54
rect 26 52 28 54
rect 10 51 28 52
rect 10 37 14 51
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 10 26 22 30
rect 6 23 7 25
rect 18 22 22 26
rect 18 21 38 22
rect 18 19 34 21
rect 36 19 38 21
rect 18 18 38 19
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 19 53 19 53 6 zn
rlabel alu0 28 20 28 20 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 52 36 52 6 b
<< end >>
