magic
tech scmos
timestamp 1199203588
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 61 70 63 74
rect 71 70 73 74
rect 29 63 31 68
rect 39 63 41 68
rect 48 46 54 48
rect 48 44 50 46
rect 52 44 54 46
rect 48 42 54 44
rect 81 63 83 68
rect 91 63 93 68
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 48 39 50 42
rect 9 37 25 39
rect 29 37 50 39
rect 61 39 63 42
rect 71 39 73 42
rect 81 39 83 42
rect 91 39 93 42
rect 61 37 73 39
rect 78 37 103 39
rect 16 35 21 37
rect 23 35 25 37
rect 16 33 25 35
rect 9 28 11 33
rect 16 31 28 33
rect 16 28 18 31
rect 26 28 28 31
rect 33 28 35 37
rect 65 35 67 37
rect 69 35 71 37
rect 65 33 71 35
rect 78 33 80 37
rect 97 35 99 37
rect 101 35 103 37
rect 97 33 103 35
rect 65 28 67 33
rect 75 31 80 33
rect 75 28 77 31
rect 85 29 91 31
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
rect 85 27 87 29
rect 89 27 91 29
rect 85 25 97 27
rect 85 22 87 25
rect 95 22 97 25
rect 65 6 67 10
rect 75 6 77 10
rect 85 8 87 13
rect 95 8 97 13
<< ndif >>
rect 2 20 9 28
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 16 28
rect 18 26 26 28
rect 18 24 21 26
rect 23 24 26 26
rect 18 16 26 24
rect 28 16 33 28
rect 35 16 44 28
rect 60 23 65 28
rect 58 21 65 23
rect 58 19 60 21
rect 62 19 65 21
rect 58 17 65 19
rect 37 11 44 16
rect 37 9 39 11
rect 41 9 44 11
rect 60 10 65 17
rect 67 26 75 28
rect 67 24 70 26
rect 72 24 75 26
rect 67 10 75 24
rect 77 22 83 28
rect 77 17 85 22
rect 77 15 80 17
rect 82 15 85 17
rect 77 13 85 15
rect 87 20 95 22
rect 87 18 90 20
rect 92 18 95 20
rect 87 13 95 18
rect 97 13 105 22
rect 77 10 83 13
rect 37 7 44 9
rect 99 11 105 13
rect 99 9 101 11
rect 103 9 105 11
rect 99 7 105 9
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 63 26 70
rect 54 68 61 70
rect 54 66 56 68
rect 58 66 61 68
rect 21 61 29 63
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 46 39 63
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 61 48 63
rect 41 59 44 61
rect 46 59 48 61
rect 41 57 48 59
rect 54 61 61 66
rect 54 59 56 61
rect 58 59 61 61
rect 54 57 61 59
rect 41 42 46 57
rect 56 42 61 57
rect 63 60 71 70
rect 63 58 66 60
rect 68 58 71 60
rect 63 53 71 58
rect 63 51 66 53
rect 68 51 71 53
rect 63 42 71 51
rect 73 63 79 70
rect 73 61 81 63
rect 73 59 76 61
rect 78 59 81 61
rect 73 42 81 59
rect 83 46 91 63
rect 83 44 86 46
rect 88 44 91 46
rect 83 42 91 44
rect 93 61 100 63
rect 93 59 96 61
rect 98 59 100 61
rect 93 42 100 59
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 68 114 79
rect 2 61 48 62
rect 2 59 4 61
rect 6 59 24 61
rect 26 59 44 61
rect 46 59 48 61
rect 2 58 48 59
rect 2 54 7 58
rect 2 52 4 54
rect 6 52 7 54
rect 2 50 7 52
rect 2 30 6 50
rect 97 38 103 46
rect 65 37 82 38
rect 65 35 67 37
rect 69 35 82 37
rect 65 34 82 35
rect 89 37 103 38
rect 89 35 99 37
rect 101 35 103 37
rect 89 34 103 35
rect 78 30 82 34
rect 2 26 24 30
rect 78 29 91 30
rect 78 27 87 29
rect 89 27 91 29
rect 78 26 91 27
rect 20 24 21 26
rect 23 24 24 26
rect 20 22 24 24
rect 20 21 64 22
rect 20 19 60 21
rect 62 19 64 21
rect 20 18 64 19
rect -2 11 114 12
rect -2 9 39 11
rect 41 9 101 11
rect 103 9 114 11
rect -2 1 114 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 9 16 11 28
rect 16 16 18 28
rect 26 16 28 28
rect 33 16 35 28
rect 65 10 67 28
rect 75 10 77 28
rect 85 13 87 22
rect 95 13 97 22
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 63
rect 39 42 41 63
rect 61 42 63 70
rect 71 42 73 70
rect 81 42 83 63
rect 91 42 93 63
<< polyct0 >>
rect 50 44 52 46
rect 21 35 23 37
<< polyct1 >>
rect 67 35 69 37
rect 99 35 101 37
rect 87 27 89 29
<< ndifct0 >>
rect 4 18 6 20
rect 70 24 72 26
rect 80 15 82 17
rect 90 18 92 20
<< ndifct1 >>
rect 21 24 23 26
rect 60 19 62 21
rect 39 9 41 11
rect 101 9 103 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 14 51 16 53
rect 14 44 16 46
rect 56 66 58 68
rect 34 44 36 46
rect 56 59 58 61
rect 66 58 68 60
rect 66 51 68 53
rect 76 59 78 61
rect 86 44 88 46
rect 96 59 98 61
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
rect 24 59 26 61
rect 44 59 46 61
<< alu0 >>
rect 54 66 56 68
rect 58 66 60 68
rect 54 61 60 66
rect 54 59 56 61
rect 58 59 60 61
rect 54 58 60 59
rect 65 60 69 62
rect 65 58 66 60
rect 68 58 69 60
rect 74 61 80 68
rect 74 59 76 61
rect 78 59 80 61
rect 74 58 80 59
rect 94 61 100 68
rect 94 59 96 61
rect 98 59 100 61
rect 94 58 100 59
rect 65 54 69 58
rect 12 53 110 54
rect 12 51 14 53
rect 16 51 66 53
rect 68 51 110 53
rect 12 50 110 51
rect 12 46 17 50
rect 12 44 14 46
rect 16 44 17 46
rect 12 42 17 44
rect 32 46 38 47
rect 32 44 34 46
rect 36 44 38 46
rect 32 38 38 44
rect 49 46 53 50
rect 84 46 90 47
rect 49 44 50 46
rect 52 44 53 46
rect 49 42 53 44
rect 57 44 86 46
rect 88 44 90 46
rect 57 42 90 44
rect 57 38 61 42
rect 19 37 61 38
rect 19 35 21 37
rect 23 35 61 37
rect 19 34 61 35
rect 57 30 61 34
rect 57 26 73 30
rect 69 24 70 26
rect 72 24 73 26
rect 69 22 73 24
rect 3 20 7 22
rect 3 18 4 20
rect 6 18 7 20
rect 106 21 110 50
rect 88 20 110 21
rect 3 12 7 18
rect 79 17 83 19
rect 88 18 90 20
rect 92 18 110 20
rect 88 17 110 18
rect 79 15 80 17
rect 82 15 83 17
rect 79 12 83 15
<< labels >>
rlabel alu0 14 48 14 48 6 bn
rlabel alu0 51 48 51 48 6 bn
rlabel alu0 35 40 35 40 6 an
rlabel alu0 40 36 40 36 6 an
rlabel alu0 71 26 71 26 6 an
rlabel alu0 67 56 67 56 6 bn
rlabel alu0 99 19 99 19 6 bn
rlabel alu0 73 44 73 44 6 an
rlabel alu0 61 52 61 52 6 bn
rlabel alu1 20 28 20 28 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 56 6 56 6 6 vss
rlabel alu1 60 20 60 20 6 z
rlabel alu1 76 36 76 36 6 b
rlabel polyct1 68 36 68 36 6 b
rlabel alu1 56 74 56 74 6 vdd
rlabel alu1 84 28 84 28 6 b
rlabel alu1 92 36 92 36 6 a
rlabel alu1 100 40 100 40 6 a
<< end >>
