magic
tech scmos
timestamp 1199541572
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 35 94 37 98
rect 47 94 49 98
rect 11 86 13 90
rect 23 85 25 89
rect 11 63 13 66
rect 7 61 13 63
rect 7 59 9 61
rect 11 59 13 61
rect 7 57 13 59
rect 23 53 25 65
rect 23 51 31 53
rect 23 49 27 51
rect 29 49 31 51
rect 23 47 31 49
rect 17 41 23 43
rect 35 41 37 55
rect 47 41 49 55
rect 17 39 19 41
rect 21 39 49 41
rect 17 37 23 39
rect 7 31 13 33
rect 7 29 9 31
rect 11 29 13 31
rect 7 27 13 29
rect 11 24 13 27
rect 23 31 31 33
rect 23 29 27 31
rect 29 29 31 31
rect 23 27 31 29
rect 23 24 25 27
rect 35 25 37 39
rect 47 25 49 39
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
<< ndif >>
rect 30 24 35 25
rect 3 21 11 24
rect 3 19 5 21
rect 7 19 11 21
rect 3 6 11 19
rect 13 6 23 24
rect 25 11 35 24
rect 25 9 29 11
rect 31 9 35 11
rect 25 6 35 9
rect 37 21 47 25
rect 37 19 41 21
rect 43 19 47 21
rect 37 6 47 19
rect 49 21 57 25
rect 49 19 53 21
rect 55 19 57 21
rect 49 11 57 19
rect 49 9 53 11
rect 55 9 57 11
rect 49 6 57 9
<< pdif >>
rect 3 91 9 93
rect 3 89 5 91
rect 7 89 9 91
rect 27 91 35 94
rect 3 86 9 89
rect 27 89 29 91
rect 31 89 35 91
rect 3 81 11 86
rect 3 79 5 81
rect 7 79 11 81
rect 3 66 11 79
rect 13 85 21 86
rect 27 85 35 89
rect 13 81 23 85
rect 13 79 17 81
rect 19 79 23 81
rect 13 66 23 79
rect 18 65 23 66
rect 25 65 35 85
rect 27 55 35 65
rect 37 81 47 94
rect 37 79 41 81
rect 43 79 47 81
rect 37 71 47 79
rect 37 69 41 71
rect 43 69 47 71
rect 37 61 47 69
rect 37 59 41 61
rect 43 59 47 61
rect 37 55 47 59
rect 49 91 57 94
rect 49 89 53 91
rect 55 89 57 91
rect 49 81 57 89
rect 49 79 53 81
rect 55 79 57 81
rect 49 71 57 79
rect 49 69 53 71
rect 55 69 57 71
rect 49 61 57 69
rect 49 59 53 61
rect 55 59 57 61
rect 49 55 57 59
<< alu1 >>
rect -2 91 62 100
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 53 91
rect 55 89 62 91
rect -2 88 62 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 77 8 79
rect 15 81 21 82
rect 15 79 17 81
rect 19 79 21 81
rect 15 78 21 79
rect 8 61 12 73
rect 8 59 9 61
rect 11 59 12 61
rect 8 31 12 59
rect 8 29 9 31
rect 11 29 12 31
rect 8 27 12 29
rect 17 42 21 78
rect 28 52 32 83
rect 25 51 32 52
rect 25 49 27 51
rect 29 49 32 51
rect 25 48 32 49
rect 17 41 23 42
rect 17 39 19 41
rect 21 39 23 41
rect 17 38 23 39
rect 17 22 21 38
rect 28 32 32 48
rect 25 31 32 32
rect 25 29 27 31
rect 29 29 32 31
rect 25 28 32 29
rect 3 21 21 22
rect 3 19 5 21
rect 7 19 21 21
rect 3 18 21 19
rect 28 17 32 28
rect 38 82 42 83
rect 38 81 45 82
rect 38 79 41 81
rect 43 79 45 81
rect 38 78 45 79
rect 52 81 56 88
rect 52 79 53 81
rect 55 79 56 81
rect 38 72 42 78
rect 38 71 45 72
rect 38 69 41 71
rect 43 69 45 71
rect 38 68 45 69
rect 52 71 56 79
rect 52 69 53 71
rect 55 69 56 71
rect 38 62 42 68
rect 38 61 45 62
rect 38 59 41 61
rect 43 59 45 61
rect 38 58 45 59
rect 52 61 56 69
rect 52 59 53 61
rect 55 59 56 61
rect 38 22 42 58
rect 52 57 56 59
rect 38 21 45 22
rect 38 19 41 21
rect 43 19 45 21
rect 38 18 45 19
rect 52 21 56 23
rect 52 19 53 21
rect 55 19 56 21
rect 38 17 42 18
rect 52 12 56 19
rect -2 11 62 12
rect -2 9 29 11
rect 31 9 53 11
rect 55 9 62 11
rect -2 0 62 9
<< nmos >>
rect 11 6 13 24
rect 23 6 25 24
rect 35 6 37 25
rect 47 6 49 25
<< pmos >>
rect 11 66 13 86
rect 23 65 25 85
rect 35 55 37 94
rect 47 55 49 94
<< polyct1 >>
rect 9 59 11 61
rect 27 49 29 51
rect 19 39 21 41
rect 9 29 11 31
rect 27 29 29 31
<< ndifct1 >>
rect 5 19 7 21
rect 29 9 31 11
rect 41 19 43 21
rect 53 19 55 21
rect 53 9 55 11
<< pdifct1 >>
rect 5 89 7 91
rect 29 89 31 91
rect 5 79 7 81
rect 17 79 19 81
rect 41 79 43 81
rect 41 69 43 71
rect 41 59 43 61
rect 53 89 55 91
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
<< labels >>
rlabel alu1 10 50 10 50 6 i0
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 40 50 40 50 6 q
rlabel alu1 30 50 30 50 6 i1
rlabel alu1 30 94 30 94 6 vdd
<< end >>
