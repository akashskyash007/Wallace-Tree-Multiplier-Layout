magic
tech scmos
timestamp 1199543874
<< ab >>
rect 0 0 240 100
<< nwell >>
rect -2 48 242 104
<< pwell >>
rect -2 -4 242 48
<< poly >>
rect 119 95 121 98
rect 155 95 157 98
rect 167 95 169 98
rect 179 95 181 98
rect 191 95 193 98
rect 203 95 205 98
rect 215 95 217 98
rect 227 95 229 98
rect 11 85 13 88
rect 23 85 25 88
rect 31 85 33 88
rect 49 85 51 88
rect 57 85 59 88
rect 83 85 85 88
rect 95 85 97 88
rect 131 85 133 88
rect 143 85 145 88
rect 119 73 121 75
rect 115 71 121 73
rect 115 69 117 71
rect 119 69 121 71
rect 115 67 121 69
rect 155 73 157 75
rect 155 71 163 73
rect 155 69 159 71
rect 161 69 163 71
rect 155 67 163 69
rect 11 51 13 65
rect 23 63 25 65
rect 17 61 25 63
rect 17 59 19 61
rect 21 59 25 61
rect 17 57 25 59
rect 31 53 33 65
rect 49 63 51 65
rect 57 63 59 65
rect 83 63 85 65
rect 47 61 53 63
rect 47 59 49 61
rect 51 59 53 61
rect 47 57 53 59
rect 57 61 63 63
rect 57 59 59 61
rect 61 59 63 61
rect 57 57 63 59
rect 83 61 91 63
rect 83 59 87 61
rect 89 59 91 61
rect 83 57 91 59
rect 27 51 33 53
rect 77 51 83 53
rect 95 51 97 65
rect 131 63 133 65
rect 127 61 133 63
rect 127 59 129 61
rect 131 59 133 61
rect 127 57 133 59
rect 127 51 133 53
rect 143 51 145 65
rect 167 63 169 75
rect 161 61 169 63
rect 161 59 163 61
rect 165 59 169 61
rect 161 57 169 59
rect 179 51 181 75
rect 191 73 193 75
rect 185 71 193 73
rect 185 69 187 71
rect 189 69 193 71
rect 185 67 193 69
rect 203 53 205 75
rect 203 51 211 53
rect 11 49 29 51
rect 31 49 51 51
rect 11 25 13 49
rect 27 47 33 49
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 17 31 25 33
rect 17 29 19 31
rect 21 29 25 31
rect 17 27 25 29
rect 23 25 25 27
rect 31 25 33 37
rect 49 25 51 49
rect 77 49 79 51
rect 81 49 129 51
rect 131 49 193 51
rect 77 47 83 49
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 57 27 63 29
rect 83 31 91 33
rect 83 29 87 31
rect 89 29 91 31
rect 83 27 91 29
rect 57 25 59 27
rect 83 25 85 27
rect 95 25 97 49
rect 127 47 133 49
rect 101 41 107 43
rect 137 41 145 43
rect 179 41 187 43
rect 101 39 103 41
rect 105 39 139 41
rect 141 39 183 41
rect 185 39 187 41
rect 101 37 107 39
rect 137 37 145 39
rect 117 31 123 33
rect 117 29 119 31
rect 121 29 123 31
rect 117 27 123 29
rect 127 31 133 33
rect 127 29 129 31
rect 131 29 133 31
rect 127 27 133 29
rect 119 25 121 27
rect 131 25 133 27
rect 143 25 145 37
rect 179 37 187 39
rect 161 31 169 33
rect 161 29 163 31
rect 165 29 169 31
rect 161 27 169 29
rect 155 21 163 23
rect 155 19 159 21
rect 161 19 163 21
rect 155 17 163 19
rect 155 15 157 17
rect 167 15 169 27
rect 179 25 181 37
rect 191 25 193 49
rect 203 49 207 51
rect 209 49 211 51
rect 203 47 211 49
rect 215 43 217 55
rect 227 43 229 55
rect 205 41 229 43
rect 205 39 207 41
rect 209 39 229 41
rect 205 37 229 39
rect 203 31 211 33
rect 203 29 207 31
rect 209 29 211 31
rect 203 27 211 29
rect 203 25 205 27
rect 215 25 217 37
rect 227 25 229 37
rect 11 12 13 15
rect 23 12 25 15
rect 31 12 33 15
rect 49 12 51 15
rect 57 12 59 15
rect 83 12 85 15
rect 95 12 97 15
rect 119 12 121 15
rect 131 12 133 15
rect 143 12 145 15
rect 179 12 181 15
rect 191 12 193 15
rect 203 12 205 15
rect 155 2 157 5
rect 167 2 169 5
rect 215 2 217 5
rect 227 2 229 5
<< ndif >>
rect 37 31 47 33
rect 37 29 39 31
rect 41 29 47 31
rect 37 25 47 29
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 25 15 31 25
rect 33 15 49 25
rect 51 15 57 25
rect 59 15 67 25
rect 75 21 83 25
rect 75 19 77 21
rect 79 19 83 21
rect 75 15 83 19
rect 85 15 95 25
rect 97 21 105 25
rect 97 19 101 21
rect 103 19 105 21
rect 97 15 105 19
rect 111 15 119 25
rect 121 15 131 25
rect 133 21 143 25
rect 133 19 137 21
rect 139 19 143 21
rect 133 15 143 19
rect 145 15 153 25
rect 171 21 179 25
rect 171 19 173 21
rect 175 19 179 21
rect 171 15 179 19
rect 181 21 191 25
rect 181 19 185 21
rect 187 19 191 21
rect 181 15 191 19
rect 193 15 203 25
rect 205 21 215 25
rect 205 19 209 21
rect 211 19 215 21
rect 205 15 215 19
rect 15 11 21 15
rect 15 9 17 11
rect 19 9 21 11
rect 61 11 67 15
rect 61 9 63 11
rect 65 9 67 11
rect 15 7 21 9
rect 61 7 67 9
rect 87 11 93 15
rect 87 9 89 11
rect 91 9 93 11
rect 87 7 93 9
rect 111 11 117 15
rect 111 9 113 11
rect 115 9 117 11
rect 111 7 117 9
rect 147 5 155 15
rect 157 11 167 15
rect 157 9 161 11
rect 163 9 167 11
rect 157 5 167 9
rect 169 5 177 15
rect 207 11 215 15
rect 207 9 209 11
rect 211 9 215 11
rect 207 5 215 9
rect 217 21 227 25
rect 217 19 221 21
rect 223 19 227 21
rect 217 5 227 19
rect 229 21 237 25
rect 229 19 233 21
rect 235 19 237 21
rect 229 11 237 19
rect 229 9 233 11
rect 235 9 237 11
rect 229 5 237 9
<< pdif >>
rect 15 91 21 93
rect 61 91 67 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 61 89 63 91
rect 65 89 67 91
rect 61 85 67 89
rect 87 91 93 93
rect 87 89 89 91
rect 91 89 93 91
rect 87 85 93 89
rect 111 91 119 95
rect 111 89 113 91
rect 115 89 119 91
rect 3 71 11 85
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 65 23 85
rect 25 65 31 85
rect 33 71 49 85
rect 33 69 39 71
rect 41 69 49 71
rect 33 65 49 69
rect 51 65 57 85
rect 59 65 67 85
rect 75 71 83 85
rect 75 69 77 71
rect 79 69 83 71
rect 75 65 83 69
rect 85 65 95 85
rect 97 71 105 85
rect 111 75 119 89
rect 121 85 129 95
rect 147 85 155 95
rect 121 75 131 85
rect 97 69 101 71
rect 103 69 105 71
rect 97 65 105 69
rect 123 65 131 75
rect 133 71 143 85
rect 133 69 137 71
rect 139 69 143 71
rect 133 65 143 69
rect 145 75 155 85
rect 157 91 167 95
rect 157 89 161 91
rect 163 89 167 91
rect 157 75 167 89
rect 169 81 179 95
rect 169 79 173 81
rect 175 79 179 81
rect 169 75 179 79
rect 181 81 191 95
rect 181 79 185 81
rect 187 79 191 81
rect 181 75 191 79
rect 193 75 203 95
rect 205 91 215 95
rect 205 89 209 91
rect 211 89 215 91
rect 205 81 215 89
rect 205 79 209 81
rect 211 79 215 81
rect 205 75 215 79
rect 145 65 153 75
rect 207 71 215 75
rect 207 69 209 71
rect 211 69 215 71
rect 207 61 215 69
rect 207 59 209 61
rect 211 59 215 61
rect 207 55 215 59
rect 217 81 227 95
rect 217 79 221 81
rect 223 79 227 81
rect 217 71 227 79
rect 217 69 221 71
rect 223 69 227 71
rect 217 61 227 69
rect 217 59 221 61
rect 223 59 227 61
rect 217 55 227 59
rect 229 91 237 95
rect 229 89 233 91
rect 235 89 237 91
rect 229 81 237 89
rect 229 79 233 81
rect 235 79 237 81
rect 229 71 237 79
rect 229 69 233 71
rect 235 69 237 71
rect 229 61 237 69
rect 229 59 233 61
rect 235 59 237 61
rect 229 55 237 59
<< alu1 >>
rect -2 95 242 100
rect -2 93 29 95
rect 31 93 49 95
rect 51 93 242 95
rect -2 91 242 93
rect -2 89 17 91
rect 19 89 63 91
rect 65 89 89 91
rect 91 89 113 91
rect 115 89 161 91
rect 163 89 209 91
rect 211 89 233 91
rect 235 89 242 91
rect -2 88 242 89
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 22 7 68
rect 18 61 22 82
rect 18 59 19 61
rect 21 59 22 61
rect 18 31 22 59
rect 28 51 32 82
rect 172 81 176 82
rect 39 79 121 81
rect 39 72 41 79
rect 119 72 121 79
rect 172 79 173 81
rect 175 79 176 81
rect 172 78 176 79
rect 184 81 188 82
rect 208 81 212 88
rect 184 79 185 81
rect 187 79 199 81
rect 184 78 188 79
rect 38 71 42 72
rect 38 69 39 71
rect 41 69 42 71
rect 38 68 42 69
rect 28 49 29 51
rect 31 49 32 51
rect 28 48 32 49
rect 28 41 32 42
rect 28 39 29 41
rect 31 39 32 41
rect 28 38 32 39
rect 18 29 19 31
rect 21 29 22 31
rect 18 28 22 29
rect 4 21 8 22
rect 29 21 31 38
rect 39 32 41 68
rect 48 61 52 62
rect 48 59 49 61
rect 51 59 52 61
rect 48 58 52 59
rect 58 61 62 72
rect 76 71 80 72
rect 76 69 77 71
rect 79 69 80 71
rect 76 68 80 69
rect 58 59 59 61
rect 61 59 62 61
rect 38 31 42 32
rect 38 29 39 31
rect 41 29 42 31
rect 38 28 42 29
rect 49 21 51 58
rect 4 19 5 21
rect 7 19 51 21
rect 58 31 62 59
rect 58 29 59 31
rect 61 29 62 31
rect 4 18 8 19
rect 58 18 62 29
rect 77 52 79 68
rect 88 62 92 72
rect 100 71 104 72
rect 100 69 101 71
rect 103 69 104 71
rect 100 68 104 69
rect 116 71 121 72
rect 116 69 117 71
rect 119 69 121 71
rect 116 68 121 69
rect 136 71 140 72
rect 158 71 162 72
rect 173 71 175 78
rect 186 71 190 72
rect 136 69 137 71
rect 139 69 151 71
rect 136 68 140 69
rect 86 61 92 62
rect 86 59 87 61
rect 89 59 92 61
rect 86 58 92 59
rect 77 51 82 52
rect 77 49 79 51
rect 81 49 82 51
rect 77 48 82 49
rect 77 22 79 48
rect 88 32 92 58
rect 86 31 92 32
rect 86 29 87 31
rect 89 29 92 31
rect 86 28 92 29
rect 76 21 80 22
rect 76 19 77 21
rect 79 19 80 21
rect 76 18 80 19
rect 88 18 92 28
rect 101 42 103 68
rect 101 41 106 42
rect 101 39 103 41
rect 105 39 106 41
rect 101 38 106 39
rect 101 22 103 38
rect 119 32 121 68
rect 128 61 132 62
rect 149 61 151 69
rect 158 69 159 71
rect 161 69 175 71
rect 158 68 162 69
rect 162 61 166 62
rect 128 59 129 61
rect 131 59 141 61
rect 128 58 132 59
rect 128 51 132 52
rect 128 49 129 51
rect 131 49 132 51
rect 128 48 132 49
rect 129 32 131 48
rect 139 42 141 59
rect 149 59 163 61
rect 165 59 166 61
rect 138 41 142 42
rect 138 39 139 41
rect 141 39 142 41
rect 138 38 142 39
rect 118 31 122 32
rect 118 29 119 31
rect 121 29 122 31
rect 118 28 122 29
rect 128 31 132 32
rect 128 29 129 31
rect 131 29 132 31
rect 128 28 132 29
rect 149 31 151 59
rect 162 58 166 59
rect 162 31 166 32
rect 149 29 163 31
rect 165 29 166 31
rect 100 21 104 22
rect 100 19 101 21
rect 103 19 104 21
rect 100 18 104 19
rect 136 21 140 22
rect 149 21 151 29
rect 162 28 166 29
rect 173 22 175 69
rect 185 69 187 71
rect 189 69 190 71
rect 185 68 190 69
rect 185 42 187 68
rect 182 41 187 42
rect 182 39 183 41
rect 185 39 187 41
rect 197 41 199 79
rect 208 79 209 81
rect 211 79 212 81
rect 208 71 212 79
rect 208 69 209 71
rect 211 69 212 71
rect 208 61 212 69
rect 208 59 209 61
rect 211 59 212 61
rect 208 58 212 59
rect 218 81 224 82
rect 218 79 221 81
rect 223 79 224 81
rect 218 78 224 79
rect 232 81 236 88
rect 232 79 233 81
rect 235 79 236 81
rect 218 72 222 78
rect 218 71 224 72
rect 218 69 221 71
rect 223 69 224 71
rect 218 68 224 69
rect 232 71 236 79
rect 232 69 233 71
rect 235 69 236 71
rect 218 62 222 68
rect 218 61 224 62
rect 218 59 221 61
rect 223 59 224 61
rect 218 58 224 59
rect 232 61 236 69
rect 232 59 233 61
rect 235 59 236 61
rect 232 58 236 59
rect 206 51 210 52
rect 218 51 222 58
rect 206 49 207 51
rect 209 49 223 51
rect 206 48 210 49
rect 206 41 210 42
rect 197 39 207 41
rect 209 39 210 41
rect 182 38 186 39
rect 136 19 137 21
rect 139 19 151 21
rect 158 21 162 22
rect 172 21 176 22
rect 158 19 159 21
rect 161 19 173 21
rect 175 19 176 21
rect 136 18 140 19
rect 158 18 162 19
rect 172 18 176 19
rect 184 21 188 22
rect 197 21 199 39
rect 206 38 210 39
rect 206 31 210 32
rect 218 31 222 49
rect 206 29 207 31
rect 209 29 223 31
rect 206 28 210 29
rect 218 22 222 29
rect 184 19 185 21
rect 187 19 199 21
rect 208 21 212 22
rect 208 19 209 21
rect 211 19 212 21
rect 184 18 188 19
rect 208 12 212 19
rect 218 21 224 22
rect 218 19 221 21
rect 223 19 224 21
rect 218 18 224 19
rect 232 21 236 22
rect 232 19 233 21
rect 235 19 236 21
rect 232 12 236 19
rect -2 11 242 12
rect -2 9 17 11
rect 19 9 63 11
rect 65 9 89 11
rect 91 9 113 11
rect 115 9 161 11
rect 163 9 209 11
rect 211 9 233 11
rect 235 9 242 11
rect -2 7 242 9
rect -2 5 29 7
rect 31 5 49 7
rect 51 5 125 7
rect 127 5 137 7
rect 139 5 185 7
rect 187 5 197 7
rect 199 5 242 7
rect -2 0 242 5
<< ptie >>
rect 27 7 53 9
rect 123 7 141 9
rect 27 5 29 7
rect 31 5 49 7
rect 51 5 53 7
rect 27 3 53 5
rect 123 5 125 7
rect 127 5 137 7
rect 139 5 141 7
rect 183 7 201 9
rect 183 5 185 7
rect 187 5 197 7
rect 199 5 201 7
rect 123 3 141 5
rect 183 3 201 5
<< ntie >>
rect 27 95 53 97
rect 27 93 29 95
rect 31 93 49 95
rect 51 93 53 95
rect 27 91 53 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 31 15 33 25
rect 49 15 51 25
rect 57 15 59 25
rect 83 15 85 25
rect 95 15 97 25
rect 119 15 121 25
rect 131 15 133 25
rect 143 15 145 25
rect 179 15 181 25
rect 191 15 193 25
rect 203 15 205 25
rect 155 5 157 15
rect 167 5 169 15
rect 215 5 217 25
rect 227 5 229 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 31 65 33 85
rect 49 65 51 85
rect 57 65 59 85
rect 83 65 85 85
rect 95 65 97 85
rect 119 75 121 95
rect 131 65 133 85
rect 143 65 145 85
rect 155 75 157 95
rect 167 75 169 95
rect 179 75 181 95
rect 191 75 193 95
rect 203 75 205 95
rect 215 55 217 95
rect 227 55 229 95
<< polyct1 >>
rect 117 69 119 71
rect 159 69 161 71
rect 19 59 21 61
rect 49 59 51 61
rect 59 59 61 61
rect 87 59 89 61
rect 129 59 131 61
rect 163 59 165 61
rect 187 69 189 71
rect 29 49 31 51
rect 29 39 31 41
rect 19 29 21 31
rect 79 49 81 51
rect 129 49 131 51
rect 59 29 61 31
rect 87 29 89 31
rect 103 39 105 41
rect 139 39 141 41
rect 183 39 185 41
rect 119 29 121 31
rect 129 29 131 31
rect 163 29 165 31
rect 159 19 161 21
rect 207 49 209 51
rect 207 39 209 41
rect 207 29 209 31
<< ndifct1 >>
rect 39 29 41 31
rect 5 19 7 21
rect 77 19 79 21
rect 101 19 103 21
rect 137 19 139 21
rect 173 19 175 21
rect 185 19 187 21
rect 209 19 211 21
rect 17 9 19 11
rect 63 9 65 11
rect 89 9 91 11
rect 113 9 115 11
rect 161 9 163 11
rect 209 9 211 11
rect 221 19 223 21
rect 233 19 235 21
rect 233 9 235 11
<< ntiect1 >>
rect 29 93 31 95
rect 49 93 51 95
<< ptiect1 >>
rect 29 5 31 7
rect 49 5 51 7
rect 125 5 127 7
rect 137 5 139 7
rect 185 5 187 7
rect 197 5 199 7
<< pdifct1 >>
rect 17 89 19 91
rect 63 89 65 91
rect 89 89 91 91
rect 113 89 115 91
rect 5 69 7 71
rect 39 69 41 71
rect 77 69 79 71
rect 101 69 103 71
rect 137 69 139 71
rect 161 89 163 91
rect 173 79 175 81
rect 185 79 187 81
rect 209 89 211 91
rect 209 79 211 81
rect 209 69 211 71
rect 209 59 211 61
rect 221 79 223 81
rect 221 69 223 71
rect 221 59 223 61
rect 233 89 235 91
rect 233 79 235 81
rect 233 69 235 71
rect 233 59 235 61
<< labels >>
rlabel alu1 20 55 20 55 6 i0
rlabel alu1 30 65 30 65 6 cmd
rlabel alu1 60 45 60 45 6 i1
rlabel alu1 90 45 90 45 6 ck
rlabel alu1 120 6 120 6 6 vss
rlabel alu1 120 94 120 94 6 vdd
rlabel alu1 220 50 220 50 6 q
<< end >>
