magic
tech scmos
timestamp 1199201950
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 69 41 74
rect 50 69 52 74
rect 60 69 62 74
rect 71 61 73 66
rect 81 61 83 65
rect 50 47 52 52
rect 9 39 11 43
rect 19 39 21 43
rect 29 39 31 47
rect 39 39 41 47
rect 50 45 56 47
rect 50 43 52 45
rect 54 43 56 45
rect 50 41 56 43
rect 60 43 62 52
rect 71 43 73 46
rect 60 41 73 43
rect 81 43 83 46
rect 81 41 87 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 19 33 31 35
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 37 46 39
rect 36 35 42 37
rect 44 35 46 37
rect 36 33 46 35
rect 36 30 38 33
rect 51 29 53 41
rect 64 36 70 41
rect 64 34 66 36
rect 68 34 70 36
rect 81 39 83 41
rect 85 39 87 41
rect 81 37 87 39
rect 81 34 83 37
rect 58 32 70 34
rect 58 29 60 32
rect 68 29 70 32
rect 75 32 83 34
rect 75 29 77 32
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
rect 51 9 53 14
rect 58 9 60 14
rect 68 13 70 18
rect 75 13 77 18
<< ndif >>
rect 3 11 12 30
rect 3 9 6 11
rect 8 10 12 11
rect 14 10 19 30
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 10 29 19
rect 31 10 36 30
rect 38 29 49 30
rect 38 21 51 29
rect 38 19 44 21
rect 46 19 51 21
rect 38 14 51 19
rect 53 14 58 29
rect 60 22 68 29
rect 60 20 63 22
rect 65 20 68 22
rect 60 18 68 20
rect 70 18 75 29
rect 77 22 88 29
rect 77 20 83 22
rect 85 20 88 22
rect 77 18 88 20
rect 60 14 65 18
rect 38 12 44 14
rect 46 12 49 14
rect 38 10 49 12
rect 8 9 10 10
rect 3 7 10 9
<< pdif >>
rect 2 67 9 69
rect 2 65 4 67
rect 6 65 9 67
rect 2 60 9 65
rect 2 58 4 60
rect 6 58 9 60
rect 2 43 9 58
rect 11 61 19 69
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 43 19 52
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 47 29 58
rect 31 61 39 69
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 47 39 52
rect 41 67 50 69
rect 41 65 44 67
rect 46 65 50 67
rect 41 60 50 65
rect 41 58 44 60
rect 46 58 50 60
rect 41 52 50 58
rect 52 56 60 69
rect 52 54 55 56
rect 57 54 60 56
rect 52 52 60 54
rect 62 67 69 69
rect 62 65 65 67
rect 67 65 69 67
rect 62 61 69 65
rect 62 60 71 61
rect 62 58 65 60
rect 67 58 71 60
rect 62 52 71 58
rect 41 47 48 52
rect 21 43 27 47
rect 64 46 71 52
rect 73 59 81 61
rect 73 57 76 59
rect 78 57 81 59
rect 73 52 81 57
rect 73 50 76 52
rect 78 50 81 52
rect 73 46 81 50
rect 83 59 90 61
rect 83 57 86 59
rect 88 57 90 59
rect 83 52 90 57
rect 83 50 86 52
rect 88 50 90 52
rect 83 46 90 50
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 33 61 39 63
rect 33 59 34 61
rect 36 59 39 61
rect 33 54 39 59
rect 2 52 14 54
rect 16 52 34 54
rect 36 52 39 54
rect 2 50 39 52
rect 2 22 6 50
rect 17 42 31 46
rect 25 37 31 42
rect 49 45 87 46
rect 49 43 52 45
rect 54 43 87 45
rect 49 42 87 43
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 81 41 87 42
rect 81 39 83 41
rect 85 39 87 41
rect 65 36 71 38
rect 65 34 66 36
rect 68 34 71 36
rect 81 34 87 39
rect 65 30 71 34
rect 65 26 87 30
rect 2 21 28 22
rect 2 19 24 21
rect 26 19 28 21
rect 2 18 28 19
rect 74 17 78 26
rect -2 11 98 12
rect -2 9 6 11
rect 8 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 51 14 53 29
rect 58 14 60 29
rect 68 18 70 29
rect 75 18 77 29
<< pmos >>
rect 9 43 11 69
rect 19 43 21 69
rect 29 47 31 69
rect 39 47 41 69
rect 50 52 52 69
rect 60 52 62 69
rect 71 46 73 61
rect 81 46 83 61
<< polyct0 >>
rect 11 35 13 37
rect 42 35 44 37
<< polyct1 >>
rect 52 43 54 45
rect 27 35 29 37
rect 66 34 68 36
rect 83 39 85 41
<< ndifct0 >>
rect 44 19 46 21
rect 63 20 65 22
rect 83 20 85 22
rect 44 12 46 14
<< ndifct1 >>
rect 6 9 8 11
rect 24 19 26 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 65 6 67
rect 4 58 6 60
rect 14 59 16 61
rect 24 65 26 67
rect 24 58 26 60
rect 44 65 46 67
rect 44 58 46 60
rect 55 54 57 56
rect 65 65 67 67
rect 65 58 67 60
rect 76 57 78 59
rect 76 50 78 52
rect 86 57 88 59
rect 86 50 88 52
<< pdifct1 >>
rect 14 52 16 54
rect 34 59 36 61
rect 34 52 36 54
<< alu0 >>
rect 2 67 8 68
rect 2 65 4 67
rect 6 65 8 67
rect 2 60 8 65
rect 22 67 28 68
rect 22 65 24 67
rect 26 65 28 67
rect 2 58 4 60
rect 6 58 8 60
rect 2 57 8 58
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 60 28 65
rect 42 67 48 68
rect 42 65 44 67
rect 46 65 48 67
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 42 60 48 65
rect 42 58 44 60
rect 46 58 48 60
rect 63 67 69 68
rect 63 65 65 67
rect 67 65 69 67
rect 63 60 69 65
rect 63 58 65 60
rect 67 58 69 60
rect 42 57 48 58
rect 54 56 58 58
rect 63 57 69 58
rect 75 59 80 61
rect 75 57 76 59
rect 78 57 80 59
rect 54 54 55 56
rect 57 54 58 56
rect 54 53 58 54
rect 75 53 80 57
rect 42 52 80 53
rect 42 50 76 52
rect 78 50 80 52
rect 42 49 80 50
rect 84 59 90 68
rect 84 57 86 59
rect 88 57 90 59
rect 84 52 90 57
rect 84 50 86 52
rect 88 50 90 52
rect 84 49 90 50
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 42 39 46 49
rect 41 37 46 39
rect 41 35 42 37
rect 44 35 46 37
rect 41 30 46 35
rect 10 26 58 30
rect 54 23 58 26
rect 54 22 67 23
rect 42 21 48 22
rect 42 19 44 21
rect 46 19 48 21
rect 54 20 63 22
rect 65 20 67 22
rect 54 19 67 20
rect 42 14 48 19
rect 81 22 87 23
rect 81 20 83 22
rect 85 20 87 22
rect 42 12 44 14
rect 46 12 48 14
rect 81 12 87 20
<< labels >>
rlabel alu0 12 32 12 32 6 an
rlabel alu0 44 39 44 39 6 an
rlabel alu0 60 21 60 21 6 an
rlabel alu0 56 53 56 53 6 an
rlabel alu0 61 51 61 51 6 an
rlabel alu0 77 55 77 55 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 44 20 44 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 36 56 36 56 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 68 32 68 32 6 a2
rlabel alu1 60 44 60 44 6 a1
rlabel alu1 68 44 68 44 6 a1
rlabel alu1 52 44 52 44 6 a1
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 76 24 76 24 6 a2
rlabel alu1 84 28 84 28 6 a2
rlabel polyct1 84 40 84 40 6 a1
rlabel alu1 76 44 76 44 6 a1
<< end >>
