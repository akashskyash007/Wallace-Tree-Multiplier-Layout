magic
tech scmos
timestamp 1199469401
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 13 94 15 98
rect 25 94 27 98
rect 33 94 35 98
rect 45 94 47 98
rect 57 94 59 98
rect 13 52 15 55
rect 25 52 27 55
rect 13 50 27 52
rect 13 48 19 50
rect 21 48 27 50
rect 13 46 27 48
rect 13 35 15 46
rect 25 35 27 46
rect 33 52 35 55
rect 45 52 47 55
rect 57 52 59 55
rect 33 50 41 52
rect 33 48 37 50
rect 39 48 41 50
rect 33 46 41 48
rect 45 50 53 52
rect 45 48 49 50
rect 51 48 53 50
rect 45 46 53 48
rect 57 50 63 52
rect 57 48 59 50
rect 61 48 63 50
rect 57 46 63 48
rect 33 35 35 46
rect 45 35 47 46
rect 57 35 59 46
rect 13 12 15 17
rect 25 12 27 17
rect 33 12 35 17
rect 45 12 47 17
rect 57 12 59 17
<< ndif >>
rect 8 31 13 35
rect 5 29 13 31
rect 5 27 7 29
rect 9 27 13 29
rect 5 21 13 27
rect 5 19 7 21
rect 9 19 13 21
rect 5 17 13 19
rect 15 17 25 35
rect 27 17 33 35
rect 35 31 45 35
rect 35 29 39 31
rect 41 29 45 31
rect 35 17 45 29
rect 47 31 57 35
rect 47 29 51 31
rect 53 29 57 31
rect 47 21 57 29
rect 47 19 51 21
rect 53 19 57 21
rect 47 17 57 19
rect 59 31 67 35
rect 59 29 63 31
rect 65 29 67 31
rect 59 21 67 29
rect 59 19 63 21
rect 65 19 67 21
rect 59 17 67 19
rect 17 11 23 17
rect 17 9 19 11
rect 21 9 23 11
rect 17 7 23 9
<< pdif >>
rect 8 83 13 94
rect 5 81 13 83
rect 5 79 7 81
rect 9 79 13 81
rect 5 73 13 79
rect 5 71 7 73
rect 9 71 13 73
rect 5 69 13 71
rect 8 55 13 69
rect 15 91 25 94
rect 15 89 19 91
rect 21 89 25 91
rect 15 81 25 89
rect 15 79 19 81
rect 21 79 25 81
rect 15 55 25 79
rect 27 55 33 94
rect 35 71 45 94
rect 35 69 39 71
rect 41 69 45 71
rect 35 61 45 69
rect 35 59 39 61
rect 41 59 45 61
rect 35 55 45 59
rect 47 81 57 94
rect 47 79 51 81
rect 53 79 57 81
rect 47 55 57 79
rect 59 91 67 94
rect 59 89 63 91
rect 65 89 67 91
rect 59 81 67 89
rect 59 79 63 81
rect 65 79 67 81
rect 59 55 67 79
<< alu1 >>
rect -2 91 72 100
rect -2 89 19 91
rect 21 89 63 91
rect 65 89 72 91
rect -2 88 72 89
rect 6 81 10 83
rect 6 79 7 81
rect 9 79 10 81
rect 6 73 10 79
rect 18 81 22 88
rect 18 79 19 81
rect 21 79 22 81
rect 18 77 22 79
rect 28 81 55 82
rect 28 79 51 81
rect 53 79 55 81
rect 28 78 55 79
rect 62 81 66 88
rect 62 79 63 81
rect 65 79 66 81
rect 6 71 7 73
rect 9 72 10 73
rect 28 72 32 78
rect 62 77 66 79
rect 9 71 32 72
rect 6 68 32 71
rect 38 71 42 73
rect 38 69 39 71
rect 41 69 42 71
rect 38 63 42 69
rect 8 52 12 63
rect 28 61 42 63
rect 28 59 39 61
rect 41 59 42 61
rect 28 57 42 59
rect 47 68 63 72
rect 8 50 23 52
rect 8 48 19 50
rect 21 48 23 50
rect 8 46 23 48
rect 8 37 12 46
rect 28 32 32 57
rect 36 50 42 53
rect 36 48 37 50
rect 39 48 42 50
rect 36 42 42 48
rect 47 50 53 68
rect 47 48 49 50
rect 51 48 53 50
rect 47 47 53 48
rect 58 50 62 63
rect 58 48 59 50
rect 61 48 62 50
rect 58 42 62 48
rect 36 37 62 42
rect 28 31 43 32
rect 5 29 11 30
rect 5 27 7 29
rect 9 27 11 29
rect 28 29 39 31
rect 41 29 43 31
rect 28 27 43 29
rect 50 31 55 33
rect 50 29 51 31
rect 53 29 55 31
rect 5 22 11 27
rect 50 22 55 29
rect 5 21 55 22
rect 5 19 7 21
rect 9 19 51 21
rect 53 19 55 21
rect 5 18 55 19
rect 62 31 66 33
rect 62 29 63 31
rect 65 29 66 31
rect 62 21 66 29
rect 62 19 63 21
rect 65 19 66 21
rect 62 12 66 19
rect -2 11 72 12
rect -2 9 19 11
rect 21 9 72 11
rect -2 7 72 9
rect -2 5 49 7
rect 51 5 59 7
rect 61 5 72 7
rect -2 0 72 5
<< ptie >>
rect 47 7 63 9
rect 47 5 49 7
rect 51 5 59 7
rect 61 5 63 7
rect 47 3 63 5
<< nmos >>
rect 13 17 15 35
rect 25 17 27 35
rect 33 17 35 35
rect 45 17 47 35
rect 57 17 59 35
<< pmos >>
rect 13 55 15 94
rect 25 55 27 94
rect 33 55 35 94
rect 45 55 47 94
rect 57 55 59 94
<< polyct1 >>
rect 19 48 21 50
rect 37 48 39 50
rect 49 48 51 50
rect 59 48 61 50
<< ndifct1 >>
rect 7 27 9 29
rect 7 19 9 21
rect 39 29 41 31
rect 51 29 53 31
rect 51 19 53 21
rect 63 29 65 31
rect 63 19 65 21
rect 19 9 21 11
<< ptiect1 >>
rect 49 5 51 7
rect 59 5 61 7
<< pdifct1 >>
rect 7 79 9 81
rect 7 71 9 73
rect 19 89 21 91
rect 19 79 21 81
rect 39 69 41 71
rect 39 59 41 61
rect 51 79 53 81
rect 63 89 65 91
rect 63 79 65 81
<< labels >>
rlabel ndifct1 8 20 8 20 6 n4
rlabel ndifct1 8 28 8 28 6 n4
rlabel pdifct1 8 72 8 72 6 n2
rlabel pdifct1 8 80 8 80 6 n2
rlabel ndifct1 52 20 52 20 6 n4
rlabel ndifct1 52 30 52 30 6 n4
rlabel pdifct1 52 80 52 80 6 n2
rlabel alu1 10 50 10 50 6 a
rlabel alu1 30 45 30 45 6 z
rlabel alu1 20 50 20 50 6 a
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 45 40 45 6 b
rlabel alu1 50 40 50 40 6 b
rlabel ndifct1 40 30 40 30 6 z
rlabel alu1 40 65 40 65 6 z
rlabel alu1 50 60 50 60 6 c
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 50 60 50 6 b
rlabel alu1 60 70 60 70 6 c
<< end >>
