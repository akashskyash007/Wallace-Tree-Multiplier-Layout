magic
tech scmos
timestamp 1199542437
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -2 48 62 104
<< pwell >>
rect -2 -4 62 48
<< poly >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 11 43 13 55
rect 23 43 25 55
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 25 43
rect 17 39 19 41
rect 21 39 25 41
rect 17 37 25 39
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 55
rect 35 41 43 43
rect 35 39 39 41
rect 41 39 43 41
rect 35 37 43 39
rect 35 25 37 37
rect 11 2 13 5
rect 23 2 25 5
rect 35 2 37 5
<< ndif >>
rect 15 31 21 33
rect 15 29 17 31
rect 19 29 21 31
rect 15 25 21 29
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 5 11 19
rect 13 5 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 5 35 19
rect 37 11 45 25
rect 37 9 41 11
rect 43 9 45 11
rect 37 5 45 9
<< pdif >>
rect 3 91 11 95
rect 3 89 5 91
rect 7 89 11 91
rect 3 55 11 89
rect 13 55 23 95
rect 25 81 35 95
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 91 45 95
rect 37 89 41 91
rect 43 89 45 91
rect 37 55 45 89
<< alu1 >>
rect -2 95 62 100
rect -2 93 53 95
rect 55 93 62 95
rect -2 91 62 93
rect -2 89 5 91
rect 7 89 41 91
rect 43 89 62 91
rect -2 88 62 89
rect 8 41 12 82
rect 8 39 9 41
rect 11 39 12 41
rect 8 38 12 39
rect 18 41 22 82
rect 18 39 19 41
rect 21 39 22 41
rect 18 38 22 39
rect 28 81 32 82
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 28 32 32 59
rect 16 31 32 32
rect 16 29 17 31
rect 19 29 32 31
rect 16 28 32 29
rect 38 41 42 82
rect 52 59 56 88
rect 52 57 53 59
rect 55 57 56 59
rect 52 56 56 57
rect 38 39 39 41
rect 41 39 42 41
rect 4 21 8 22
rect 28 21 32 22
rect 4 19 5 21
rect 7 19 29 21
rect 31 19 32 21
rect 4 18 8 19
rect 28 18 32 19
rect 38 18 42 39
rect 52 35 56 36
rect 52 33 53 35
rect 55 33 56 35
rect 52 12 56 33
rect -2 11 62 12
rect -2 9 41 11
rect 43 9 62 11
rect -2 7 62 9
rect -2 5 53 7
rect 55 5 62 7
rect -2 0 62 5
<< ptie >>
rect 51 35 57 37
rect 51 33 53 35
rect 55 33 57 35
rect 51 25 57 33
rect 51 7 57 15
rect 51 5 53 7
rect 55 5 57 7
rect 51 3 57 5
<< ntie >>
rect 51 95 57 97
rect 51 93 53 95
rect 55 93 57 95
rect 51 85 57 93
rect 51 59 57 67
rect 51 57 53 59
rect 55 57 57 59
rect 51 55 57 57
<< nmos >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 5 37 25
<< pmos >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 39 39 41 41
<< ndifct1 >>
rect 17 29 19 31
rect 5 19 7 21
rect 29 19 31 21
rect 41 9 43 11
<< ntiect1 >>
rect 53 93 55 95
rect 53 57 55 59
<< ptiect1 >>
rect 53 33 55 35
rect 53 5 55 7
<< pdifct1 >>
rect 5 89 7 91
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
rect 41 89 43 91
<< labels >>
rlabel alu1 10 60 10 60 6 i0
rlabel alu1 20 60 20 60 6 i1
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 40 50 40 50 6 i2
rlabel alu1 30 55 30 55 6 nq
rlabel alu1 30 94 30 94 6 vdd
<< end >>
