magic
tech scmos
timestamp 1199543590
<< ab >>
rect 0 0 160 100
<< nwell >>
rect -2 48 162 104
<< pwell >>
rect -2 -4 162 48
<< poly >>
rect 11 95 13 98
rect 23 95 25 98
rect 47 95 49 98
rect 59 95 61 98
rect 71 95 73 98
rect 83 95 85 98
rect 111 95 113 98
rect 123 95 125 98
rect 135 95 137 98
rect 147 95 149 98
rect 11 53 13 55
rect 7 51 13 53
rect 7 49 9 51
rect 11 49 13 51
rect 7 47 13 49
rect 11 25 13 47
rect 23 53 25 55
rect 47 53 49 55
rect 59 53 61 55
rect 71 53 73 55
rect 83 53 85 55
rect 111 53 113 55
rect 23 51 33 53
rect 23 49 29 51
rect 31 49 33 51
rect 23 47 33 49
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 57 51 63 53
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 67 51 73 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 77 51 85 53
rect 107 51 113 53
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 107 49 109 51
rect 111 49 113 51
rect 107 47 113 49
rect 123 53 125 55
rect 123 51 129 53
rect 123 49 125 51
rect 127 49 129 51
rect 123 47 129 49
rect 23 25 25 47
rect 51 25 53 47
rect 59 25 61 47
rect 71 25 73 47
rect 79 25 81 47
rect 93 41 99 43
rect 135 41 137 55
rect 147 41 149 55
rect 93 39 95 41
rect 97 39 149 41
rect 93 37 99 39
rect 111 31 117 33
rect 111 29 113 31
rect 115 29 117 31
rect 111 27 117 29
rect 115 25 117 27
rect 123 31 129 33
rect 123 29 125 31
rect 127 29 129 31
rect 123 27 129 29
rect 123 25 125 27
rect 135 25 137 39
rect 147 25 149 39
rect 11 2 13 5
rect 23 2 25 5
rect 51 2 53 5
rect 59 2 61 5
rect 71 2 73 5
rect 79 2 81 5
rect 115 2 117 5
rect 123 2 125 5
rect 135 2 137 5
rect 147 2 149 5
<< ndif >>
rect 3 11 11 25
rect 3 9 5 11
rect 7 9 11 11
rect 3 5 11 9
rect 13 5 23 25
rect 25 21 33 25
rect 25 19 29 21
rect 31 19 33 21
rect 25 5 33 19
rect 43 11 51 25
rect 43 9 45 11
rect 47 9 51 11
rect 43 5 51 9
rect 53 5 59 25
rect 61 21 71 25
rect 61 19 65 21
rect 67 19 71 21
rect 61 5 71 19
rect 73 5 79 25
rect 81 11 89 25
rect 107 21 115 25
rect 107 19 109 21
rect 111 19 115 21
rect 81 9 85 11
rect 87 9 89 11
rect 81 5 89 9
rect 107 5 115 19
rect 117 5 123 25
rect 125 11 135 25
rect 125 9 129 11
rect 131 9 135 11
rect 125 5 135 9
rect 137 21 147 25
rect 137 19 141 21
rect 143 19 147 21
rect 137 5 147 19
rect 149 21 157 25
rect 149 19 153 21
rect 155 19 157 21
rect 149 11 157 19
rect 149 9 153 11
rect 155 9 157 11
rect 149 5 157 9
<< pdif >>
rect 3 81 11 95
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 55 11 69
rect 13 71 23 95
rect 13 69 17 71
rect 19 69 23 71
rect 13 55 23 69
rect 25 81 33 95
rect 25 79 29 81
rect 31 79 33 81
rect 25 71 33 79
rect 25 69 29 71
rect 31 69 33 71
rect 25 55 33 69
rect 39 81 47 95
rect 39 79 41 81
rect 43 79 47 81
rect 39 55 47 79
rect 49 71 59 95
rect 49 69 53 71
rect 55 69 59 71
rect 49 55 59 69
rect 61 81 71 95
rect 61 79 65 81
rect 67 79 71 81
rect 61 71 71 79
rect 61 69 65 71
rect 67 69 71 71
rect 61 55 71 69
rect 73 71 83 95
rect 73 69 77 71
rect 79 69 83 71
rect 73 55 83 69
rect 85 81 93 95
rect 85 79 89 81
rect 91 79 93 81
rect 85 55 93 79
rect 103 91 111 95
rect 103 89 105 91
rect 107 89 111 91
rect 103 81 111 89
rect 103 79 105 81
rect 107 79 111 81
rect 103 55 111 79
rect 113 81 123 95
rect 113 79 117 81
rect 119 79 123 81
rect 113 55 123 79
rect 125 91 135 95
rect 125 89 129 91
rect 131 89 135 91
rect 125 81 135 89
rect 125 79 129 81
rect 131 79 135 81
rect 125 55 135 79
rect 137 81 147 95
rect 137 79 141 81
rect 143 79 147 81
rect 137 71 147 79
rect 137 69 141 71
rect 143 69 147 71
rect 137 61 147 69
rect 137 59 141 61
rect 143 59 147 61
rect 137 55 147 59
rect 149 91 157 95
rect 149 89 153 91
rect 155 89 157 91
rect 149 81 157 89
rect 149 79 153 81
rect 155 79 157 81
rect 149 71 157 79
rect 149 69 153 71
rect 155 69 157 71
rect 149 55 157 69
<< alu1 >>
rect -2 91 162 100
rect -2 89 105 91
rect 107 89 129 91
rect 131 89 153 91
rect 155 89 162 91
rect -2 88 162 89
rect 4 81 8 82
rect 28 81 32 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 32 81
rect 4 78 8 79
rect 28 78 32 79
rect 40 81 44 82
rect 64 81 68 82
rect 88 81 92 82
rect 40 79 41 81
rect 43 79 65 81
rect 67 79 89 81
rect 91 79 92 81
rect 40 78 44 79
rect 64 78 68 79
rect 88 78 92 79
rect 104 81 108 88
rect 104 79 105 81
rect 107 79 108 81
rect 104 78 108 79
rect 116 81 120 82
rect 116 79 117 81
rect 119 79 120 81
rect 116 78 120 79
rect 128 81 132 88
rect 128 79 129 81
rect 131 79 132 81
rect 128 78 132 79
rect 138 81 144 82
rect 138 79 141 81
rect 143 79 144 81
rect 138 78 144 79
rect 152 81 156 88
rect 152 79 153 81
rect 155 79 156 81
rect 5 72 7 78
rect 29 72 31 78
rect 65 72 67 78
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 16 71 20 72
rect 28 71 32 72
rect 52 71 56 72
rect 16 69 17 71
rect 19 69 21 71
rect 16 68 21 69
rect 28 69 29 71
rect 31 69 53 71
rect 55 69 56 71
rect 28 68 32 69
rect 52 68 56 69
rect 64 71 68 72
rect 64 69 65 71
rect 67 69 68 71
rect 64 68 68 69
rect 76 71 80 72
rect 117 71 119 78
rect 138 72 142 78
rect 76 69 77 71
rect 79 69 119 71
rect 76 68 80 69
rect 8 51 12 62
rect 8 49 9 51
rect 11 49 12 51
rect 8 18 12 49
rect 19 21 21 68
rect 28 51 32 62
rect 28 49 29 51
rect 31 49 32 51
rect 28 28 32 49
rect 48 51 52 62
rect 48 49 49 51
rect 51 49 52 51
rect 48 28 52 49
rect 58 51 62 62
rect 58 49 59 51
rect 61 49 62 51
rect 58 28 62 49
rect 68 51 72 62
rect 68 49 69 51
rect 71 49 72 51
rect 68 28 72 49
rect 78 51 82 62
rect 78 49 79 51
rect 81 49 82 51
rect 78 28 82 49
rect 108 51 112 62
rect 128 52 132 72
rect 108 49 109 51
rect 111 49 112 51
rect 94 41 98 42
rect 94 39 95 41
rect 97 39 98 41
rect 94 38 98 39
rect 28 21 32 22
rect 64 21 68 22
rect 95 21 97 38
rect 108 32 112 49
rect 124 51 132 52
rect 124 49 125 51
rect 127 49 132 51
rect 124 48 132 49
rect 128 32 132 48
rect 108 31 116 32
rect 108 29 113 31
rect 115 29 116 31
rect 108 28 116 29
rect 124 31 132 32
rect 124 29 125 31
rect 127 29 132 31
rect 124 28 132 29
rect 138 71 144 72
rect 138 69 141 71
rect 143 69 144 71
rect 138 68 144 69
rect 152 71 156 79
rect 152 69 153 71
rect 155 69 156 71
rect 152 68 156 69
rect 138 62 142 68
rect 138 61 144 62
rect 138 59 141 61
rect 143 59 144 61
rect 138 58 144 59
rect 138 22 142 58
rect 108 21 112 22
rect 19 19 29 21
rect 31 19 65 21
rect 67 19 109 21
rect 111 19 112 21
rect 28 18 32 19
rect 64 18 68 19
rect 108 18 112 19
rect 138 21 144 22
rect 138 19 141 21
rect 143 19 144 21
rect 138 18 144 19
rect 152 21 156 22
rect 152 19 153 21
rect 155 19 156 21
rect 152 12 156 19
rect -2 11 162 12
rect -2 9 5 11
rect 7 9 45 11
rect 47 9 85 11
rect 87 9 129 11
rect 131 9 153 11
rect 155 9 162 11
rect -2 7 97 9
rect 99 7 162 9
rect -2 0 162 7
<< ptie >>
rect 95 9 101 17
rect 95 7 97 9
rect 99 7 101 9
rect 95 5 101 7
<< nmos >>
rect 11 5 13 25
rect 23 5 25 25
rect 51 5 53 25
rect 59 5 61 25
rect 71 5 73 25
rect 79 5 81 25
rect 115 5 117 25
rect 123 5 125 25
rect 135 5 137 25
rect 147 5 149 25
<< pmos >>
rect 11 55 13 95
rect 23 55 25 95
rect 47 55 49 95
rect 59 55 61 95
rect 71 55 73 95
rect 83 55 85 95
rect 111 55 113 95
rect 123 55 125 95
rect 135 55 137 95
rect 147 55 149 95
<< polyct1 >>
rect 9 49 11 51
rect 29 49 31 51
rect 49 49 51 51
rect 59 49 61 51
rect 69 49 71 51
rect 79 49 81 51
rect 109 49 111 51
rect 125 49 127 51
rect 95 39 97 41
rect 113 29 115 31
rect 125 29 127 31
<< ndifct1 >>
rect 5 9 7 11
rect 29 19 31 21
rect 45 9 47 11
rect 65 19 67 21
rect 109 19 111 21
rect 85 9 87 11
rect 129 9 131 11
rect 141 19 143 21
rect 153 19 155 21
rect 153 9 155 11
<< ptiect1 >>
rect 97 7 99 9
<< pdifct1 >>
rect 5 79 7 81
rect 5 69 7 71
rect 17 69 19 71
rect 29 79 31 81
rect 29 69 31 71
rect 41 79 43 81
rect 53 69 55 71
rect 65 79 67 81
rect 65 69 67 71
rect 77 69 79 71
rect 89 79 91 81
rect 105 89 107 91
rect 105 79 107 81
rect 117 79 119 81
rect 129 89 131 91
rect 129 79 131 81
rect 141 79 143 81
rect 141 69 143 71
rect 141 59 143 61
rect 153 89 155 91
rect 153 79 155 81
rect 153 69 155 71
<< labels >>
rlabel alu1 10 40 10 40 6 i7
rlabel alu1 50 45 50 45 6 i5
rlabel alu1 30 45 30 45 6 i6
rlabel alu1 80 6 80 6 6 vss
rlabel alu1 80 45 80 45 6 i2
rlabel alu1 70 45 70 45 6 i3
rlabel alu1 60 45 60 45 6 i4
rlabel alu1 80 94 80 94 6 vdd
rlabel alu1 110 45 110 45 6 i1
rlabel alu1 130 50 130 50 6 i0
rlabel alu1 140 50 140 50 6 q
<< end >>
