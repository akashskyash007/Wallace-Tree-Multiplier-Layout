magic
tech scmos
timestamp 1199203371
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< labels >>
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 16 74 16 74 6 vdd
<< end >>
