magic
tech scmos
timestamp 1199203046
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 13 68 15 73
rect 20 68 22 73
rect 27 68 29 73
rect 34 68 36 73
rect 44 61 46 65
rect 51 61 53 65
rect 58 61 60 65
rect 65 61 67 65
rect 13 40 15 43
rect 2 38 15 40
rect 2 36 4 38
rect 6 36 11 38
rect 2 34 11 36
rect 9 22 11 34
rect 20 33 22 43
rect 27 40 29 43
rect 34 40 36 43
rect 44 40 46 43
rect 27 37 30 40
rect 34 38 46 40
rect 17 31 23 33
rect 17 29 19 31
rect 21 29 23 31
rect 17 27 23 29
rect 28 31 30 37
rect 28 29 34 31
rect 28 27 30 29
rect 32 27 34 29
rect 19 22 21 27
rect 28 25 34 27
rect 31 22 33 25
rect 41 22 43 38
rect 51 31 53 43
rect 58 34 60 43
rect 65 40 67 43
rect 65 38 73 40
rect 67 36 69 38
rect 71 36 73 38
rect 67 34 73 36
rect 47 29 53 31
rect 47 27 49 29
rect 51 27 53 29
rect 57 32 63 34
rect 57 30 59 32
rect 61 30 63 32
rect 57 28 63 30
rect 47 25 53 27
rect 57 21 63 23
rect 57 19 59 21
rect 61 19 63 21
rect 57 17 63 19
rect 9 11 11 16
rect 19 11 21 16
rect 31 11 33 16
rect 41 13 43 16
rect 57 13 59 17
rect 41 11 59 13
<< ndif >>
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 20 19 22
rect 11 18 14 20
rect 16 18 19 20
rect 11 16 19 18
rect 21 16 31 22
rect 33 20 41 22
rect 33 18 36 20
rect 38 18 41 20
rect 33 16 41 18
rect 43 20 50 22
rect 43 18 46 20
rect 48 18 50 20
rect 43 16 50 18
rect 23 11 29 16
rect 23 9 25 11
rect 27 9 29 11
rect 23 7 29 9
<< pdif >>
rect 4 71 11 73
rect 4 69 7 71
rect 9 69 11 71
rect 4 68 11 69
rect 4 43 13 68
rect 15 43 20 68
rect 22 43 27 68
rect 29 43 34 68
rect 36 61 41 68
rect 36 53 44 61
rect 36 51 39 53
rect 41 51 44 53
rect 36 43 44 51
rect 46 43 51 61
rect 53 43 58 61
rect 60 43 65 61
rect 67 59 74 61
rect 67 57 70 59
rect 72 57 74 59
rect 67 52 74 57
rect 67 50 70 52
rect 72 50 74 52
rect 67 43 74 50
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 71 82 79
rect -2 69 7 71
rect 9 69 82 71
rect -2 68 82 69
rect 2 58 62 62
rect 2 38 6 58
rect 10 53 43 54
rect 10 51 39 53
rect 41 51 43 53
rect 10 50 43 51
rect 2 36 4 38
rect 2 34 6 36
rect 10 22 14 50
rect 58 46 62 58
rect 18 42 53 46
rect 58 42 73 46
rect 18 31 22 42
rect 49 38 53 42
rect 67 38 73 42
rect 18 29 19 31
rect 21 29 22 31
rect 33 30 39 38
rect 49 34 62 38
rect 67 36 69 38
rect 71 36 73 38
rect 67 35 73 36
rect 58 32 62 34
rect 58 30 59 32
rect 61 30 62 32
rect 18 27 22 29
rect 28 29 53 30
rect 28 27 30 29
rect 32 27 49 29
rect 51 27 53 29
rect 58 28 62 30
rect 28 26 53 27
rect 66 23 70 31
rect 10 20 40 22
rect 10 18 14 20
rect 16 18 36 20
rect 38 18 40 20
rect 10 17 40 18
rect 58 21 70 23
rect 58 19 59 21
rect 61 19 70 21
rect 58 17 70 19
rect -2 11 82 12
rect -2 9 25 11
rect 27 9 82 11
rect -2 1 82 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 9 16 11 22
rect 19 16 21 22
rect 31 16 33 22
rect 41 16 43 22
<< pmos >>
rect 13 43 15 68
rect 20 43 22 68
rect 27 43 29 68
rect 34 43 36 68
rect 44 43 46 61
rect 51 43 53 61
rect 58 43 60 61
rect 65 43 67 61
<< polyct1 >>
rect 4 36 6 38
rect 19 29 21 31
rect 30 27 32 29
rect 69 36 71 38
rect 49 27 51 29
rect 59 30 61 32
rect 59 19 61 21
<< ndifct0 >>
rect 4 18 6 20
rect 46 18 48 20
<< ndifct1 >>
rect 14 18 16 20
rect 36 18 38 20
rect 25 9 27 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 70 57 72 59
rect 70 50 72 52
<< pdifct1 >>
rect 7 69 9 71
rect 39 51 41 53
<< alu0 >>
rect 6 34 7 40
rect 68 59 74 68
rect 68 57 70 59
rect 72 57 74 59
rect 68 52 74 57
rect 68 50 70 52
rect 72 50 74 52
rect 68 49 74 50
rect 3 20 7 22
rect 3 18 4 20
rect 6 18 7 20
rect 3 12 7 18
rect 45 20 49 22
rect 45 18 46 20
rect 48 18 49 20
rect 45 12 49 18
<< labels >>
rlabel alu1 4 48 4 48 6 a
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 32 12 32 6 z
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 36 20 36 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 60 12 60 6 a
rlabel alu1 28 60 28 60 6 a
rlabel alu1 20 60 20 60 6 a
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 44 28 44 28 6 c
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 32 36 32 6 c
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 44 36 44 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 60 44 60 6 a
rlabel alu1 36 60 36 60 6 a
rlabel alu1 40 74 40 74 6 vdd
rlabel polyct1 60 20 60 20 6 d
rlabel alu1 52 36 52 36 6 b
rlabel alu1 60 52 60 52 6 a
rlabel alu1 52 60 52 60 6 a
rlabel alu1 68 24 68 24 6 d
rlabel alu1 68 44 68 44 6 a
<< end >>
