magic
tech scmos
timestamp 1199470274
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -5 48 105 105
<< pwell >>
rect -5 -5 105 48
<< poly >>
rect 15 93 17 98
rect 23 93 25 98
rect 35 93 37 98
rect 43 93 45 98
rect 55 93 57 98
rect 63 93 65 98
rect 75 93 77 98
rect 83 93 85 98
rect 15 47 17 56
rect 23 53 25 56
rect 35 53 37 56
rect 43 53 45 56
rect 55 53 57 56
rect 63 53 65 56
rect 75 53 77 56
rect 23 51 37 53
rect 41 51 47 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 41 49 43 51
rect 45 49 47 51
rect 41 47 47 49
rect 53 51 59 53
rect 63 51 77 53
rect 83 53 85 56
rect 83 51 93 53
rect 53 49 55 51
rect 57 49 59 51
rect 53 47 59 49
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 87 49 89 51
rect 91 49 93 51
rect 87 47 93 49
rect 15 45 23 47
rect 15 44 19 45
rect 17 43 19 44
rect 21 43 23 45
rect 17 41 23 43
rect 31 39 33 47
rect 43 39 45 47
rect 55 39 57 47
rect 67 39 69 47
rect 31 2 33 6
rect 43 2 45 6
rect 55 2 57 6
rect 67 2 69 6
<< ndif >>
rect 26 23 31 39
rect 23 21 31 23
rect 23 19 25 21
rect 27 19 31 21
rect 23 17 31 19
rect 26 6 31 17
rect 33 31 43 39
rect 33 29 37 31
rect 39 29 43 31
rect 33 6 43 29
rect 45 21 55 39
rect 45 19 49 21
rect 51 19 55 21
rect 45 6 55 19
rect 57 11 67 39
rect 57 9 61 11
rect 63 9 67 11
rect 57 6 67 9
rect 69 33 74 39
rect 69 31 77 33
rect 69 29 73 31
rect 75 29 77 31
rect 69 23 77 29
rect 69 21 73 23
rect 75 21 77 23
rect 69 19 77 21
rect 69 6 74 19
<< pdif >>
rect 6 91 15 93
rect 6 89 9 91
rect 11 89 15 91
rect 6 81 15 89
rect 6 79 9 81
rect 11 79 15 81
rect 6 56 15 79
rect 17 56 23 93
rect 25 81 35 93
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 56 35 69
rect 37 56 43 93
rect 45 91 55 93
rect 45 89 49 91
rect 51 89 55 91
rect 45 81 55 89
rect 45 79 49 81
rect 51 79 55 81
rect 45 56 55 79
rect 57 56 63 93
rect 65 71 75 93
rect 65 69 69 71
rect 71 69 75 71
rect 65 61 75 69
rect 65 59 69 61
rect 71 59 75 61
rect 65 56 75 59
rect 77 56 83 93
rect 85 91 94 93
rect 85 89 89 91
rect 91 89 94 91
rect 85 81 94 89
rect 85 79 89 81
rect 91 79 94 81
rect 85 71 94 79
rect 85 69 89 71
rect 91 69 94 71
rect 85 56 94 69
<< alu1 >>
rect -2 91 102 100
rect -2 89 9 91
rect 11 89 49 91
rect 51 89 89 91
rect 91 89 102 91
rect -2 88 102 89
rect 8 81 12 88
rect 8 79 9 81
rect 11 79 12 81
rect 8 77 12 79
rect 28 81 32 83
rect 28 79 29 81
rect 31 79 32 81
rect 28 72 32 79
rect 48 81 52 88
rect 48 79 49 81
rect 51 79 52 81
rect 48 77 52 79
rect 88 81 92 88
rect 88 79 89 81
rect 91 79 92 81
rect 7 71 73 72
rect 7 69 29 71
rect 31 69 69 71
rect 71 69 73 71
rect 7 68 73 69
rect 7 32 12 68
rect 18 58 42 63
rect 67 61 73 68
rect 67 59 69 61
rect 71 59 73 61
rect 67 58 73 59
rect 18 45 22 58
rect 38 53 42 58
rect 78 53 82 73
rect 88 71 92 79
rect 88 69 89 71
rect 91 69 92 71
rect 88 67 92 69
rect 18 43 19 45
rect 21 43 22 45
rect 18 37 22 43
rect 27 51 33 52
rect 27 49 29 51
rect 31 49 33 51
rect 27 42 33 49
rect 38 51 47 53
rect 38 49 43 51
rect 45 49 47 51
rect 38 47 47 49
rect 53 51 63 53
rect 53 49 55 51
rect 57 49 63 51
rect 53 47 63 49
rect 68 51 82 53
rect 68 49 69 51
rect 71 49 82 51
rect 68 47 82 49
rect 87 51 93 62
rect 87 49 89 51
rect 91 49 93 51
rect 57 42 63 47
rect 87 42 93 49
rect 27 38 53 42
rect 57 38 93 42
rect 7 31 43 32
rect 7 29 37 31
rect 39 29 43 31
rect 7 28 43 29
rect 47 28 53 38
rect 72 31 76 33
rect 72 29 73 31
rect 75 29 76 31
rect 72 23 76 29
rect 72 22 73 23
rect 23 21 73 22
rect 75 21 76 23
rect 23 19 25 21
rect 27 19 49 21
rect 51 19 76 21
rect 23 18 76 19
rect -2 11 102 12
rect -2 9 61 11
rect 63 9 102 11
rect -2 7 102 9
rect -2 5 83 7
rect 85 5 93 7
rect 95 5 102 7
rect -2 0 102 5
<< ptie >>
rect 81 7 97 9
rect 81 5 83 7
rect 85 5 93 7
rect 95 5 97 7
rect 81 3 97 5
<< nmos >>
rect 31 6 33 39
rect 43 6 45 39
rect 55 6 57 39
rect 67 6 69 39
<< pmos >>
rect 15 56 17 93
rect 23 56 25 93
rect 35 56 37 93
rect 43 56 45 93
rect 55 56 57 93
rect 63 56 65 93
rect 75 56 77 93
rect 83 56 85 93
<< polyct1 >>
rect 29 49 31 51
rect 43 49 45 51
rect 55 49 57 51
rect 69 49 71 51
rect 89 49 91 51
rect 19 43 21 45
<< ndifct1 >>
rect 25 19 27 21
rect 37 29 39 31
rect 49 19 51 21
rect 61 9 63 11
rect 73 29 75 31
rect 73 21 75 23
<< ptiect1 >>
rect 83 5 85 7
rect 93 5 95 7
<< pdifct1 >>
rect 9 89 11 91
rect 9 79 11 81
rect 29 79 31 81
rect 29 69 31 71
rect 49 89 51 91
rect 49 79 51 81
rect 69 69 71 71
rect 69 59 71 61
rect 89 89 91 91
rect 89 79 91 81
rect 89 69 91 71
<< labels >>
rlabel ndifct1 26 20 26 20 6 n3
rlabel ndifct1 50 20 50 20 6 n3
rlabel ndifct1 74 22 74 22 6 n3
rlabel ndifct1 74 30 74 30 6 n3
rlabel alu1 10 50 10 50 6 z
rlabel alu1 20 30 20 30 6 z
rlabel alu1 30 30 30 30 6 z
rlabel alu1 20 50 20 50 6 b1
rlabel alu1 30 45 30 45 6 b2
rlabel alu1 30 60 30 60 6 b1
rlabel alu1 20 70 20 70 6 z
rlabel alu1 30 75 30 75 6 z
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 40 30 40 30 6 z
rlabel alu1 50 35 50 35 6 b2
rlabel alu1 40 40 40 40 6 b2
rlabel alu1 40 55 40 55 6 b1
rlabel alu1 40 70 40 70 6 z
rlabel alu1 50 70 50 70 6 z
rlabel alu1 50 94 50 94 6 vdd
rlabel alu1 70 40 70 40 6 a1
rlabel alu1 60 45 60 45 6 a1
rlabel polyct1 70 50 70 50 6 a2
rlabel alu1 60 70 60 70 6 z
rlabel alu1 70 65 70 65 6 z
rlabel alu1 80 40 80 40 6 a1
rlabel polyct1 90 50 90 50 6 a1
rlabel alu1 80 60 80 60 6 a2
<< end >>
