magic
tech scmos
timestamp 1199469133
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 11 93 13 98
rect 33 93 35 98
rect 45 93 47 98
rect 57 93 59 98
rect 11 52 13 55
rect 33 52 35 55
rect 45 52 47 55
rect 57 52 59 55
rect 11 50 22 52
rect 15 48 18 50
rect 20 48 22 50
rect 15 46 22 48
rect 33 50 41 52
rect 33 48 37 50
rect 39 48 41 50
rect 33 46 41 48
rect 45 50 53 52
rect 45 48 49 50
rect 51 48 53 50
rect 45 46 53 48
rect 57 50 63 52
rect 57 48 59 50
rect 61 48 63 50
rect 57 46 63 48
rect 15 35 17 46
rect 33 35 35 46
rect 45 35 47 46
rect 57 40 59 46
rect 53 38 59 40
rect 53 35 55 38
rect 33 20 35 25
rect 15 11 17 16
rect 45 13 47 18
rect 53 13 55 18
<< ndif >>
rect 7 33 15 35
rect 7 31 9 33
rect 11 31 15 33
rect 7 25 15 31
rect 7 23 9 25
rect 11 23 15 25
rect 7 21 15 23
rect 10 16 15 21
rect 17 31 33 35
rect 17 29 21 31
rect 23 29 33 31
rect 17 25 33 29
rect 35 33 45 35
rect 35 31 39 33
rect 41 31 45 33
rect 35 25 45 31
rect 17 21 31 25
rect 17 19 21 21
rect 23 19 31 21
rect 17 16 31 19
rect 40 18 45 25
rect 47 18 53 35
rect 55 31 64 35
rect 55 29 59 31
rect 61 29 64 31
rect 55 22 64 29
rect 55 20 59 22
rect 61 20 64 22
rect 55 18 64 20
<< pdif >>
rect 6 73 11 93
rect 3 71 11 73
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 57 11 59
rect 6 55 11 57
rect 13 91 21 93
rect 13 89 17 91
rect 19 89 21 91
rect 13 81 21 89
rect 13 79 17 81
rect 19 79 21 81
rect 13 75 21 79
rect 13 55 19 75
rect 28 69 33 93
rect 25 67 33 69
rect 25 65 27 67
rect 29 65 33 67
rect 25 59 33 65
rect 25 57 27 59
rect 29 57 33 59
rect 25 55 33 57
rect 35 81 45 93
rect 35 79 39 81
rect 41 79 45 81
rect 35 55 45 79
rect 47 91 57 93
rect 47 89 51 91
rect 53 89 57 91
rect 47 55 57 89
rect 59 83 64 93
rect 59 81 67 83
rect 59 79 63 81
rect 65 79 67 81
rect 59 77 67 79
rect 59 55 64 77
<< alu1 >>
rect -2 91 72 100
rect -2 89 17 91
rect 19 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 16 81 20 88
rect 16 79 17 81
rect 19 79 20 81
rect 16 77 20 79
rect 37 81 67 82
rect 37 79 39 81
rect 41 79 63 81
rect 65 79 67 81
rect 37 78 67 79
rect 4 71 22 73
rect 4 69 5 71
rect 7 69 22 71
rect 4 67 22 69
rect 26 67 30 69
rect 8 63 12 67
rect 4 61 12 63
rect 4 59 5 61
rect 7 59 12 61
rect 4 57 12 59
rect 8 33 12 57
rect 26 65 27 67
rect 29 65 30 67
rect 26 59 30 65
rect 26 57 27 59
rect 29 57 30 59
rect 26 51 30 57
rect 38 68 53 73
rect 38 52 42 68
rect 58 63 62 73
rect 16 50 30 51
rect 16 48 18 50
rect 20 48 30 50
rect 16 47 30 48
rect 26 42 30 47
rect 36 50 42 52
rect 36 48 37 50
rect 39 48 42 50
rect 36 46 42 48
rect 48 57 62 63
rect 48 50 52 57
rect 48 48 49 50
rect 51 48 52 50
rect 48 46 52 48
rect 57 50 63 52
rect 57 48 59 50
rect 61 48 63 50
rect 57 42 63 48
rect 26 38 42 42
rect 38 33 42 38
rect 8 31 9 33
rect 11 31 12 33
rect 8 25 12 31
rect 8 23 9 25
rect 11 23 12 25
rect 8 17 12 23
rect 20 31 24 33
rect 20 29 21 31
rect 23 29 24 31
rect 38 31 39 33
rect 41 31 42 33
rect 38 29 42 31
rect 47 38 63 42
rect 20 21 24 29
rect 20 19 21 21
rect 23 19 24 21
rect 20 12 24 19
rect 47 18 53 38
rect 58 31 62 33
rect 58 29 59 31
rect 61 29 62 31
rect 58 22 62 29
rect 58 20 59 22
rect 61 20 62 22
rect 58 12 62 20
rect -2 7 72 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 72 7
rect -2 0 72 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< nmos >>
rect 15 16 17 35
rect 33 25 35 35
rect 45 18 47 35
rect 53 18 55 35
<< pmos >>
rect 11 55 13 93
rect 33 55 35 93
rect 45 55 47 93
rect 57 55 59 93
<< polyct1 >>
rect 18 48 20 50
rect 37 48 39 50
rect 49 48 51 50
rect 59 48 61 50
<< ndifct1 >>
rect 9 31 11 33
rect 9 23 11 25
rect 21 29 23 31
rect 39 31 41 33
rect 21 19 23 21
rect 59 29 61 31
rect 59 20 61 22
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 5 69 7 71
rect 5 59 7 61
rect 17 89 19 91
rect 17 79 19 81
rect 27 65 29 67
rect 27 57 29 59
rect 39 79 41 81
rect 51 89 53 91
rect 63 79 65 81
<< labels >>
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 70 20 70 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 23 49 23 49 6 zn
rlabel alu1 28 53 28 53 6 zn
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 50 30 50 30 6 a1
rlabel alu1 40 35 40 35 6 zn
rlabel alu1 50 55 50 55 6 a2
rlabel alu1 40 60 40 60 6 b
rlabel alu1 50 70 50 70 6 b
rlabel alu1 60 45 60 45 6 a1
rlabel alu1 60 65 60 65 6 a2
rlabel alu1 52 80 52 80 6 n2
<< end >>
