magic
tech scmos
timestamp 1199541682
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -5 48 55 105
<< pwell >>
rect -5 -5 55 48
<< poly >>
rect 17 94 19 98
rect 25 94 27 98
rect 37 76 39 80
rect 17 43 19 55
rect 13 41 21 43
rect 13 39 17 41
rect 19 39 21 41
rect 13 37 21 39
rect 25 41 27 55
rect 37 53 39 56
rect 31 51 39 53
rect 31 49 33 51
rect 35 49 39 51
rect 31 47 39 49
rect 41 41 47 43
rect 25 39 43 41
rect 45 39 47 41
rect 13 25 15 37
rect 25 25 27 39
rect 41 37 47 39
rect 31 31 39 33
rect 31 29 33 31
rect 35 29 39 31
rect 31 27 39 29
rect 37 24 39 27
rect 13 11 15 15
rect 25 11 27 15
rect 37 10 39 14
<< ndif >>
rect 5 15 13 25
rect 15 21 25 25
rect 15 19 19 21
rect 21 19 25 21
rect 15 15 25 19
rect 27 24 32 25
rect 27 15 37 24
rect 5 11 11 15
rect 29 14 37 15
rect 39 21 47 24
rect 39 19 43 21
rect 45 19 47 21
rect 39 14 47 19
rect 29 11 35 14
rect 5 9 7 11
rect 9 9 11 11
rect 5 7 11 9
rect 29 9 31 11
rect 33 9 35 11
rect 29 7 35 9
<< pdif >>
rect 12 85 17 94
rect 5 81 17 85
rect 5 79 7 81
rect 9 79 17 81
rect 5 71 17 79
rect 5 69 7 71
rect 9 69 17 71
rect 5 61 17 69
rect 5 59 7 61
rect 9 59 17 61
rect 5 55 17 59
rect 19 55 25 94
rect 27 91 35 94
rect 27 89 31 91
rect 33 89 35 91
rect 27 76 35 89
rect 27 56 37 76
rect 39 71 47 76
rect 39 69 43 71
rect 45 69 47 71
rect 39 61 47 69
rect 39 59 43 61
rect 45 59 47 61
rect 39 56 47 59
rect 27 55 32 56
<< alu1 >>
rect -2 95 52 100
rect -2 93 43 95
rect 45 93 52 95
rect -2 91 52 93
rect -2 89 31 91
rect 33 89 52 91
rect -2 88 52 89
rect 8 82 12 83
rect 5 81 12 82
rect 5 79 7 81
rect 9 79 12 81
rect 5 78 12 79
rect 8 72 12 78
rect 5 71 12 72
rect 5 69 7 71
rect 9 69 12 71
rect 5 68 12 69
rect 8 62 12 68
rect 5 61 12 62
rect 5 59 7 61
rect 9 59 12 61
rect 5 58 12 59
rect 8 52 12 58
rect 4 47 12 52
rect 4 33 8 47
rect 18 42 22 83
rect 15 41 22 42
rect 15 39 17 41
rect 19 39 22 41
rect 15 38 22 39
rect 4 28 12 33
rect 8 22 12 28
rect 18 27 22 38
rect 28 52 32 83
rect 42 71 46 73
rect 42 69 43 71
rect 45 69 46 71
rect 42 61 46 69
rect 42 59 43 61
rect 45 59 46 61
rect 28 51 37 52
rect 28 49 33 51
rect 35 49 37 51
rect 28 48 37 49
rect 28 32 32 48
rect 42 41 46 59
rect 42 39 43 41
rect 45 39 46 41
rect 28 31 37 32
rect 28 29 33 31
rect 35 29 37 31
rect 28 28 37 29
rect 8 21 23 22
rect 8 19 19 21
rect 21 19 23 21
rect 8 18 23 19
rect 8 17 12 18
rect 28 17 32 28
rect 42 21 46 39
rect 42 19 43 21
rect 45 19 46 21
rect 42 17 46 19
rect -2 11 52 12
rect -2 9 7 11
rect 9 9 31 11
rect 33 9 52 11
rect -2 0 52 9
<< ntie >>
rect 41 95 47 97
rect 41 93 43 95
rect 45 93 47 95
rect 41 86 47 93
<< nmos >>
rect 13 15 15 25
rect 25 15 27 25
rect 37 14 39 24
<< pmos >>
rect 17 55 19 94
rect 25 55 27 94
rect 37 56 39 76
<< polyct1 >>
rect 17 39 19 41
rect 33 49 35 51
rect 43 39 45 41
rect 33 29 35 31
<< ndifct1 >>
rect 19 19 21 21
rect 43 19 45 21
rect 7 9 9 11
rect 31 9 33 11
<< ntiect1 >>
rect 43 93 45 95
<< pdifct1 >>
rect 7 79 9 81
rect 7 69 9 71
rect 7 59 9 61
rect 31 89 33 91
rect 43 69 45 71
rect 43 59 45 61
<< labels >>
rlabel ndifct1 20 20 20 20 6 q
rlabel alu1 10 25 10 25 6 q
rlabel alu1 10 65 10 65 6 q
rlabel alu1 20 55 20 55 6 i0
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 50 30 50 6 i1
rlabel alu1 25 94 25 94 6 vdd
<< end >>
