magic
tech scmos
timestamp 1199541576
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -2 48 62 104
<< pwell >>
rect -2 -4 62 48
<< poly >>
rect 47 95 49 98
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 11 43 13 65
rect 23 63 25 65
rect 19 61 25 63
rect 19 53 21 61
rect 35 53 37 65
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 27 51 37 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 11 35 13 37
rect 19 35 21 47
rect 27 35 29 47
rect 47 43 49 55
rect 37 41 49 43
rect 37 39 39 41
rect 41 39 49 41
rect 37 37 49 39
rect 47 25 49 37
rect 11 12 13 15
rect 19 12 21 15
rect 27 12 29 15
rect 47 2 49 5
<< ndif >>
rect 3 21 11 35
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 19 35
rect 21 15 27 35
rect 29 25 37 35
rect 29 15 47 25
rect 31 11 47 15
rect 31 9 33 11
rect 35 9 41 11
rect 43 9 47 11
rect 31 5 47 9
rect 49 21 57 25
rect 49 19 53 21
rect 55 19 57 21
rect 49 5 57 19
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 39 91 47 95
rect 39 89 41 91
rect 43 89 47 91
rect 39 85 47 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 65 11 79
rect 13 65 23 85
rect 25 81 35 85
rect 25 79 29 81
rect 31 79 35 81
rect 25 65 35 79
rect 37 65 47 85
rect 39 55 47 65
rect 49 81 57 95
rect 49 79 53 81
rect 55 79 57 81
rect 49 71 57 79
rect 49 69 53 71
rect 55 69 57 71
rect 49 61 57 69
rect 49 59 53 61
rect 55 59 57 61
rect 49 55 57 59
<< alu1 >>
rect -2 91 62 100
rect -2 89 17 91
rect 19 89 41 91
rect 43 89 62 91
rect -2 88 62 89
rect 4 81 8 82
rect 28 81 32 82
rect 48 81 56 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 41 81
rect 4 78 8 79
rect 28 78 32 79
rect 8 41 12 72
rect 8 39 9 41
rect 11 39 12 41
rect 8 28 12 39
rect 18 51 22 72
rect 18 49 19 51
rect 21 49 22 51
rect 18 28 22 49
rect 28 51 32 72
rect 28 49 29 51
rect 31 49 32 51
rect 28 28 32 49
rect 39 42 41 79
rect 48 79 53 81
rect 55 79 56 81
rect 48 78 56 79
rect 48 72 52 78
rect 48 71 56 72
rect 48 69 53 71
rect 55 69 56 71
rect 48 68 56 69
rect 48 62 52 68
rect 48 61 56 62
rect 48 59 53 61
rect 55 59 56 61
rect 48 58 56 59
rect 38 41 42 42
rect 38 39 39 41
rect 41 39 42 41
rect 38 38 42 39
rect 4 21 8 22
rect 39 21 41 38
rect 4 19 5 21
rect 7 19 41 21
rect 48 22 52 58
rect 48 21 56 22
rect 48 19 53 21
rect 55 19 56 21
rect 4 18 8 19
rect 48 18 56 19
rect -2 11 62 12
rect -2 9 33 11
rect 35 9 41 11
rect 43 9 62 11
rect -2 7 62 9
rect -2 5 5 7
rect 7 5 13 7
rect 15 5 21 7
rect 23 5 62 7
rect -2 0 62 5
<< ptie >>
rect 3 7 25 9
rect 3 5 5 7
rect 7 5 13 7
rect 15 5 21 7
rect 23 5 25 7
rect 3 3 25 5
<< nmos >>
rect 11 15 13 35
rect 19 15 21 35
rect 27 15 29 35
rect 47 5 49 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 55 49 95
<< polyct1 >>
rect 19 49 21 51
rect 29 49 31 51
rect 9 39 11 41
rect 39 39 41 41
<< ndifct1 >>
rect 5 19 7 21
rect 33 9 35 11
rect 41 9 43 11
rect 53 19 55 21
<< ptiect1 >>
rect 5 5 7 7
rect 13 5 15 7
rect 21 5 23 7
<< pdifct1 >>
rect 17 89 19 91
rect 41 89 43 91
rect 5 79 7 81
rect 29 79 31 81
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
<< labels >>
rlabel alu1 10 50 10 50 6 i0
rlabel polyct1 20 50 20 50 6 i1
rlabel alu1 30 6 30 6 6 vss
rlabel polyct1 30 50 30 50 6 i2
rlabel alu1 30 94 30 94 6 vdd
rlabel alu1 50 50 50 50 6 q
<< end >>
