magic
tech scmos
timestamp 1199203155
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 13 70 15 74
rect 21 70 23 74
rect 31 70 33 74
rect 39 70 41 74
rect 13 40 15 43
rect 21 40 23 43
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 19 38 25 40
rect 31 39 33 43
rect 39 40 41 43
rect 19 36 21 38
rect 23 36 25 38
rect 19 34 25 36
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 9 30 11 34
rect 19 30 21 34
rect 29 33 35 35
rect 39 38 48 40
rect 39 36 44 38
rect 46 36 48 38
rect 39 34 48 36
rect 29 27 31 33
rect 41 27 43 34
rect 9 11 11 16
rect 19 11 21 16
rect 29 11 31 16
rect 41 11 43 16
<< ndif >>
rect 4 22 9 30
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 16 19 26
rect 21 27 26 30
rect 21 20 29 27
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 31 16 41 27
rect 43 22 48 27
rect 43 20 50 22
rect 43 18 46 20
rect 48 18 50 20
rect 43 16 50 18
rect 33 11 39 16
rect 33 9 35 11
rect 37 9 39 11
rect 33 7 39 9
<< pdif >>
rect 5 68 13 70
rect 5 66 8 68
rect 10 66 13 68
rect 5 43 13 66
rect 15 43 21 70
rect 23 61 31 70
rect 23 59 26 61
rect 28 59 31 61
rect 23 43 31 59
rect 33 43 39 70
rect 41 68 48 70
rect 41 66 44 68
rect 46 66 48 68
rect 41 61 48 66
rect 41 59 44 61
rect 46 59 48 61
rect 41 43 48 59
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 61 30 62
rect 2 59 26 61
rect 28 59 30 61
rect 2 58 30 59
rect 2 29 6 58
rect 34 54 38 63
rect 10 50 23 54
rect 34 50 47 54
rect 10 38 14 50
rect 10 36 11 38
rect 13 36 14 38
rect 10 33 14 36
rect 18 42 39 46
rect 18 38 24 42
rect 43 38 47 50
rect 18 36 21 38
rect 23 36 24 38
rect 18 33 24 36
rect 29 37 39 38
rect 29 35 31 37
rect 33 35 39 37
rect 29 34 39 35
rect 43 36 44 38
rect 46 36 47 38
rect 43 34 47 36
rect 33 30 39 34
rect 2 28 18 29
rect 2 26 14 28
rect 16 26 18 28
rect 33 26 47 30
rect 2 25 18 26
rect -2 11 58 12
rect -2 9 35 11
rect 37 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 27
rect 41 16 43 27
<< pmos >>
rect 13 43 15 70
rect 21 43 23 70
rect 31 43 33 70
rect 39 43 41 70
<< polyct1 >>
rect 11 36 13 38
rect 21 36 23 38
rect 31 35 33 37
rect 44 36 46 38
<< ndifct0 >>
rect 4 18 6 20
rect 24 18 26 20
rect 46 18 48 20
<< ndifct1 >>
rect 14 26 16 28
rect 35 9 37 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 8 66 10 68
rect 44 66 46 68
rect 44 59 46 61
<< pdifct1 >>
rect 26 59 28 61
<< alu0 >>
rect 6 66 8 68
rect 10 66 12 68
rect 6 65 12 66
rect 42 66 44 68
rect 46 66 48 68
rect 42 61 48 66
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 2 20 50 21
rect 2 18 4 20
rect 6 18 24 20
rect 26 18 46 20
rect 48 18 50 20
rect 2 17 50 18
<< labels >>
rlabel alu0 26 19 26 19 6 n3
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 36 20 36 6 b2
rlabel alu1 12 40 12 40 6 b1
rlabel alu1 20 52 20 52 6 b1
rlabel alu1 20 60 20 60 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 32 36 32 6 a2
rlabel alu1 36 44 36 44 6 b2
rlabel alu1 28 44 28 44 6 b2
rlabel alu1 36 60 36 60 6 a1
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 44 52 44 52 6 a1
<< end >>
