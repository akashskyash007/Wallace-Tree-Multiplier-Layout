magic
tech scmos
timestamp 1199202370
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 61 61 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 37 42 39
rect 20 30 22 37
rect 29 35 37 37
rect 39 35 42 37
rect 29 33 42 35
rect 49 37 61 39
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 30 30 32 33
rect 40 30 42 33
rect 50 30 52 33
rect 20 10 22 15
rect 30 10 32 15
rect 40 9 42 14
rect 50 9 52 14
<< ndif >>
rect 13 27 20 30
rect 13 25 15 27
rect 17 25 20 27
rect 13 19 20 25
rect 13 17 15 19
rect 17 17 20 19
rect 13 15 20 17
rect 22 28 30 30
rect 22 26 25 28
rect 27 26 30 28
rect 22 21 30 26
rect 22 19 25 21
rect 27 19 30 21
rect 22 15 30 19
rect 32 19 40 30
rect 32 17 35 19
rect 37 17 40 19
rect 32 15 40 17
rect 34 14 40 15
rect 42 28 50 30
rect 42 26 45 28
rect 47 26 50 28
rect 42 21 50 26
rect 42 19 45 21
rect 47 19 50 21
rect 42 14 50 19
rect 52 18 59 30
rect 52 16 55 18
rect 57 16 59 18
rect 52 14 59 16
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 42 9 52
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 60 29 66
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 53 39 70
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 60 49 66
rect 41 58 44 60
rect 46 58 49 60
rect 41 42 49 58
rect 51 61 56 70
rect 51 53 59 61
rect 51 51 54 53
rect 56 51 59 53
rect 51 46 59 51
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 59 68 61
rect 61 57 64 59
rect 66 57 68 59
rect 61 52 68 57
rect 61 50 64 52
rect 66 50 68 52
rect 61 42 68 50
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 33 53 38 55
rect 33 51 34 53
rect 36 51 38 53
rect 33 46 38 51
rect 9 44 14 46
rect 16 44 34 46
rect 36 44 54 46
rect 56 44 63 46
rect 9 42 63 44
rect 26 30 30 42
rect 35 37 63 38
rect 35 35 37 37
rect 39 35 51 37
rect 53 35 63 37
rect 35 34 63 35
rect 23 28 47 30
rect 23 26 25 28
rect 27 26 45 28
rect 23 21 27 26
rect 23 19 25 21
rect 23 17 27 19
rect 42 21 47 26
rect 42 19 45 21
rect 42 17 47 19
rect 58 25 63 34
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 20 15 22 30
rect 30 15 32 30
rect 40 14 42 30
rect 50 14 52 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 61
<< polyct1 >>
rect 37 35 39 37
rect 51 35 53 37
<< ndifct0 >>
rect 15 25 17 27
rect 15 17 17 19
rect 35 17 37 19
rect 55 16 57 18
<< ndifct1 >>
rect 25 26 27 28
rect 25 19 27 21
rect 45 26 47 28
rect 45 19 47 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 4 52 6 54
rect 14 51 16 53
rect 24 66 26 68
rect 24 58 26 60
rect 44 66 46 68
rect 44 58 46 60
rect 54 51 56 53
rect 64 57 66 59
rect 64 50 66 52
<< pdifct1 >>
rect 14 44 16 46
rect 34 51 36 53
rect 34 44 36 46
rect 54 44 56 46
<< alu0 >>
rect 3 66 4 68
rect 6 66 7 68
rect 3 61 7 66
rect 3 59 4 61
rect 6 59 7 61
rect 3 54 7 59
rect 23 66 24 68
rect 26 66 27 68
rect 23 60 27 66
rect 23 58 24 60
rect 26 58 27 60
rect 23 56 27 58
rect 43 66 44 68
rect 46 66 47 68
rect 43 60 47 66
rect 43 58 44 60
rect 46 58 47 60
rect 43 56 47 58
rect 62 59 68 68
rect 62 57 64 59
rect 66 57 68 59
rect 3 52 4 54
rect 6 52 7 54
rect 3 50 7 52
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 13 46 17 51
rect 53 53 57 55
rect 53 51 54 53
rect 56 51 57 53
rect 53 46 57 51
rect 62 52 68 57
rect 62 50 64 52
rect 66 50 68 52
rect 62 49 68 50
rect 14 27 18 29
rect 14 25 15 27
rect 17 25 18 27
rect 14 19 18 25
rect 14 17 15 19
rect 17 17 18 19
rect 27 17 28 26
rect 34 19 38 21
rect 34 17 35 19
rect 37 17 38 19
rect 47 17 48 30
rect 54 18 58 20
rect 14 12 18 17
rect 34 12 38 17
rect 54 16 55 18
rect 57 16 58 18
rect 54 12 58 16
<< labels >>
rlabel alu1 12 44 12 44 6 z
rlabel alu1 28 36 28 36 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 28 36 28 6 z
rlabel alu1 44 36 44 36 6 a
rlabel polyct1 52 36 52 36 6 a
rlabel alu1 44 24 44 24 6 z
rlabel alu1 44 44 44 44 6 z
rlabel alu1 52 44 52 44 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 32 60 32 6 a
rlabel alu1 60 44 60 44 6 z
<< end >>
