magic
tech scmos
timestamp 1199202918
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 37 28 39
rect 22 35 24 37
rect 26 35 28 37
rect 22 33 28 35
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 33 37 45 39
rect 49 37 55 39
rect 33 35 35 37
rect 37 35 39 37
rect 33 33 39 35
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 9 27 15 29
rect 23 28 25 33
rect 35 28 37 33
rect 49 29 51 33
rect 13 24 15 27
rect 45 27 51 29
rect 45 24 47 27
rect 35 12 37 17
rect 45 12 47 17
rect 13 6 15 11
rect 23 6 25 11
<< ndif >>
rect 18 24 23 28
rect 4 11 13 24
rect 15 21 23 24
rect 15 19 18 21
rect 20 19 23 21
rect 15 11 23 19
rect 25 17 35 28
rect 37 24 42 28
rect 37 21 45 24
rect 37 19 40 21
rect 42 19 45 21
rect 37 17 45 19
rect 47 21 55 24
rect 47 19 50 21
rect 52 19 55 21
rect 47 17 55 19
rect 25 11 33 17
rect 4 9 7 11
rect 9 9 11 11
rect 4 7 11 9
rect 27 9 29 11
rect 31 9 33 11
rect 27 7 33 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 42 16 70
rect 18 68 26 70
rect 18 66 21 68
rect 23 66 26 68
rect 18 61 26 66
rect 18 59 21 61
rect 23 59 26 61
rect 18 42 26 59
rect 28 42 33 70
rect 35 61 43 70
rect 35 59 38 61
rect 40 59 43 61
rect 35 54 43 59
rect 35 52 38 54
rect 40 52 43 54
rect 35 42 43 52
rect 45 42 50 70
rect 52 68 60 70
rect 52 66 55 68
rect 57 66 60 68
rect 52 61 60 66
rect 52 59 55 61
rect 57 59 60 61
rect 52 42 60 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 37 61 41 63
rect 37 59 38 61
rect 40 59 41 61
rect 37 54 41 59
rect 2 53 38 54
rect 2 51 4 53
rect 6 52 38 53
rect 40 52 41 54
rect 6 51 41 52
rect 2 50 41 51
rect 2 46 6 50
rect 2 44 4 46
rect 2 22 6 44
rect 22 42 55 46
rect 22 37 28 42
rect 22 35 24 37
rect 26 35 28 37
rect 22 34 28 35
rect 33 37 39 38
rect 33 35 35 37
rect 37 35 39 37
rect 10 31 14 33
rect 10 29 11 31
rect 13 30 14 31
rect 33 30 39 35
rect 49 37 55 42
rect 49 35 51 37
rect 53 35 55 37
rect 49 34 55 35
rect 13 29 39 30
rect 10 26 39 29
rect 2 21 44 22
rect 2 19 18 21
rect 20 19 40 21
rect 42 19 44 21
rect 2 18 44 19
rect -2 11 66 12
rect -2 9 7 11
rect 9 9 29 11
rect 31 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 13 11 15 24
rect 23 11 25 28
rect 35 17 37 28
rect 45 17 47 24
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
<< polyct1 >>
rect 24 35 26 37
rect 35 35 37 37
rect 51 35 53 37
rect 11 29 13 31
<< ndifct0 >>
rect 50 19 52 21
<< ndifct1 >>
rect 18 19 20 21
rect 40 19 42 21
rect 7 9 9 11
rect 29 9 31 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 21 66 23 68
rect 21 59 23 61
rect 55 66 57 68
rect 55 59 57 61
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 38 59 40 61
rect 38 52 40 54
<< alu0 >>
rect 19 66 21 68
rect 23 66 25 68
rect 19 61 25 66
rect 53 66 55 68
rect 57 66 59 68
rect 19 59 21 61
rect 23 59 25 61
rect 19 58 25 59
rect 53 61 59 66
rect 53 59 55 61
rect 57 59 59 61
rect 53 58 59 59
rect 6 42 7 50
rect 49 21 53 23
rect 49 19 50 21
rect 52 19 53 21
rect 49 12 53 19
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 28 28 28 6 b
rlabel alu1 28 44 28 44 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 32 36 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 36 52 36 52 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 40 52 40 6 a
<< end >>
