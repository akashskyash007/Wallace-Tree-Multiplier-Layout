magic
tech scmos
timestamp 1199202821
<< ab >>
rect 0 0 144 72
<< nwell >>
rect -5 32 149 77
<< pwell >>
rect -5 -5 149 32
<< poly >>
rect 20 65 22 70
rect 30 65 32 70
rect 40 65 42 70
rect 50 65 52 70
rect 70 65 72 70
rect 80 65 82 70
rect 100 65 102 70
rect 110 65 112 70
rect 120 65 122 70
rect 20 35 22 38
rect 30 35 32 38
rect 40 35 42 38
rect 10 33 42 35
rect 10 31 12 33
rect 14 31 19 33
rect 21 31 42 33
rect 10 29 42 31
rect 10 26 12 29
rect 20 26 22 29
rect 30 26 32 29
rect 40 26 42 29
rect 50 35 52 38
rect 70 35 72 38
rect 80 35 82 38
rect 100 35 102 38
rect 110 35 112 38
rect 120 35 122 38
rect 50 33 92 35
rect 50 31 52 33
rect 54 31 59 33
rect 61 31 92 33
rect 50 29 92 31
rect 50 26 52 29
rect 60 26 62 29
rect 70 26 72 29
rect 80 26 82 29
rect 90 26 92 29
rect 100 33 132 35
rect 100 31 120 33
rect 122 31 128 33
rect 130 31 132 33
rect 100 29 132 31
rect 100 26 102 29
rect 110 26 112 29
rect 120 26 122 29
rect 130 26 132 29
rect 80 11 82 16
rect 90 11 92 16
rect 10 2 12 6
rect 20 2 22 6
rect 30 2 32 6
rect 40 2 42 6
rect 50 2 52 6
rect 60 2 62 6
rect 70 2 72 6
rect 100 2 102 6
rect 110 2 112 6
rect 120 2 122 6
rect 130 2 132 6
<< ndif >>
rect 3 24 10 26
rect 3 22 5 24
rect 7 22 10 24
rect 3 17 10 22
rect 3 15 5 17
rect 7 15 10 17
rect 3 13 10 15
rect 5 6 10 13
rect 12 17 20 26
rect 12 15 15 17
rect 17 15 20 17
rect 12 10 20 15
rect 12 8 15 10
rect 17 8 20 10
rect 12 6 20 8
rect 22 24 30 26
rect 22 22 25 24
rect 27 22 30 24
rect 22 17 30 22
rect 22 15 25 17
rect 27 15 30 17
rect 22 6 30 15
rect 32 10 40 26
rect 32 8 35 10
rect 37 8 40 10
rect 32 6 40 8
rect 42 17 50 26
rect 42 15 45 17
rect 47 15 50 17
rect 42 6 50 15
rect 52 24 60 26
rect 52 22 55 24
rect 57 22 60 24
rect 52 6 60 22
rect 62 17 70 26
rect 62 15 65 17
rect 67 15 70 17
rect 62 6 70 15
rect 72 24 80 26
rect 72 22 75 24
rect 77 22 80 24
rect 72 16 80 22
rect 82 20 90 26
rect 82 18 85 20
rect 87 18 90 20
rect 82 16 90 18
rect 92 24 100 26
rect 92 22 95 24
rect 97 22 100 24
rect 92 16 100 22
rect 72 6 77 16
rect 95 6 100 16
rect 102 24 110 26
rect 102 22 105 24
rect 107 22 110 24
rect 102 6 110 22
rect 112 16 120 26
rect 112 14 115 16
rect 117 14 120 16
rect 112 6 120 14
rect 122 24 130 26
rect 122 22 125 24
rect 127 22 130 24
rect 122 6 130 22
rect 132 24 139 26
rect 132 22 135 24
rect 137 22 139 24
rect 132 17 139 22
rect 132 15 135 17
rect 137 15 139 17
rect 132 13 139 15
rect 132 6 137 13
<< pdif >>
rect 13 63 20 65
rect 13 61 15 63
rect 17 61 20 63
rect 13 56 20 61
rect 13 54 15 56
rect 17 54 20 56
rect 13 38 20 54
rect 22 49 30 65
rect 22 47 25 49
rect 27 47 30 49
rect 22 42 30 47
rect 22 40 25 42
rect 27 40 30 42
rect 22 38 30 40
rect 32 63 40 65
rect 32 61 35 63
rect 37 61 40 63
rect 32 56 40 61
rect 32 54 35 56
rect 37 54 40 56
rect 32 38 40 54
rect 42 49 50 65
rect 42 47 45 49
rect 47 47 50 49
rect 42 42 50 47
rect 42 40 45 42
rect 47 40 50 42
rect 42 38 50 40
rect 52 63 70 65
rect 52 61 55 63
rect 57 61 65 63
rect 67 61 70 63
rect 52 56 70 61
rect 52 54 55 56
rect 57 54 65 56
rect 67 54 70 56
rect 52 38 70 54
rect 72 49 80 65
rect 72 47 75 49
rect 77 47 80 49
rect 72 42 80 47
rect 72 40 75 42
rect 77 40 80 42
rect 72 38 80 40
rect 82 63 89 65
rect 82 61 85 63
rect 87 61 89 63
rect 82 56 89 61
rect 82 54 85 56
rect 87 54 89 56
rect 82 38 89 54
rect 95 51 100 65
rect 93 49 100 51
rect 93 47 95 49
rect 97 47 100 49
rect 93 42 100 47
rect 93 40 95 42
rect 97 40 100 42
rect 93 38 100 40
rect 102 63 110 65
rect 102 61 105 63
rect 107 61 110 63
rect 102 56 110 61
rect 102 54 105 56
rect 107 54 110 56
rect 102 38 110 54
rect 112 49 120 65
rect 112 47 115 49
rect 117 47 120 49
rect 112 42 120 47
rect 112 40 115 42
rect 117 40 120 42
rect 112 38 120 40
rect 122 63 130 65
rect 122 61 125 63
rect 127 61 130 63
rect 122 56 130 61
rect 122 54 125 56
rect 127 54 130 56
rect 122 38 130 54
<< alu1 >>
rect -2 67 146 72
rect -2 65 5 67
rect 7 65 137 67
rect 139 65 146 67
rect -2 64 146 65
rect 2 34 6 51
rect 24 49 28 51
rect 24 47 25 49
rect 27 47 28 49
rect 24 42 28 47
rect 44 49 48 51
rect 44 47 45 49
rect 47 47 48 49
rect 44 42 48 47
rect 74 49 78 59
rect 74 47 75 49
rect 77 47 78 49
rect 74 42 78 47
rect 94 49 98 51
rect 94 47 95 49
rect 97 47 98 49
rect 94 42 98 47
rect 114 49 118 51
rect 114 47 115 49
rect 117 47 118 49
rect 114 42 118 47
rect 24 40 25 42
rect 27 40 45 42
rect 47 40 75 42
rect 77 40 95 42
rect 97 40 115 42
rect 117 40 118 42
rect 24 38 118 40
rect 2 33 23 34
rect 2 31 12 33
rect 14 31 19 33
rect 21 31 23 33
rect 2 29 23 31
rect 41 33 63 34
rect 41 31 52 33
rect 54 31 59 33
rect 61 31 63 33
rect 41 30 63 31
rect 41 22 47 30
rect 106 26 110 38
rect 129 34 135 42
rect 118 33 135 34
rect 118 31 120 33
rect 122 31 128 33
rect 130 31 135 33
rect 118 30 135 31
rect 103 24 129 26
rect 103 22 105 24
rect 107 22 125 24
rect 127 22 129 24
rect 103 21 129 22
rect -2 7 146 8
rect -2 5 85 7
rect 87 5 146 7
rect -2 0 146 5
<< ptie >>
rect 81 7 91 9
rect 81 5 85 7
rect 87 5 91 7
rect 81 3 91 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 135 67 141 69
rect 135 65 137 67
rect 139 65 141 67
rect 3 40 9 65
rect 135 40 141 65
<< nmos >>
rect 10 6 12 26
rect 20 6 22 26
rect 30 6 32 26
rect 40 6 42 26
rect 50 6 52 26
rect 60 6 62 26
rect 70 6 72 26
rect 80 16 82 26
rect 90 16 92 26
rect 100 6 102 26
rect 110 6 112 26
rect 120 6 122 26
rect 130 6 132 26
<< pmos >>
rect 20 38 22 65
rect 30 38 32 65
rect 40 38 42 65
rect 50 38 52 65
rect 70 38 72 65
rect 80 38 82 65
rect 100 38 102 65
rect 110 38 112 65
rect 120 38 122 65
<< polyct1 >>
rect 12 31 14 33
rect 19 31 21 33
rect 52 31 54 33
rect 59 31 61 33
rect 120 31 122 33
rect 128 31 130 33
<< ndifct0 >>
rect 5 22 7 24
rect 5 15 7 17
rect 15 15 17 17
rect 15 8 17 10
rect 25 22 27 24
rect 25 15 27 17
rect 35 8 37 10
rect 45 15 47 17
rect 55 22 57 24
rect 65 15 67 17
rect 75 22 77 24
rect 85 18 87 20
rect 95 22 97 24
rect 115 14 117 16
rect 135 22 137 24
rect 135 15 137 17
<< ndifct1 >>
rect 105 22 107 24
rect 125 22 127 24
<< ntiect1 >>
rect 5 65 7 67
rect 137 65 139 67
<< ptiect1 >>
rect 85 5 87 7
<< pdifct0 >>
rect 15 61 17 63
rect 15 54 17 56
rect 35 61 37 63
rect 35 54 37 56
rect 55 61 57 63
rect 65 61 67 63
rect 55 54 57 56
rect 65 54 67 56
rect 85 61 87 63
rect 85 54 87 56
rect 105 61 107 63
rect 105 54 107 56
rect 125 61 127 63
rect 125 54 127 56
<< pdifct1 >>
rect 25 47 27 49
rect 25 40 27 42
rect 45 47 47 49
rect 45 40 47 42
rect 75 47 77 49
rect 75 40 77 42
rect 95 47 97 49
rect 95 40 97 42
rect 115 47 117 49
rect 115 40 117 42
<< alu0 >>
rect 14 63 18 64
rect 14 61 15 63
rect 17 61 18 63
rect 14 56 18 61
rect 14 54 15 56
rect 17 54 18 56
rect 14 52 18 54
rect 34 63 38 64
rect 34 61 35 63
rect 37 61 38 63
rect 34 56 38 61
rect 34 54 35 56
rect 37 54 38 56
rect 34 52 38 54
rect 54 63 58 64
rect 54 61 55 63
rect 57 61 58 63
rect 54 56 58 61
rect 54 54 55 56
rect 57 54 58 56
rect 54 52 58 54
rect 64 63 68 64
rect 64 61 65 63
rect 67 61 68 63
rect 64 56 68 61
rect 84 63 88 64
rect 84 61 85 63
rect 87 61 88 63
rect 64 54 65 56
rect 67 54 68 56
rect 64 52 68 54
rect 84 56 88 61
rect 84 54 85 56
rect 87 54 88 56
rect 84 52 88 54
rect 104 63 108 64
rect 104 61 105 63
rect 107 61 108 63
rect 104 56 108 61
rect 104 54 105 56
rect 107 54 108 56
rect 104 52 108 54
rect 124 63 128 64
rect 124 61 125 63
rect 127 61 128 63
rect 124 56 128 61
rect 124 54 125 56
rect 127 54 128 56
rect 124 52 128 54
rect 4 24 28 26
rect 4 22 5 24
rect 7 22 25 24
rect 27 22 28 24
rect 75 26 98 30
rect 75 25 79 26
rect 53 24 79 25
rect 53 22 55 24
rect 57 22 75 24
rect 77 22 79 24
rect 94 24 98 26
rect 94 22 95 24
rect 97 22 98 24
rect 4 17 8 22
rect 24 18 28 22
rect 53 21 79 22
rect 84 20 88 22
rect 84 18 85 20
rect 87 18 88 20
rect 4 15 5 17
rect 7 15 8 17
rect 4 13 8 15
rect 13 17 19 18
rect 13 15 15 17
rect 17 15 19 17
rect 13 10 19 15
rect 24 17 88 18
rect 24 15 25 17
rect 27 15 45 17
rect 47 15 65 17
rect 67 15 88 17
rect 24 14 88 15
rect 94 17 98 22
rect 134 24 138 26
rect 134 22 135 24
rect 137 22 138 24
rect 134 17 138 22
rect 94 16 135 17
rect 94 14 115 16
rect 117 15 135 16
rect 137 15 138 17
rect 117 14 138 15
rect 94 13 138 14
rect 13 8 15 10
rect 17 8 19 10
rect 33 10 39 11
rect 33 8 35 10
rect 37 8 39 10
<< labels >>
rlabel alu0 6 19 6 19 6 n1
rlabel alu0 26 20 26 20 6 n1
rlabel alu0 56 16 56 16 6 n1
rlabel alu0 96 21 96 21 6 n2
rlabel alu0 66 23 66 23 6 n2
rlabel ndifct0 116 15 116 15 6 n2
rlabel alu0 136 19 136 19 6 n2
rlabel alu1 12 32 12 32 6 a
rlabel polyct1 20 32 20 32 6 a
rlabel alu1 4 40 4 40 6 a
rlabel alu1 52 32 52 32 6 b
rlabel alu1 44 28 44 28 6 b
rlabel alu1 28 40 28 40 6 z
rlabel alu1 44 40 44 40 6 z
rlabel alu1 52 40 52 40 6 z
rlabel alu1 36 40 36 40 6 z
rlabel alu1 72 4 72 4 6 vss
rlabel polyct1 60 32 60 32 6 b
rlabel alu1 60 40 60 40 6 z
rlabel alu1 84 40 84 40 6 z
rlabel alu1 68 40 68 40 6 z
rlabel pdifct1 76 48 76 48 6 z
rlabel alu1 72 68 72 68 6 vdd
rlabel alu1 108 32 108 32 6 z
rlabel alu1 92 40 92 40 6 z
rlabel alu1 100 40 100 40 6 z
rlabel alu1 116 24 116 24 6 z
rlabel alu1 124 24 124 24 6 z
rlabel alu1 124 32 124 32 6 c
rlabel alu1 132 36 132 36 6 c
rlabel pdifct1 116 48 116 48 6 z
<< end >>
