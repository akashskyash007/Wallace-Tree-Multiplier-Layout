magic
tech scmos
timestamp 1199202478
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 9 72 94 74
rect 9 62 11 72
rect 19 62 21 67
rect 29 62 31 67
rect 39 62 41 72
rect 50 64 52 68
rect 63 64 65 68
rect 73 64 75 68
rect 83 64 85 68
rect 92 65 94 72
rect 92 63 103 65
rect 101 60 103 63
rect 9 37 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 17 37 31 39
rect 39 37 41 42
rect 50 39 52 44
rect 63 41 65 44
rect 73 41 75 44
rect 63 39 75 41
rect 83 41 85 44
rect 83 39 97 41
rect 48 37 54 39
rect 17 35 19 37
rect 21 35 31 37
rect 48 35 50 37
rect 52 35 54 37
rect 17 33 35 35
rect 33 30 35 33
rect 45 33 54 35
rect 63 38 69 39
rect 63 36 65 38
rect 67 36 69 38
rect 63 34 69 36
rect 91 37 93 39
rect 95 37 97 39
rect 91 35 97 37
rect 101 35 103 44
rect 45 30 47 33
rect 66 30 68 34
rect 76 33 87 35
rect 76 30 78 33
rect 85 31 87 33
rect 101 33 110 35
rect 101 31 106 33
rect 108 31 110 33
rect 85 29 110 31
rect 96 26 98 29
rect 96 11 98 16
rect 33 6 35 10
rect 45 6 47 10
rect 66 6 68 10
rect 76 6 78 10
<< ndif >>
rect 24 21 33 30
rect 24 19 27 21
rect 29 19 33 21
rect 24 14 33 19
rect 24 12 27 14
rect 29 12 33 14
rect 24 10 33 12
rect 35 21 45 30
rect 35 19 38 21
rect 40 19 45 21
rect 35 10 45 19
rect 47 28 54 30
rect 47 26 50 28
rect 52 26 54 28
rect 47 21 54 26
rect 47 19 50 21
rect 52 19 54 21
rect 47 17 54 19
rect 47 10 52 17
rect 58 14 66 30
rect 58 12 61 14
rect 63 12 66 14
rect 58 10 66 12
rect 68 28 76 30
rect 68 26 71 28
rect 73 26 76 28
rect 68 10 76 26
rect 78 23 83 30
rect 89 24 96 26
rect 78 21 85 23
rect 78 19 81 21
rect 83 19 85 21
rect 89 22 91 24
rect 93 22 96 24
rect 89 20 96 22
rect 78 17 85 19
rect 78 10 83 17
rect 91 16 96 20
rect 98 16 107 26
rect 100 11 107 16
rect 100 9 102 11
rect 104 9 107 11
rect 100 7 107 9
<< pdif >>
rect 43 62 50 64
rect 4 55 9 62
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 46 19 62
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 60 29 62
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 46 39 62
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 60 45 62
rect 47 60 50 62
rect 41 44 50 60
rect 52 48 63 64
rect 52 46 58 48
rect 60 46 63 48
rect 52 44 63 46
rect 65 62 73 64
rect 65 60 68 62
rect 70 60 73 62
rect 65 44 73 60
rect 75 48 83 64
rect 75 46 78 48
rect 80 46 83 48
rect 75 44 83 46
rect 85 50 90 64
rect 94 58 101 60
rect 94 56 96 58
rect 98 56 101 58
rect 94 54 101 56
rect 85 48 92 50
rect 85 46 88 48
rect 90 46 92 48
rect 85 44 92 46
rect 96 44 101 54
rect 103 58 110 60
rect 103 56 106 58
rect 108 56 110 58
rect 103 50 110 56
rect 103 48 106 50
rect 108 48 110 50
rect 103 44 110 48
rect 41 42 46 44
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 68 114 79
rect 42 62 49 63
rect 42 60 45 62
rect 47 60 49 62
rect 42 59 49 60
rect 42 54 46 59
rect 2 53 46 54
rect 2 51 4 53
rect 6 51 46 53
rect 2 50 46 51
rect 2 46 7 50
rect 2 44 4 46
rect 6 44 7 46
rect 2 41 7 44
rect 18 37 22 39
rect 18 35 19 37
rect 21 35 22 37
rect 18 23 22 35
rect 10 17 22 23
rect 42 30 46 50
rect 85 48 92 49
rect 85 46 88 48
rect 90 46 92 48
rect 85 45 92 46
rect 57 38 70 39
rect 57 36 65 38
rect 67 36 70 38
rect 57 33 70 36
rect 42 28 53 30
rect 42 26 50 28
rect 52 26 53 28
rect 57 26 63 33
rect 85 39 89 45
rect 42 25 53 26
rect 82 35 89 39
rect 48 22 53 25
rect 82 22 86 35
rect 48 21 86 22
rect 48 19 50 21
rect 52 19 81 21
rect 83 19 86 21
rect 105 33 110 39
rect 105 31 106 33
rect 108 31 110 33
rect 105 23 110 31
rect 48 18 86 19
rect 98 17 110 23
rect -2 11 114 12
rect -2 9 102 11
rect 104 9 114 11
rect -2 1 114 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 33 10 35 30
rect 45 10 47 30
rect 66 10 68 30
rect 76 10 78 30
rect 96 16 98 26
<< pmos >>
rect 9 42 11 62
rect 19 42 21 62
rect 29 42 31 62
rect 39 42 41 62
rect 50 44 52 64
rect 63 44 65 64
rect 73 44 75 64
rect 83 44 85 64
rect 101 44 103 60
<< polyct0 >>
rect 50 35 52 37
rect 93 37 95 39
<< polyct1 >>
rect 19 35 21 37
rect 65 36 67 38
rect 106 31 108 33
<< ndifct0 >>
rect 27 19 29 21
rect 27 12 29 14
rect 38 19 40 21
rect 61 12 63 14
rect 71 26 73 28
rect 91 22 93 24
<< ndifct1 >>
rect 50 26 52 28
rect 50 19 52 21
rect 81 19 83 21
rect 102 9 104 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 14 44 16 46
rect 24 58 26 60
rect 34 44 36 46
rect 58 46 60 48
rect 68 60 70 62
rect 78 46 80 48
rect 96 56 98 58
rect 106 56 108 58
rect 106 48 108 50
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 45 60 47 62
rect 88 46 90 48
<< alu0 >>
rect 22 60 28 68
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 66 62 72 68
rect 66 60 68 62
rect 70 60 72 62
rect 66 59 72 60
rect 95 58 99 60
rect 95 56 96 58
rect 98 56 99 58
rect 12 46 38 47
rect 12 44 14 46
rect 16 44 34 46
rect 36 44 38 46
rect 12 43 38 44
rect 26 21 30 23
rect 26 19 27 21
rect 29 19 30 21
rect 26 14 30 19
rect 34 22 38 43
rect 49 52 99 56
rect 49 37 53 52
rect 56 48 82 49
rect 56 46 58 48
rect 60 46 78 48
rect 80 46 82 48
rect 56 45 82 46
rect 49 35 50 37
rect 52 35 53 37
rect 49 33 53 35
rect 74 29 78 45
rect 95 41 99 52
rect 105 58 109 68
rect 105 56 106 58
rect 108 56 109 58
rect 105 50 109 56
rect 105 48 106 50
rect 108 48 109 50
rect 105 46 109 48
rect 69 28 78 29
rect 69 26 71 28
rect 73 26 78 28
rect 69 25 78 26
rect 92 39 99 41
rect 92 37 93 39
rect 95 37 99 39
rect 92 30 96 37
rect 34 21 42 22
rect 34 19 38 21
rect 40 19 42 21
rect 34 18 42 19
rect 90 26 96 30
rect 90 24 94 26
rect 90 22 91 24
rect 93 22 94 24
rect 90 20 94 22
rect 26 12 27 14
rect 29 12 30 14
rect 59 14 65 15
rect 59 12 61 14
rect 63 12 65 14
<< labels >>
rlabel alu0 51 44 51 44 6 sn
rlabel alu0 36 32 36 32 6 a0n
rlabel alu0 25 45 25 45 6 a0n
rlabel alu0 73 27 73 27 6 a1n
rlabel alu0 69 47 69 47 6 a1n
rlabel alu0 92 25 92 25 6 sn
rlabel alu0 97 48 97 48 6 sn
rlabel alu0 94 33 94 33 6 sn
rlabel alu1 12 20 12 20 6 a0
rlabel alu1 20 28 20 28 6 a0
rlabel alu1 4 44 4 44 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 44 44 44 44 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 56 6 56 6 6 vss
rlabel alu1 68 20 68 20 6 z
rlabel alu1 76 20 76 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 60 32 60 32 6 a1
rlabel alu1 68 36 68 36 6 a1
rlabel alu1 56 74 56 74 6 vdd
rlabel alu1 100 20 100 20 6 s
rlabel alu1 84 32 84 32 6 z
rlabel alu1 108 28 108 28 6 s
<< end >>
