magic
tech scmos
timestamp 1199543043
<< ab >>
rect 0 0 170 100
<< nwell >>
rect -5 48 175 105
<< pwell >>
rect -5 -5 175 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 47 94 49 98
rect 59 94 61 98
rect 71 94 73 98
rect 83 94 85 98
rect 109 94 111 98
rect 121 94 123 98
rect 133 94 135 98
rect 145 94 147 98
rect 11 53 13 56
rect 7 51 13 53
rect 7 49 9 51
rect 11 49 13 51
rect 7 47 13 49
rect 11 25 13 47
rect 23 53 25 56
rect 47 53 49 56
rect 59 53 61 56
rect 71 53 73 56
rect 83 53 85 56
rect 157 75 159 79
rect 23 51 33 53
rect 23 49 29 51
rect 31 49 33 51
rect 23 47 33 49
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 57 51 63 53
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 67 51 73 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 77 51 85 53
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 23 25 25 47
rect 51 25 53 47
rect 59 25 61 47
rect 71 25 73 47
rect 79 25 81 47
rect 109 43 111 55
rect 121 43 123 55
rect 107 41 113 43
rect 107 39 109 41
rect 111 39 113 41
rect 107 37 113 39
rect 121 41 127 43
rect 121 39 123 41
rect 125 39 127 41
rect 121 37 127 39
rect 133 41 135 55
rect 145 43 147 55
rect 145 41 153 43
rect 133 39 149 41
rect 151 39 153 41
rect 109 29 111 37
rect 109 27 115 29
rect 113 24 115 27
rect 121 24 123 37
rect 133 25 135 39
rect 145 37 153 39
rect 145 25 147 37
rect 157 33 159 55
rect 151 31 159 33
rect 151 29 153 31
rect 155 29 159 31
rect 151 27 159 29
rect 157 24 159 27
rect 157 10 159 14
rect 11 2 13 6
rect 23 2 25 6
rect 51 2 53 6
rect 59 2 61 6
rect 71 2 73 6
rect 79 2 81 6
rect 113 2 115 6
rect 121 2 123 6
rect 133 2 135 6
rect 145 2 147 6
<< ndif >>
rect 3 11 11 25
rect 3 9 5 11
rect 7 9 11 11
rect 3 6 11 9
rect 13 6 23 25
rect 25 21 33 25
rect 25 19 29 21
rect 31 19 33 21
rect 25 6 33 19
rect 43 11 51 25
rect 43 9 45 11
rect 47 9 51 11
rect 43 6 51 9
rect 53 6 59 25
rect 61 21 71 25
rect 61 19 65 21
rect 67 19 71 21
rect 61 6 71 19
rect 73 6 79 25
rect 81 11 89 25
rect 137 31 143 33
rect 137 29 139 31
rect 141 29 143 31
rect 137 25 143 29
rect 128 24 133 25
rect 81 9 85 11
rect 87 9 89 11
rect 81 6 89 9
rect 105 21 113 24
rect 105 19 107 21
rect 109 19 113 21
rect 105 6 113 19
rect 115 6 121 24
rect 123 11 133 24
rect 123 9 127 11
rect 129 9 133 11
rect 123 6 133 9
rect 135 6 145 25
rect 147 24 152 25
rect 147 14 157 24
rect 159 21 167 24
rect 159 19 163 21
rect 165 19 167 21
rect 159 14 167 19
rect 147 11 155 14
rect 147 9 151 11
rect 153 9 155 11
rect 147 6 155 9
<< pdif >>
rect 3 81 11 94
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 56 11 69
rect 13 71 23 94
rect 13 69 17 71
rect 19 69 23 71
rect 13 56 23 69
rect 25 81 33 94
rect 25 79 29 81
rect 31 79 33 81
rect 25 71 33 79
rect 25 69 29 71
rect 31 69 33 71
rect 25 56 33 69
rect 39 81 47 94
rect 39 79 41 81
rect 43 79 47 81
rect 39 56 47 79
rect 49 71 59 94
rect 49 69 53 71
rect 55 69 59 71
rect 49 56 59 69
rect 61 81 71 94
rect 61 79 65 81
rect 67 79 71 81
rect 61 71 71 79
rect 61 69 65 71
rect 67 69 71 71
rect 61 56 71 69
rect 73 71 83 94
rect 73 69 77 71
rect 79 69 83 71
rect 73 56 83 69
rect 85 81 93 94
rect 85 79 89 81
rect 91 79 93 81
rect 85 56 93 79
rect 101 91 109 94
rect 101 89 103 91
rect 105 89 109 91
rect 101 81 109 89
rect 101 79 103 81
rect 105 79 109 81
rect 101 55 109 79
rect 111 81 121 94
rect 111 79 115 81
rect 117 79 121 81
rect 111 55 121 79
rect 123 91 133 94
rect 123 89 127 91
rect 129 89 133 91
rect 123 81 133 89
rect 123 79 127 81
rect 129 79 133 81
rect 123 55 133 79
rect 135 81 145 94
rect 135 79 139 81
rect 141 79 145 81
rect 135 71 145 79
rect 135 69 139 71
rect 141 69 145 71
rect 135 61 145 69
rect 135 59 139 61
rect 141 59 145 61
rect 135 55 145 59
rect 147 91 155 94
rect 147 89 151 91
rect 153 89 155 91
rect 147 81 155 89
rect 147 79 151 81
rect 153 79 155 81
rect 147 75 155 79
rect 147 71 157 75
rect 147 69 151 71
rect 153 69 157 71
rect 147 55 157 69
rect 159 71 167 75
rect 159 69 163 71
rect 165 69 167 71
rect 159 59 167 69
rect 159 57 163 59
rect 165 57 167 59
rect 159 55 167 57
<< alu1 >>
rect -2 93 172 100
rect -2 91 163 93
rect 165 91 172 93
rect -2 89 103 91
rect 105 89 127 91
rect 129 89 151 91
rect 153 89 172 91
rect -2 88 172 89
rect 4 82 8 83
rect 28 82 32 83
rect 4 81 32 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 32 81
rect 4 78 32 79
rect 39 81 93 82
rect 39 79 41 81
rect 43 79 65 81
rect 67 79 89 81
rect 91 79 93 81
rect 39 78 93 79
rect 102 81 106 88
rect 102 79 103 81
rect 105 79 106 81
rect 4 71 8 78
rect 28 72 32 78
rect 4 69 5 71
rect 7 69 8 71
rect 4 67 8 69
rect 15 71 22 72
rect 15 69 17 71
rect 19 69 22 71
rect 15 68 22 69
rect 8 51 12 63
rect 8 49 9 51
rect 11 49 12 51
rect 8 17 12 49
rect 18 22 22 68
rect 28 71 57 72
rect 28 69 29 71
rect 31 69 53 71
rect 55 69 57 71
rect 28 68 57 69
rect 64 71 68 78
rect 102 77 106 79
rect 114 81 118 83
rect 114 79 115 81
rect 117 79 118 81
rect 114 72 118 79
rect 126 81 130 88
rect 126 79 127 81
rect 129 79 130 81
rect 126 77 130 79
rect 138 81 142 83
rect 138 79 139 81
rect 141 79 142 81
rect 64 69 65 71
rect 67 69 68 71
rect 28 67 32 68
rect 64 67 68 69
rect 75 71 118 72
rect 75 69 77 71
rect 79 69 118 71
rect 75 68 118 69
rect 28 51 32 63
rect 28 49 29 51
rect 31 49 32 51
rect 28 27 32 49
rect 48 51 52 63
rect 48 49 49 51
rect 51 49 52 51
rect 48 27 52 49
rect 58 51 62 63
rect 58 49 59 51
rect 61 49 62 51
rect 58 27 62 49
rect 68 51 72 63
rect 68 49 69 51
rect 71 49 72 51
rect 68 27 72 49
rect 78 51 82 63
rect 78 49 79 51
rect 81 49 82 51
rect 78 27 82 49
rect 108 41 112 63
rect 128 42 132 73
rect 108 39 109 41
rect 111 39 112 41
rect 108 27 112 39
rect 121 41 132 42
rect 121 39 123 41
rect 125 39 132 41
rect 121 38 132 39
rect 128 27 132 38
rect 138 71 142 79
rect 138 69 139 71
rect 141 69 142 71
rect 138 61 142 69
rect 150 81 154 88
rect 150 79 151 81
rect 153 79 154 81
rect 150 71 154 79
rect 150 69 151 71
rect 153 69 154 71
rect 150 67 154 69
rect 162 71 166 73
rect 162 69 163 71
rect 165 69 166 71
rect 138 59 139 61
rect 141 59 142 61
rect 138 31 142 59
rect 162 59 166 69
rect 162 57 163 59
rect 165 57 166 59
rect 162 42 166 57
rect 147 41 166 42
rect 147 39 149 41
rect 151 39 166 41
rect 147 38 166 39
rect 138 29 139 31
rect 141 29 142 31
rect 138 27 142 29
rect 152 31 156 33
rect 152 29 153 31
rect 155 29 156 31
rect 152 22 156 29
rect 18 21 156 22
rect 18 19 29 21
rect 31 19 65 21
rect 67 19 107 21
rect 109 19 156 21
rect 18 18 156 19
rect 162 21 166 38
rect 162 19 163 21
rect 165 19 166 21
rect 162 17 166 19
rect -2 11 172 12
rect -2 9 5 11
rect 7 9 45 11
rect 47 9 85 11
rect 87 9 127 11
rect 129 9 151 11
rect 153 9 172 11
rect -2 0 172 9
<< ntie >>
rect 161 93 167 95
rect 161 91 163 93
rect 165 91 167 93
rect 161 84 167 91
<< nmos >>
rect 11 6 13 25
rect 23 6 25 25
rect 51 6 53 25
rect 59 6 61 25
rect 71 6 73 25
rect 79 6 81 25
rect 113 6 115 24
rect 121 6 123 24
rect 133 6 135 25
rect 145 6 147 25
rect 157 14 159 24
<< pmos >>
rect 11 56 13 94
rect 23 56 25 94
rect 47 56 49 94
rect 59 56 61 94
rect 71 56 73 94
rect 83 56 85 94
rect 109 55 111 94
rect 121 55 123 94
rect 133 55 135 94
rect 145 55 147 94
rect 157 55 159 75
<< polyct1 >>
rect 9 49 11 51
rect 29 49 31 51
rect 49 49 51 51
rect 59 49 61 51
rect 69 49 71 51
rect 79 49 81 51
rect 109 39 111 41
rect 123 39 125 41
rect 149 39 151 41
rect 153 29 155 31
<< ndifct1 >>
rect 5 9 7 11
rect 29 19 31 21
rect 45 9 47 11
rect 65 19 67 21
rect 139 29 141 31
rect 85 9 87 11
rect 107 19 109 21
rect 127 9 129 11
rect 163 19 165 21
rect 151 9 153 11
<< ntiect1 >>
rect 163 91 165 93
<< pdifct1 >>
rect 5 79 7 81
rect 5 69 7 71
rect 17 69 19 71
rect 29 79 31 81
rect 29 69 31 71
rect 41 79 43 81
rect 53 69 55 71
rect 65 79 67 81
rect 65 69 67 71
rect 77 69 79 71
rect 89 79 91 81
rect 103 89 105 91
rect 103 79 105 81
rect 115 79 117 81
rect 127 89 129 91
rect 127 79 129 81
rect 139 79 141 81
rect 139 69 141 71
rect 139 59 141 61
rect 151 89 153 91
rect 151 79 153 81
rect 151 69 153 71
rect 163 69 165 71
rect 163 57 165 59
<< labels >>
rlabel alu1 30 45 30 45 6 i6
rlabel alu1 10 40 10 40 6 i7
rlabel alu1 80 45 80 45 6 i2
rlabel alu1 70 45 70 45 6 i3
rlabel alu1 60 45 60 45 6 i4
rlabel alu1 50 45 50 45 6 i5
rlabel alu1 85 6 85 6 6 vss
rlabel alu1 110 45 110 45 6 i1
rlabel alu1 85 94 85 94 6 vdd
rlabel alu1 130 50 130 50 6 i0
rlabel alu1 140 55 140 55 6 nq
<< end >>
