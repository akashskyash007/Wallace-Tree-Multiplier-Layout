magic
tech scmos
timestamp 1199201996
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 56 41 61
rect 49 56 51 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 9 33 31 35
rect 14 31 27 33
rect 29 31 31 33
rect 14 29 31 31
rect 37 33 51 35
rect 37 31 43 33
rect 45 31 47 33
rect 37 29 47 31
rect 14 26 16 29
rect 24 26 26 29
rect 37 26 39 29
rect 14 2 16 6
rect 24 2 26 6
rect 37 2 39 7
<< ndif >>
rect 6 17 14 26
rect 6 15 9 17
rect 11 15 14 17
rect 6 10 14 15
rect 6 8 9 10
rect 11 8 14 10
rect 6 6 14 8
rect 16 24 24 26
rect 16 22 19 24
rect 21 22 24 24
rect 16 17 24 22
rect 16 15 19 17
rect 21 15 24 17
rect 16 6 24 15
rect 26 17 37 26
rect 26 15 31 17
rect 33 15 37 17
rect 26 10 37 15
rect 26 8 31 10
rect 33 8 37 10
rect 26 7 37 8
rect 39 24 46 26
rect 39 22 42 24
rect 44 22 46 24
rect 39 17 46 22
rect 39 15 42 17
rect 44 15 46 17
rect 39 13 46 15
rect 39 7 44 13
rect 26 6 35 7
<< pdif >>
rect 4 51 9 65
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 62 19 65
rect 11 60 14 62
rect 16 60 19 62
rect 11 54 19 60
rect 11 52 14 54
rect 16 52 19 54
rect 11 38 19 52
rect 21 49 29 65
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 56 37 65
rect 31 54 39 56
rect 31 52 34 54
rect 36 52 39 54
rect 31 38 39 52
rect 41 49 49 56
rect 41 47 44 49
rect 46 47 49 49
rect 41 42 49 47
rect 41 40 44 42
rect 46 40 49 42
rect 41 38 49 40
rect 51 54 58 56
rect 51 52 54 54
rect 56 52 58 54
rect 51 46 58 52
rect 51 44 54 46
rect 56 44 58 46
rect 51 38 58 44
<< alu1 >>
rect -2 67 66 72
rect -2 65 45 67
rect 47 65 53 67
rect 55 65 66 67
rect -2 64 66 65
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 23 49 27 51
rect 23 47 24 49
rect 26 47 27 49
rect 23 42 27 47
rect 2 40 4 42
rect 6 40 24 42
rect 26 40 27 42
rect 2 38 27 40
rect 2 37 14 38
rect 9 26 14 37
rect 41 33 55 34
rect 41 31 43 33
rect 45 31 55 33
rect 41 30 55 31
rect 9 24 23 26
rect 9 22 19 24
rect 21 22 23 24
rect 49 22 55 30
rect 18 17 23 22
rect 18 15 19 17
rect 21 15 23 17
rect 18 13 23 15
rect -2 7 66 8
rect -2 5 53 7
rect 55 5 66 7
rect -2 0 66 5
<< ptie >>
rect 51 7 57 24
rect 51 5 53 7
rect 55 5 57 7
rect 51 3 57 5
<< ntie >>
rect 43 67 57 69
rect 43 65 45 67
rect 47 65 53 67
rect 55 65 57 67
rect 43 63 57 65
<< nmos >>
rect 14 6 16 26
rect 24 6 26 26
rect 37 7 39 26
<< pmos >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 56
rect 49 38 51 56
<< polyct0 >>
rect 27 31 29 33
<< polyct1 >>
rect 43 31 45 33
<< ndifct0 >>
rect 9 15 11 17
rect 9 8 11 10
rect 31 15 33 17
rect 31 8 33 10
rect 42 22 44 24
rect 42 15 44 17
<< ndifct1 >>
rect 19 22 21 24
rect 19 15 21 17
<< ntiect1 >>
rect 45 65 47 67
rect 53 65 55 67
<< ptiect1 >>
rect 53 5 55 7
<< pdifct0 >>
rect 14 60 16 62
rect 14 52 16 54
rect 34 52 36 54
rect 44 47 46 49
rect 44 40 46 42
rect 54 52 56 54
rect 54 44 56 46
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 24 47 26 49
rect 24 40 26 42
<< alu0 >>
rect 13 62 17 64
rect 13 60 14 62
rect 16 60 17 62
rect 13 54 17 60
rect 13 52 14 54
rect 16 52 17 54
rect 13 50 17 52
rect 33 54 37 64
rect 33 52 34 54
rect 36 52 37 54
rect 33 50 37 52
rect 53 54 57 64
rect 53 52 54 54
rect 56 52 57 54
rect 43 49 47 51
rect 43 47 44 49
rect 46 47 47 49
rect 43 42 47 47
rect 53 46 57 52
rect 53 44 54 46
rect 56 44 57 46
rect 53 42 57 44
rect 33 40 44 42
rect 46 40 47 42
rect 33 38 47 40
rect 33 34 37 38
rect 25 33 37 34
rect 25 31 27 33
rect 29 31 37 33
rect 25 30 37 31
rect 33 26 37 30
rect 33 24 45 26
rect 33 22 42 24
rect 44 22 45 24
rect 7 17 13 18
rect 7 15 9 17
rect 11 15 13 17
rect 7 10 13 15
rect 29 17 35 18
rect 29 15 31 17
rect 33 15 35 17
rect 7 8 9 10
rect 11 8 13 10
rect 29 10 35 15
rect 41 17 45 22
rect 41 15 42 17
rect 44 15 45 17
rect 41 13 45 15
rect 29 8 31 10
rect 33 8 35 10
<< labels >>
rlabel alu0 31 32 31 32 6 an
rlabel alu0 43 19 43 19 6 an
rlabel alu0 45 44 45 44 6 an
rlabel alu1 12 32 12 32 6 z
rlabel alu1 4 44 4 44 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel polyct1 44 32 44 32 6 a
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 28 52 28 6 a
<< end >>
