magic
tech scmos
timestamp 1199447821
<< ab >>
rect -13 0 317 72
<< alu1 >>
rect -10 65 -6 70
rect -10 63 -9 65
rect -7 63 -6 65
rect -10 49 -6 63
rect -10 47 -9 49
rect -7 47 -6 49
rect -10 33 -6 47
rect -10 31 -9 33
rect -7 31 -6 33
rect -10 17 -6 31
rect -10 15 -9 17
rect -7 15 -6 17
rect -10 8 -6 15
rect -12 4 316 8
rect -10 2 -6 4
<< alu2 >>
rect -13 65 317 66
rect -13 63 -9 65
rect -7 63 317 65
rect -13 62 317 63
rect -13 49 317 50
rect -13 47 -9 49
rect -7 47 317 49
rect -13 46 317 47
rect -13 33 317 34
rect -13 31 -9 33
rect -7 31 317 33
rect -13 30 317 31
rect -13 17 317 18
rect -13 15 -9 17
rect -7 15 3 17
rect 5 15 19 17
rect 21 15 35 17
rect 37 15 51 17
rect 53 15 67 17
rect 69 15 83 17
rect 85 15 99 17
rect 101 15 115 17
rect 117 15 131 17
rect 133 15 147 17
rect 149 15 163 17
rect 165 15 179 17
rect 181 15 195 17
rect 197 15 211 17
rect 213 15 227 17
rect 229 15 243 17
rect 245 15 259 17
rect 261 15 275 17
rect 277 15 291 17
rect 293 15 307 17
rect 309 15 317 17
rect -13 14 317 15
<< alu3 >>
rect 2 57 6 70
rect 2 55 3 57
rect 5 55 6 57
rect 2 41 6 55
rect 2 39 3 41
rect 5 39 6 41
rect 2 25 6 39
rect 2 23 3 25
rect 5 23 6 25
rect 2 17 6 23
rect 2 15 3 17
rect 5 15 6 17
rect 2 9 6 15
rect 2 7 3 9
rect 5 7 6 9
rect 2 2 6 7
rect 18 17 22 70
rect 18 15 19 17
rect 21 15 22 17
rect 18 2 22 15
rect 34 17 38 70
rect 34 15 35 17
rect 37 15 38 17
rect 34 2 38 15
rect 50 17 54 70
rect 50 15 51 17
rect 53 15 54 17
rect 50 2 54 15
rect 66 17 70 70
rect 66 15 67 17
rect 69 15 70 17
rect 66 2 70 15
rect 82 17 86 70
rect 82 15 83 17
rect 85 15 86 17
rect 82 2 86 15
rect 98 17 102 70
rect 98 15 99 17
rect 101 15 102 17
rect 98 2 102 15
rect 114 17 118 70
rect 114 15 115 17
rect 117 15 118 17
rect 114 2 118 15
rect 130 17 134 70
rect 130 15 131 17
rect 133 15 134 17
rect 130 2 134 15
rect 146 17 150 70
rect 146 15 147 17
rect 149 15 150 17
rect 146 2 150 15
rect 162 17 166 70
rect 162 15 163 17
rect 165 15 166 17
rect 162 2 166 15
rect 178 17 182 70
rect 178 15 179 17
rect 181 15 182 17
rect 178 2 182 15
rect 194 17 198 70
rect 194 15 195 17
rect 197 15 198 17
rect 194 2 198 15
rect 210 17 214 70
rect 210 15 211 17
rect 213 15 214 17
rect 210 2 214 15
rect 226 17 230 70
rect 226 15 227 17
rect 229 15 230 17
rect 226 2 230 15
rect 242 17 246 70
rect 242 15 243 17
rect 245 15 246 17
rect 242 2 246 15
rect 258 17 262 70
rect 258 15 259 17
rect 261 15 262 17
rect 258 2 262 15
rect 274 17 278 70
rect 274 15 275 17
rect 277 15 278 17
rect 274 2 278 15
rect 290 17 294 70
rect 290 15 291 17
rect 293 15 294 17
rect 290 2 294 15
rect 306 17 310 70
rect 306 15 307 17
rect 309 15 310 17
rect 306 2 310 15
<< alu4 >>
rect -13 57 317 58
rect -13 55 3 57
rect 5 55 317 57
rect -13 54 317 55
rect -13 41 317 42
rect -13 39 3 41
rect 5 39 317 41
rect -13 38 317 39
rect -13 25 317 26
rect -13 23 3 25
rect 5 23 317 25
rect -13 22 317 23
rect -13 9 317 10
rect -13 7 -5 9
rect -3 7 3 9
rect 5 7 11 9
rect 13 7 27 9
rect 29 7 43 9
rect 45 7 59 9
rect 61 7 75 9
rect 77 7 91 9
rect 93 7 107 9
rect 109 7 123 9
rect 125 7 139 9
rect 141 7 155 9
rect 157 7 171 9
rect 173 7 187 9
rect 189 7 203 9
rect 205 7 219 9
rect 221 7 235 9
rect 237 7 251 9
rect 253 7 267 9
rect 269 7 283 9
rect 285 7 299 9
rect 301 7 317 9
rect -13 6 317 7
<< alu5 >>
rect -6 9 -2 70
rect -6 7 -5 9
rect -3 7 -2 9
rect -6 2 -2 7
rect 10 9 14 70
rect 10 7 11 9
rect 13 7 14 9
rect 10 2 14 7
rect 26 9 30 70
rect 26 7 27 9
rect 29 7 30 9
rect 26 2 30 7
rect 42 9 46 70
rect 42 7 43 9
rect 45 7 46 9
rect 42 2 46 7
rect 58 9 62 70
rect 58 7 59 9
rect 61 7 62 9
rect 58 2 62 7
rect 74 9 78 70
rect 74 7 75 9
rect 77 7 78 9
rect 74 2 78 7
rect 90 9 94 70
rect 90 7 91 9
rect 93 7 94 9
rect 90 2 94 7
rect 106 9 110 70
rect 106 7 107 9
rect 109 7 110 9
rect 106 2 110 7
rect 122 9 126 70
rect 122 7 123 9
rect 125 7 126 9
rect 122 2 126 7
rect 138 9 142 70
rect 138 7 139 9
rect 141 7 142 9
rect 138 2 142 7
rect 154 9 158 70
rect 154 7 155 9
rect 157 7 158 9
rect 154 2 158 7
rect 170 9 174 70
rect 170 7 171 9
rect 173 7 174 9
rect 170 2 174 7
rect 186 9 190 70
rect 186 7 187 9
rect 189 7 190 9
rect 186 2 190 7
rect 202 9 206 70
rect 202 7 203 9
rect 205 7 206 9
rect 202 2 206 7
rect 218 9 222 70
rect 218 7 219 9
rect 221 7 222 9
rect 218 2 222 7
rect 234 9 238 70
rect 234 7 235 9
rect 237 7 238 9
rect 234 2 238 7
rect 250 9 254 70
rect 250 7 251 9
rect 253 7 254 9
rect 250 2 254 7
rect 266 9 270 70
rect 266 7 267 9
rect 269 7 270 9
rect 266 2 270 7
rect 282 9 286 70
rect 282 7 283 9
rect 285 7 286 9
rect 282 2 286 7
rect 298 9 302 70
rect 298 7 299 9
rect 301 7 302 9
rect 298 2 302 7
<< via1 >>
rect -9 63 -7 65
rect -9 47 -7 49
rect -9 31 -7 33
rect -9 15 -7 17
<< via2 >>
rect 3 15 5 17
rect 19 15 21 17
rect 35 15 37 17
rect 51 15 53 17
rect 67 15 69 17
rect 83 15 85 17
rect 99 15 101 17
rect 115 15 117 17
rect 131 15 133 17
rect 147 15 149 17
rect 163 15 165 17
rect 179 15 181 17
rect 195 15 197 17
rect 211 15 213 17
rect 227 15 229 17
rect 243 15 245 17
rect 259 15 261 17
rect 275 15 277 17
rect 291 15 293 17
rect 307 15 309 17
<< via3 >>
rect 3 55 5 57
rect 3 39 5 41
rect 3 23 5 25
rect 3 7 5 9
<< via4 >>
rect -5 7 -3 9
rect 11 7 13 9
rect 27 7 29 9
rect 43 7 45 9
rect 59 7 61 9
rect 75 7 77 9
rect 91 7 93 9
rect 107 7 109 9
rect 123 7 125 9
rect 139 7 141 9
rect 155 7 157 9
rect 171 7 173 9
rect 187 7 189 9
rect 203 7 205 9
rect 219 7 221 9
rect 235 7 237 9
rect 251 7 253 9
rect 267 7 269 9
rect 283 7 285 9
rect 299 7 301 9
<< end >>
