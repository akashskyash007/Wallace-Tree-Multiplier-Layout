magic
tech scmos
timestamp 1199201922
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 54 11 59
rect 19 54 21 59
rect 30 55 32 60
rect 40 55 42 60
rect 9 29 11 46
rect 19 43 21 46
rect 19 41 25 43
rect 19 39 21 41
rect 23 39 25 41
rect 19 37 25 39
rect 9 27 15 29
rect 9 25 11 27
rect 13 25 15 27
rect 9 23 15 25
rect 12 20 14 23
rect 19 20 21 37
rect 30 29 32 46
rect 40 43 42 46
rect 39 41 47 43
rect 39 39 43 41
rect 45 39 47 41
rect 39 37 47 39
rect 25 27 34 29
rect 25 25 27 27
rect 29 25 34 27
rect 25 23 34 25
rect 32 20 34 23
rect 39 20 41 37
rect 12 8 14 13
rect 19 8 21 13
rect 32 8 34 13
rect 39 8 41 13
<< ndif >>
rect 5 18 12 20
rect 5 16 7 18
rect 9 16 12 18
rect 5 13 12 16
rect 14 13 19 20
rect 21 17 32 20
rect 21 15 27 17
rect 29 15 32 17
rect 21 13 32 15
rect 34 13 39 20
rect 41 18 48 20
rect 41 16 44 18
rect 46 16 48 18
rect 41 13 48 16
<< pdif >>
rect 23 54 30 55
rect 2 52 9 54
rect 2 50 4 52
rect 6 50 9 52
rect 2 46 9 50
rect 11 50 19 54
rect 11 48 14 50
rect 16 48 19 50
rect 11 46 19 48
rect 21 52 30 54
rect 21 50 25 52
rect 27 50 30 52
rect 21 46 30 50
rect 32 50 40 55
rect 32 48 35 50
rect 37 48 40 50
rect 32 46 40 48
rect 42 52 50 55
rect 42 50 46 52
rect 48 50 50 52
rect 42 46 50 50
<< alu1 >>
rect -2 67 58 72
rect -2 65 5 67
rect 7 65 13 67
rect 15 65 58 67
rect -2 64 58 65
rect 10 50 17 52
rect 10 48 14 50
rect 16 48 17 50
rect 10 46 17 48
rect 10 43 14 46
rect 2 39 14 43
rect 2 19 6 39
rect 41 41 54 43
rect 41 39 43 41
rect 45 39 54 41
rect 41 38 54 39
rect 10 27 14 35
rect 26 27 30 35
rect 10 25 11 27
rect 13 25 22 27
rect 10 23 22 25
rect 2 18 14 19
rect 2 16 7 18
rect 9 16 14 18
rect 2 13 14 16
rect 18 13 22 23
rect 26 25 27 27
rect 29 25 38 27
rect 26 21 38 25
rect 50 21 54 38
rect -2 7 58 8
rect -2 5 49 7
rect 51 5 58 7
rect -2 0 58 5
<< ptie >>
rect 47 7 53 9
rect 47 5 49 7
rect 51 5 53 7
rect 47 3 53 5
<< ntie >>
rect 3 67 17 69
rect 3 65 5 67
rect 7 65 13 67
rect 15 65 17 67
rect 3 63 17 65
<< nmos >>
rect 12 13 14 20
rect 19 13 21 20
rect 32 13 34 20
rect 39 13 41 20
<< pmos >>
rect 9 46 11 54
rect 19 46 21 54
rect 30 46 32 55
rect 40 46 42 55
<< polyct0 >>
rect 21 39 23 41
<< polyct1 >>
rect 11 25 13 27
rect 43 39 45 41
rect 27 25 29 27
<< ndifct0 >>
rect 27 15 29 17
rect 44 16 46 18
<< ndifct1 >>
rect 7 16 9 18
<< ntiect1 >>
rect 5 65 7 67
rect 13 65 15 67
<< ptiect1 >>
rect 49 5 51 7
<< pdifct0 >>
rect 4 50 6 52
rect 25 50 27 52
rect 35 48 37 50
rect 46 50 48 52
<< pdifct1 >>
rect 14 48 16 50
<< alu0 >>
rect 3 52 7 64
rect 24 52 28 64
rect 45 52 49 64
rect 3 50 4 52
rect 6 50 7 52
rect 3 48 7 50
rect 24 50 25 52
rect 27 50 28 52
rect 24 48 28 50
rect 34 50 38 52
rect 34 48 35 50
rect 37 48 38 50
rect 45 50 46 52
rect 48 50 49 52
rect 45 48 49 50
rect 34 42 38 48
rect 19 41 38 42
rect 19 39 21 41
rect 23 39 38 41
rect 19 38 38 39
rect 34 34 38 38
rect 34 30 47 34
rect 43 18 47 30
rect 25 17 31 18
rect 25 15 27 17
rect 29 15 31 17
rect 25 8 31 15
rect 43 16 44 18
rect 46 16 47 18
rect 43 14 47 16
<< labels >>
rlabel alu0 45 24 45 24 6 an
rlabel alu0 28 40 28 40 6 an
rlabel alu1 4 28 4 28 6 z
rlabel alu1 20 20 20 20 6 b
rlabel alu1 12 16 12 16 6 z
rlabel alu1 12 32 12 32 6 b
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 28 28 28 6 a1
rlabel alu1 36 24 36 24 6 a1
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 52 32 52 32 6 a2
rlabel polyct1 44 40 44 40 6 a2
<< end >>
