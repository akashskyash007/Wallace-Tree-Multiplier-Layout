magic
tech scmos
timestamp 1199202546
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 10 62 16 64
rect 10 60 12 62
rect 14 60 16 62
rect 10 58 16 60
rect 10 56 12 58
rect 9 53 12 56
rect 29 55 31 60
rect 9 50 11 53
rect 19 50 21 54
rect 9 30 11 42
rect 19 39 21 42
rect 16 37 23 39
rect 16 35 19 37
rect 21 35 23 37
rect 16 33 23 35
rect 16 30 18 33
rect 29 31 31 45
rect 9 18 11 23
rect 16 18 18 23
rect 28 29 34 31
rect 28 27 30 29
rect 32 27 34 29
rect 28 25 34 27
rect 28 22 30 25
rect 28 11 30 16
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 23 9 26
rect 11 23 16 30
rect 18 23 26 30
rect 20 22 26 23
rect 20 16 28 22
rect 30 20 37 22
rect 30 18 33 20
rect 35 18 37 20
rect 30 16 37 18
rect 20 11 26 16
rect 20 9 22 11
rect 24 9 26 11
rect 20 7 26 9
<< pdif >>
rect 2 71 8 73
rect 2 69 4 71
rect 6 69 8 71
rect 2 58 8 69
rect 21 60 27 62
rect 21 58 23 60
rect 25 58 27 60
rect 2 50 7 58
rect 21 56 27 58
rect 23 55 27 56
rect 23 50 29 55
rect 2 42 9 50
rect 11 46 19 50
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 45 29 50
rect 31 53 38 55
rect 31 51 34 53
rect 36 51 38 53
rect 31 49 38 51
rect 31 45 36 49
rect 21 42 27 45
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 71 42 79
rect -2 69 4 71
rect 6 69 42 71
rect -2 68 42 69
rect 2 62 16 63
rect 2 60 12 62
rect 14 60 16 62
rect 2 57 16 60
rect 2 41 6 57
rect 10 46 23 47
rect 10 44 14 46
rect 16 44 23 46
rect 10 42 23 44
rect 10 31 14 42
rect 2 28 14 31
rect 2 26 4 28
rect 6 26 14 28
rect 2 25 14 26
rect 34 31 38 47
rect 26 29 38 31
rect 26 27 30 29
rect 32 27 38 29
rect 26 25 38 27
rect -2 11 42 12
rect -2 9 22 11
rect 24 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 23 11 30
rect 16 23 18 30
rect 28 16 30 22
<< pmos >>
rect 9 42 11 50
rect 19 42 21 50
rect 29 45 31 55
<< polyct0 >>
rect 19 35 21 37
<< polyct1 >>
rect 12 60 14 62
rect 30 27 32 29
<< ndifct0 >>
rect 33 18 35 20
<< ndifct1 >>
rect 4 26 6 28
rect 22 9 24 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 23 58 25 60
rect 34 51 36 53
<< pdifct1 >>
rect 4 69 6 71
rect 14 44 16 46
<< alu0 >>
rect 21 60 27 68
rect 21 58 23 60
rect 25 58 27 60
rect 21 57 27 58
rect 26 53 38 54
rect 26 51 34 53
rect 36 51 38 53
rect 26 50 38 51
rect 26 39 30 50
rect 18 37 30 39
rect 18 35 19 37
rect 21 35 30 37
rect 18 21 22 35
rect 18 20 37 21
rect 18 18 33 20
rect 35 18 37 20
rect 18 17 37 18
<< labels >>
rlabel alu0 20 28 20 28 6 an
rlabel alu0 27 19 27 19 6 an
rlabel alu0 32 52 32 52 6 an
rlabel alu1 4 28 4 28 6 z
rlabel alu1 4 52 4 52 6 b
rlabel alu1 12 36 12 36 6 z
rlabel alu1 12 60 12 60 6 b
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 28 28 28 6 a
rlabel alu1 20 44 20 44 6 z
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 36 36 36 6 a
<< end >>
