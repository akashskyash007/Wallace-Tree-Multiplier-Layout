magic
tech scmos
timestamp 1199470035
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -5 48 55 105
<< pwell >>
rect -5 -5 55 48
<< poly >>
rect 15 94 17 98
rect 23 94 25 98
rect 37 77 39 82
rect 15 43 17 55
rect 23 52 25 55
rect 37 52 39 55
rect 23 49 27 52
rect 13 41 21 43
rect 13 39 17 41
rect 19 39 21 41
rect 13 37 21 39
rect 25 42 27 49
rect 32 50 39 52
rect 32 48 34 50
rect 36 48 39 50
rect 32 46 39 48
rect 25 40 32 42
rect 25 38 28 40
rect 30 38 32 40
rect 13 28 15 37
rect 25 36 32 38
rect 25 28 27 36
rect 37 28 39 46
rect 13 12 15 17
rect 25 12 27 17
rect 37 12 39 17
<< ndif >>
rect 4 17 13 28
rect 15 21 25 28
rect 15 19 19 21
rect 21 19 25 21
rect 15 17 25 19
rect 27 21 37 28
rect 27 19 31 21
rect 33 19 37 21
rect 27 17 37 19
rect 39 26 47 28
rect 39 24 43 26
rect 45 24 47 26
rect 39 22 47 24
rect 39 17 44 22
rect 4 11 11 17
rect 4 9 7 11
rect 9 9 11 11
rect 4 7 11 9
<< pdif >>
rect 10 69 15 94
rect 7 67 15 69
rect 7 65 9 67
rect 11 65 15 67
rect 7 59 15 65
rect 7 57 9 59
rect 11 57 15 59
rect 7 55 15 57
rect 17 55 23 94
rect 25 91 35 94
rect 25 89 29 91
rect 31 89 35 91
rect 25 81 35 89
rect 25 79 29 81
rect 31 79 35 81
rect 25 77 35 79
rect 25 71 37 77
rect 25 69 29 71
rect 31 69 37 71
rect 25 55 37 69
rect 39 69 44 77
rect 39 67 47 69
rect 39 65 43 67
rect 45 65 47 67
rect 39 59 47 65
rect 39 57 43 59
rect 45 57 47 59
rect 39 55 47 57
<< alu1 >>
rect -2 95 52 100
rect -2 93 43 95
rect 45 93 52 95
rect -2 91 52 93
rect -2 89 29 91
rect 31 89 52 91
rect -2 88 52 89
rect 28 81 32 88
rect 28 79 29 81
rect 31 79 32 81
rect 8 67 12 73
rect 8 65 9 67
rect 11 65 12 67
rect 8 59 12 65
rect 8 57 9 59
rect 11 57 12 59
rect 18 63 22 73
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 67 32 69
rect 42 67 46 69
rect 42 65 43 67
rect 45 65 46 67
rect 18 57 32 63
rect 8 23 12 57
rect 18 44 22 53
rect 28 51 32 57
rect 42 59 46 65
rect 42 57 43 59
rect 45 57 46 59
rect 28 50 38 51
rect 28 48 34 50
rect 36 48 38 50
rect 28 47 38 48
rect 16 41 22 44
rect 42 41 46 57
rect 16 39 17 41
rect 19 39 22 41
rect 16 38 22 39
rect 18 32 22 38
rect 26 40 46 41
rect 26 38 28 40
rect 30 38 46 40
rect 26 37 46 38
rect 18 27 33 32
rect 42 26 46 37
rect 42 24 43 26
rect 45 24 46 26
rect 8 21 22 23
rect 8 19 19 21
rect 21 19 22 21
rect 8 17 22 19
rect 30 21 34 23
rect 42 22 46 24
rect 30 19 31 21
rect 33 19 34 21
rect 30 12 34 19
rect -2 11 52 12
rect -2 9 7 11
rect 9 9 52 11
rect -2 7 52 9
rect -2 5 19 7
rect 21 5 29 7
rect 31 5 52 7
rect -2 0 52 5
<< ptie >>
rect 17 7 33 9
rect 17 5 19 7
rect 21 5 29 7
rect 31 5 33 7
rect 17 3 33 5
<< ntie >>
rect 41 95 47 97
rect 41 93 43 95
rect 45 93 47 95
rect 41 91 47 93
<< nmos >>
rect 13 17 15 28
rect 25 17 27 28
rect 37 17 39 28
<< pmos >>
rect 15 55 17 94
rect 23 55 25 94
rect 37 55 39 77
<< polyct1 >>
rect 17 39 19 41
rect 34 48 36 50
rect 28 38 30 40
<< ndifct1 >>
rect 19 19 21 21
rect 31 19 33 21
rect 43 24 45 26
rect 7 9 9 11
<< ntiect1 >>
rect 43 93 45 95
<< ptiect1 >>
rect 19 5 21 7
rect 29 5 31 7
<< pdifct1 >>
rect 9 65 11 67
rect 9 57 11 59
rect 29 89 31 91
rect 29 79 31 81
rect 29 69 31 71
rect 43 65 45 67
rect 43 57 45 59
<< labels >>
rlabel polyct1 29 39 29 39 6 an
rlabel ndifct1 44 25 44 25 6 an
rlabel pdifct1 44 66 44 66 6 an
rlabel ndifct1 20 20 20 20 6 z
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 65 20 65 6 a
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 30 30 30 6 b
rlabel alu1 30 55 30 55 6 a
rlabel alu1 25 94 25 94 6 vdd
<< end >>
