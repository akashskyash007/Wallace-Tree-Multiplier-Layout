magic
tech scmos
timestamp 1199202094
<< ab >>
rect 0 0 112 72
<< nwell >>
rect -5 32 117 77
<< pwell >>
rect -5 -5 117 32
<< poly >>
rect 25 68 110 70
rect 15 59 17 64
rect 25 60 27 68
rect 56 65 58 68
rect 35 60 37 64
rect 77 60 79 64
rect 87 60 89 68
rect 97 60 99 64
rect 56 40 58 43
rect 56 38 61 40
rect 15 35 17 38
rect 2 33 17 35
rect 25 35 27 38
rect 25 33 30 35
rect 2 31 4 33
rect 6 31 17 33
rect 2 29 17 31
rect 12 22 14 29
rect 28 27 30 33
rect 35 34 37 38
rect 59 36 61 38
rect 59 34 65 36
rect 77 35 79 38
rect 35 32 55 34
rect 43 30 51 32
rect 53 30 55 32
rect 43 28 55 30
rect 59 32 61 34
rect 63 32 65 34
rect 59 30 65 32
rect 73 33 79 35
rect 87 33 89 38
rect 97 35 99 38
rect 94 33 99 35
rect 73 31 75 33
rect 77 31 79 33
rect 22 22 24 27
rect 28 25 34 27
rect 32 22 34 25
rect 12 7 14 12
rect 22 4 24 12
rect 32 8 34 12
rect 43 4 45 28
rect 59 26 61 30
rect 73 29 79 31
rect 94 29 96 33
rect 108 29 110 68
rect 73 27 83 29
rect 81 24 83 27
rect 91 27 96 29
rect 101 27 110 29
rect 91 24 93 27
rect 101 24 103 27
rect 59 11 61 16
rect 81 9 83 14
rect 91 4 93 14
rect 101 9 103 14
rect 22 2 93 4
<< ndif >>
rect 3 16 12 22
rect 3 14 6 16
rect 8 14 12 16
rect 3 12 12 14
rect 14 20 22 22
rect 14 18 17 20
rect 19 18 22 20
rect 14 12 22 18
rect 24 20 32 22
rect 24 18 27 20
rect 29 18 32 20
rect 24 12 32 18
rect 34 19 39 22
rect 34 17 41 19
rect 34 15 37 17
rect 39 15 41 17
rect 34 12 41 15
rect 52 24 59 26
rect 52 22 54 24
rect 56 22 59 24
rect 52 20 59 22
rect 54 16 59 20
rect 61 24 66 26
rect 61 18 81 24
rect 61 16 72 18
rect 74 16 81 18
rect 63 14 81 16
rect 83 22 91 24
rect 83 20 86 22
rect 88 20 91 22
rect 83 14 91 20
rect 93 18 101 24
rect 93 16 96 18
rect 98 16 101 18
rect 93 14 101 16
rect 103 22 110 24
rect 103 20 106 22
rect 108 20 110 22
rect 103 18 110 20
rect 103 14 108 18
<< pdif >>
rect 20 59 25 60
rect 7 57 15 59
rect 7 55 10 57
rect 12 55 15 57
rect 7 50 15 55
rect 7 48 10 50
rect 12 48 15 50
rect 7 38 15 48
rect 17 49 25 59
rect 17 47 20 49
rect 22 47 25 49
rect 17 42 25 47
rect 17 40 20 42
rect 22 40 25 42
rect 17 38 25 40
rect 27 49 35 60
rect 27 47 30 49
rect 32 47 35 49
rect 27 42 35 47
rect 27 40 30 42
rect 32 40 35 42
rect 27 38 35 40
rect 37 51 42 60
rect 37 49 44 51
rect 51 49 56 65
rect 37 47 40 49
rect 42 47 44 49
rect 37 42 44 47
rect 49 47 56 49
rect 49 45 51 47
rect 53 45 56 47
rect 49 43 56 45
rect 58 63 75 65
rect 58 61 64 63
rect 66 61 75 63
rect 58 60 75 61
rect 58 43 77 60
rect 37 40 40 42
rect 42 40 44 42
rect 37 38 44 40
rect 67 38 77 43
rect 79 49 87 60
rect 79 47 82 49
rect 84 47 87 49
rect 79 42 87 47
rect 79 40 82 42
rect 84 40 87 42
rect 79 38 87 40
rect 89 49 97 60
rect 89 47 92 49
rect 94 47 97 49
rect 89 42 97 47
rect 89 40 92 42
rect 94 40 97 42
rect 89 38 97 40
rect 99 58 106 60
rect 99 56 102 58
rect 104 56 106 58
rect 99 51 106 56
rect 99 49 102 51
rect 104 49 106 51
rect 99 47 106 49
rect 99 38 104 47
<< alu1 >>
rect -2 67 114 72
rect -2 65 5 67
rect 7 65 114 67
rect -2 64 114 65
rect 2 37 14 43
rect 2 33 7 37
rect 2 31 4 33
rect 6 31 7 33
rect 2 21 7 31
rect 26 49 33 51
rect 26 47 30 49
rect 32 47 33 49
rect 26 42 33 47
rect 26 40 30 42
rect 32 40 33 42
rect 26 38 33 40
rect 26 27 30 38
rect 65 46 78 50
rect 26 21 38 27
rect 26 20 30 21
rect 26 18 27 20
rect 29 18 30 20
rect 57 35 63 42
rect 57 34 70 35
rect 57 32 61 34
rect 63 32 70 34
rect 57 29 70 32
rect 74 33 78 46
rect 74 31 75 33
rect 77 31 78 33
rect 74 29 78 31
rect 90 49 95 51
rect 90 47 92 49
rect 94 47 95 49
rect 90 42 95 47
rect 90 40 92 42
rect 94 40 95 42
rect 90 35 95 40
rect 90 29 102 35
rect 26 13 30 18
rect 98 19 102 29
rect 94 18 102 19
rect 94 16 96 18
rect 98 16 102 18
rect 94 13 102 16
rect -2 0 114 8
<< ptie >>
rect 47 10 53 12
rect 47 8 49 10
rect 51 8 53 10
rect 47 6 53 8
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 12 12 14 22
rect 22 12 24 22
rect 32 12 34 22
rect 59 16 61 26
rect 81 14 83 24
rect 91 14 93 24
rect 101 14 103 24
<< pmos >>
rect 15 38 17 59
rect 25 38 27 60
rect 35 38 37 60
rect 56 43 58 65
rect 77 38 79 60
rect 87 38 89 60
rect 97 38 99 60
<< polyct0 >>
rect 51 30 53 32
<< polyct1 >>
rect 4 31 6 33
rect 61 32 63 34
rect 75 31 77 33
<< ndifct0 >>
rect 6 14 8 16
rect 17 18 19 20
rect 37 15 39 17
rect 54 22 56 24
rect 72 16 74 18
rect 86 20 88 22
rect 106 20 108 22
<< ndifct1 >>
rect 27 18 29 20
rect 96 16 98 18
<< ntiect1 >>
rect 5 65 7 67
<< ptiect0 >>
rect 49 8 51 10
<< pdifct0 >>
rect 10 55 12 57
rect 10 48 12 50
rect 20 47 22 49
rect 20 40 22 42
rect 40 47 42 49
rect 51 45 53 47
rect 64 61 66 63
rect 40 40 42 42
rect 82 47 84 49
rect 82 40 84 42
rect 102 56 104 58
rect 102 49 104 51
<< pdifct1 >>
rect 30 47 32 49
rect 30 40 32 42
rect 92 47 94 49
rect 92 40 94 42
<< alu0 >>
rect 9 57 13 64
rect 62 63 68 64
rect 62 61 64 63
rect 66 61 68 63
rect 62 60 68 61
rect 9 55 10 57
rect 12 55 13 57
rect 9 50 13 55
rect 9 48 10 50
rect 12 48 13 50
rect 9 46 13 48
rect 19 57 52 59
rect 72 58 106 59
rect 72 57 102 58
rect 19 56 102 57
rect 104 56 106 58
rect 19 55 106 56
rect 19 49 23 55
rect 48 53 76 55
rect 100 52 106 55
rect 100 51 109 52
rect 19 47 20 49
rect 22 47 23 49
rect 19 42 23 47
rect 19 40 20 42
rect 22 40 23 42
rect 19 34 23 40
rect 16 30 23 34
rect 39 49 43 51
rect 39 47 40 49
rect 42 47 43 49
rect 39 42 43 47
rect 39 40 40 42
rect 42 40 43 42
rect 16 20 20 30
rect 16 18 17 20
rect 19 18 20 20
rect 4 16 10 17
rect 16 16 20 18
rect 39 35 43 40
rect 50 47 54 49
rect 50 45 51 47
rect 53 45 54 47
rect 39 31 46 35
rect 42 18 46 31
rect 50 32 54 45
rect 50 30 51 32
rect 53 30 54 32
rect 50 25 54 30
rect 81 49 85 51
rect 81 47 82 49
rect 84 47 85 49
rect 81 42 85 47
rect 81 40 82 42
rect 84 40 85 42
rect 81 26 85 40
rect 100 49 102 51
rect 104 49 109 51
rect 100 48 109 49
rect 50 24 58 25
rect 50 22 54 24
rect 56 22 58 24
rect 50 21 58 22
rect 62 22 89 26
rect 62 18 66 22
rect 85 20 86 22
rect 88 20 89 22
rect 4 14 6 16
rect 8 14 10 16
rect 4 8 10 14
rect 35 17 66 18
rect 35 15 37 17
rect 39 15 66 17
rect 35 14 66 15
rect 70 18 76 19
rect 85 18 89 20
rect 105 22 109 48
rect 105 20 106 22
rect 108 20 109 22
rect 105 18 109 20
rect 70 16 72 18
rect 74 16 76 18
rect 47 10 53 11
rect 47 8 49 10
rect 51 8 53 10
rect 70 8 76 16
<< labels >>
rlabel alu0 18 25 18 25 6 a0n
rlabel alu0 21 44 21 44 6 a0n
rlabel alu0 52 35 52 35 6 sn
rlabel pdifct0 41 41 41 41 6 a1n
rlabel alu0 50 16 50 16 6 a1n
rlabel alu0 75 24 75 24 6 a1n
rlabel alu0 83 36 83 36 6 a1n
rlabel alu0 107 35 107 35 6 a0n
rlabel alu0 89 57 89 57 6 a0n
rlabel alu1 4 32 4 32 6 a0
rlabel alu1 12 40 12 40 6 a0
rlabel alu1 28 32 28 32 6 z0
rlabel alu1 36 24 36 24 6 z0
rlabel alu1 56 4 56 4 6 vss
rlabel alu1 68 32 68 32 6 s
rlabel alu1 76 36 76 36 6 a1
rlabel alu1 60 36 60 36 6 s
rlabel alu1 68 48 68 48 6 a1
rlabel alu1 56 68 56 68 6 vdd
rlabel alu1 100 24 100 24 6 z1
rlabel alu1 92 40 92 40 6 z1
<< end >>
