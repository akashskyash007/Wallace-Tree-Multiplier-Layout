magic
tech scmos
timestamp 1199201783
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 37 70 39 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 2 37 11 39
rect 2 35 4 37
rect 6 35 11 37
rect 2 33 11 35
rect 9 30 11 33
rect 16 37 23 39
rect 16 35 19 37
rect 21 35 23 37
rect 16 33 23 35
rect 27 37 33 39
rect 27 35 29 37
rect 31 35 33 37
rect 27 33 33 35
rect 16 30 18 33
rect 27 28 29 33
rect 37 31 39 42
rect 37 29 43 31
rect 37 28 39 29
rect 26 25 29 28
rect 36 27 39 28
rect 41 27 43 29
rect 36 25 43 27
rect 26 22 28 25
rect 36 22 38 25
rect 9 16 11 21
rect 16 17 18 21
rect 26 11 28 16
rect 36 11 38 16
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 21 9 24
rect 11 21 16 30
rect 18 22 24 30
rect 18 21 26 22
rect 20 16 26 21
rect 28 20 36 22
rect 28 18 31 20
rect 33 18 36 20
rect 28 16 36 18
rect 38 16 46 22
rect 20 15 24 16
rect 18 13 24 15
rect 18 11 20 13
rect 22 11 24 13
rect 40 11 46 16
rect 18 9 24 11
rect 40 9 42 11
rect 44 9 46 11
rect 40 7 46 9
<< pdif >>
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 42 9 58
rect 11 46 19 70
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 62 29 70
rect 21 60 24 62
rect 26 60 29 62
rect 21 42 29 60
rect 31 42 37 70
rect 39 68 46 70
rect 39 66 42 68
rect 44 66 46 68
rect 39 61 46 66
rect 39 59 42 61
rect 44 59 46 61
rect 39 42 46 59
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 2 50 15 55
rect 2 37 6 50
rect 25 46 31 54
rect 21 42 31 46
rect 21 39 25 42
rect 2 35 4 37
rect 2 33 6 35
rect 10 22 14 39
rect 18 37 25 39
rect 18 35 19 37
rect 21 35 25 37
rect 18 33 25 35
rect 42 38 46 55
rect 33 34 46 38
rect 33 29 46 30
rect 33 27 39 29
rect 41 27 46 29
rect 33 26 46 27
rect 10 20 36 22
rect 10 18 31 20
rect 33 18 36 20
rect 10 17 36 18
rect 42 17 46 26
rect -2 11 20 12
rect 22 11 50 12
rect -2 9 42 11
rect 44 9 50 11
rect -2 1 50 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 9 21 11 30
rect 16 21 18 30
rect 26 16 28 22
rect 36 16 38 22
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 37 42 39 70
<< polyct0 >>
rect 29 35 31 37
<< polyct1 >>
rect 4 35 6 37
rect 19 35 21 37
rect 39 27 41 29
<< ndifct0 >>
rect 4 26 6 28
rect 20 12 22 13
<< ndifct1 >>
rect 31 18 33 20
rect 20 11 22 12
rect 42 9 44 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 4 60 6 62
rect 14 44 16 46
rect 24 60 26 62
rect 42 66 44 68
rect 42 59 44 61
<< alu0 >>
rect 40 66 42 68
rect 44 66 46 68
rect 2 62 28 63
rect 2 60 4 62
rect 6 60 24 62
rect 26 60 28 62
rect 2 59 28 60
rect 40 61 46 66
rect 40 59 42 61
rect 44 59 46 61
rect 40 58 46 59
rect 11 46 18 47
rect 11 44 14 46
rect 16 44 18 46
rect 11 43 18 44
rect 11 39 15 43
rect 6 33 7 39
rect 2 28 10 29
rect 2 26 4 28
rect 6 26 10 28
rect 2 25 10 26
rect 14 35 15 39
rect 28 38 42 39
rect 28 37 33 38
rect 28 35 29 37
rect 31 35 33 37
rect 28 34 33 35
rect 28 33 37 34
rect 18 13 24 14
rect 18 12 20 13
rect 22 12 24 13
<< labels >>
rlabel alu0 15 61 15 61 6 n2
rlabel alu1 4 44 4 44 6 c2
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 28 12 28 6 z
rlabel polyct1 20 36 20 36 6 c1
rlabel alu1 12 52 12 52 6 c2
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 48 28 48 6 c1
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 44 20 44 20 6 a
rlabel alu1 36 36 36 36 6 b
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 48 44 48 6 b
<< end >>
