magic
tech scmos
timestamp 1199543826
<< ab >>
rect 0 0 180 100
<< nwell >>
rect -2 48 182 104
<< pwell >>
rect -2 -4 182 48
<< poly >>
rect 47 95 49 98
rect 59 95 61 98
rect 95 95 97 98
rect 107 95 109 98
rect 119 95 121 98
rect 131 95 133 98
rect 143 95 145 98
rect 155 95 157 98
rect 167 95 169 98
rect 11 85 13 88
rect 23 85 25 88
rect 71 85 73 88
rect 83 85 85 88
rect 47 73 49 75
rect 47 71 53 73
rect 47 69 49 71
rect 51 69 53 71
rect 47 67 53 69
rect 11 63 13 65
rect 11 61 19 63
rect 11 59 15 61
rect 17 59 19 61
rect 11 57 19 59
rect 3 51 9 53
rect 23 51 25 65
rect 59 63 61 75
rect 95 73 97 75
rect 95 71 103 73
rect 95 69 99 71
rect 101 69 103 71
rect 95 67 103 69
rect 71 63 73 65
rect 37 61 43 63
rect 57 61 63 63
rect 37 59 39 61
rect 41 59 59 61
rect 61 59 63 61
rect 37 57 43 59
rect 57 57 63 59
rect 67 61 73 63
rect 67 59 69 61
rect 71 59 73 61
rect 67 57 73 59
rect 67 51 73 53
rect 83 51 85 65
rect 107 63 109 75
rect 101 61 109 63
rect 101 59 103 61
rect 105 59 109 61
rect 101 57 109 59
rect 119 51 121 75
rect 131 73 133 75
rect 125 71 133 73
rect 125 69 127 71
rect 129 69 133 71
rect 125 67 133 69
rect 143 53 145 75
rect 143 51 151 53
rect 3 49 5 51
rect 7 49 69 51
rect 71 49 133 51
rect 3 47 9 49
rect 11 31 19 33
rect 11 29 15 31
rect 17 29 19 31
rect 11 27 19 29
rect 11 25 13 27
rect 23 25 25 49
rect 67 47 73 49
rect 29 41 35 43
rect 77 41 85 43
rect 119 41 127 43
rect 29 39 31 41
rect 33 39 79 41
rect 81 39 123 41
rect 125 39 127 41
rect 29 37 35 39
rect 77 37 85 39
rect 47 31 53 33
rect 47 29 49 31
rect 51 29 53 31
rect 47 27 53 29
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 57 27 63 29
rect 67 31 73 33
rect 67 29 69 31
rect 71 29 73 31
rect 67 27 73 29
rect 47 25 49 27
rect 59 25 61 27
rect 71 25 73 27
rect 83 25 85 37
rect 119 37 127 39
rect 101 31 109 33
rect 101 29 103 31
rect 105 29 109 31
rect 101 27 109 29
rect 95 21 103 23
rect 95 19 99 21
rect 101 19 103 21
rect 95 17 103 19
rect 95 15 97 17
rect 107 15 109 27
rect 119 25 121 37
rect 131 25 133 49
rect 143 49 147 51
rect 149 49 151 51
rect 143 47 151 49
rect 155 43 157 55
rect 167 43 169 55
rect 145 41 169 43
rect 145 39 147 41
rect 149 39 169 41
rect 145 37 169 39
rect 143 31 151 33
rect 143 29 147 31
rect 149 29 151 31
rect 143 27 151 29
rect 143 25 145 27
rect 155 25 157 37
rect 167 25 169 37
rect 11 12 13 15
rect 23 12 25 15
rect 47 12 49 15
rect 59 12 61 15
rect 71 12 73 15
rect 83 12 85 15
rect 119 12 121 15
rect 131 12 133 15
rect 143 12 145 15
rect 95 2 97 5
rect 107 2 109 5
rect 155 2 157 5
rect 167 2 169 5
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 25 21 33 25
rect 25 19 29 21
rect 31 19 33 21
rect 25 15 33 19
rect 39 21 47 25
rect 39 19 41 21
rect 43 19 47 21
rect 39 15 47 19
rect 49 15 59 25
rect 61 15 71 25
rect 73 21 83 25
rect 73 19 77 21
rect 79 19 83 21
rect 73 15 83 19
rect 85 15 93 25
rect 111 21 119 25
rect 111 19 113 21
rect 115 19 119 21
rect 111 15 119 19
rect 121 21 131 25
rect 121 19 125 21
rect 127 19 131 21
rect 121 15 131 19
rect 133 15 143 25
rect 145 21 155 25
rect 145 19 149 21
rect 151 19 155 21
rect 145 15 155 19
rect 15 11 21 15
rect 15 9 17 11
rect 19 9 21 11
rect 51 11 57 15
rect 51 9 53 11
rect 55 9 57 11
rect 15 7 21 9
rect 51 7 57 9
rect 87 5 95 15
rect 97 11 107 15
rect 97 9 101 11
rect 103 9 107 11
rect 97 5 107 9
rect 109 5 117 15
rect 147 11 155 15
rect 147 9 149 11
rect 151 9 155 11
rect 147 5 155 9
rect 157 21 167 25
rect 157 19 161 21
rect 163 19 167 21
rect 157 5 167 19
rect 169 21 177 25
rect 169 19 173 21
rect 175 19 177 21
rect 169 11 177 19
rect 169 9 173 11
rect 175 9 177 11
rect 169 5 177 9
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 65 23 85
rect 25 71 33 85
rect 39 81 47 95
rect 39 79 41 81
rect 43 79 47 81
rect 39 75 47 79
rect 49 91 59 95
rect 49 89 53 91
rect 55 89 59 91
rect 49 75 59 89
rect 61 85 69 95
rect 87 85 95 95
rect 61 75 71 85
rect 25 69 29 71
rect 31 69 33 71
rect 25 65 33 69
rect 63 65 71 75
rect 73 71 83 85
rect 73 69 77 71
rect 79 69 83 71
rect 73 65 83 69
rect 85 75 95 85
rect 97 91 107 95
rect 97 89 101 91
rect 103 89 107 91
rect 97 75 107 89
rect 109 81 119 95
rect 109 79 113 81
rect 115 79 119 81
rect 109 75 119 79
rect 121 81 131 95
rect 121 79 125 81
rect 127 79 131 81
rect 121 75 131 79
rect 133 75 143 95
rect 145 91 155 95
rect 145 89 149 91
rect 151 89 155 91
rect 145 81 155 89
rect 145 79 149 81
rect 151 79 155 81
rect 145 75 155 79
rect 85 65 93 75
rect 147 71 155 75
rect 147 69 149 71
rect 151 69 155 71
rect 147 61 155 69
rect 147 59 149 61
rect 151 59 155 61
rect 147 55 155 59
rect 157 81 167 95
rect 157 79 161 81
rect 163 79 167 81
rect 157 71 167 79
rect 157 69 161 71
rect 163 69 167 71
rect 157 61 167 69
rect 157 59 161 61
rect 163 59 167 61
rect 157 55 167 59
rect 169 91 177 95
rect 169 89 173 91
rect 175 89 177 91
rect 169 81 177 89
rect 169 79 173 81
rect 175 79 177 81
rect 169 71 177 79
rect 169 69 173 71
rect 175 69 177 71
rect 169 61 177 69
rect 169 59 173 61
rect 175 59 177 61
rect 169 55 177 59
<< alu1 >>
rect -2 91 182 100
rect -2 89 17 91
rect 19 89 53 91
rect 55 89 101 91
rect 103 89 149 91
rect 151 89 173 91
rect 175 89 182 91
rect -2 88 182 89
rect 4 81 8 82
rect 4 79 5 81
rect 7 79 8 81
rect 4 78 8 79
rect 5 72 7 78
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 52 7 68
rect 18 62 22 82
rect 40 81 44 82
rect 58 81 62 82
rect 40 79 41 81
rect 43 79 44 81
rect 40 78 44 79
rect 50 79 62 81
rect 28 71 32 72
rect 28 69 29 71
rect 31 69 32 71
rect 28 68 32 69
rect 14 61 22 62
rect 14 59 15 61
rect 17 59 22 61
rect 14 58 22 59
rect 4 51 8 52
rect 4 49 5 51
rect 7 49 8 51
rect 4 48 8 49
rect 5 22 7 48
rect 18 32 22 58
rect 14 31 22 32
rect 14 29 15 31
rect 17 29 22 31
rect 14 28 22 29
rect 4 21 8 22
rect 4 19 5 21
rect 7 19 8 21
rect 4 18 8 19
rect 18 18 22 28
rect 29 42 31 68
rect 40 62 42 78
rect 50 72 52 79
rect 58 78 62 79
rect 112 81 116 82
rect 112 79 113 81
rect 115 79 116 81
rect 112 78 116 79
rect 124 81 128 82
rect 148 81 152 88
rect 124 79 125 81
rect 127 79 139 81
rect 124 78 128 79
rect 38 61 42 62
rect 38 59 39 61
rect 41 59 42 61
rect 38 58 42 59
rect 29 41 34 42
rect 29 39 31 41
rect 33 39 34 41
rect 29 38 34 39
rect 29 22 31 38
rect 40 22 42 58
rect 48 71 52 72
rect 48 69 49 71
rect 51 69 52 71
rect 48 31 52 69
rect 76 71 80 72
rect 98 71 102 72
rect 113 71 115 78
rect 126 71 130 72
rect 76 69 77 71
rect 79 69 91 71
rect 76 68 80 69
rect 58 61 62 62
rect 58 59 59 61
rect 61 59 62 61
rect 58 58 62 59
rect 68 61 72 62
rect 89 61 91 69
rect 98 69 99 71
rect 101 69 115 71
rect 98 68 102 69
rect 102 61 106 62
rect 68 59 69 61
rect 71 59 81 61
rect 68 58 72 59
rect 59 32 61 58
rect 68 51 72 52
rect 68 49 69 51
rect 71 49 72 51
rect 68 48 72 49
rect 69 32 71 48
rect 79 42 81 59
rect 89 59 103 61
rect 105 59 106 61
rect 78 41 82 42
rect 78 39 79 41
rect 81 39 82 41
rect 78 38 82 39
rect 48 29 49 31
rect 51 29 52 31
rect 48 28 52 29
rect 58 31 62 32
rect 58 29 59 31
rect 61 29 62 31
rect 58 28 62 29
rect 68 31 72 32
rect 68 29 69 31
rect 71 29 72 31
rect 68 28 72 29
rect 89 31 91 59
rect 102 58 106 59
rect 102 31 106 32
rect 89 29 103 31
rect 105 29 106 31
rect 28 21 32 22
rect 28 19 29 21
rect 31 19 32 21
rect 28 18 32 19
rect 40 21 44 22
rect 40 19 41 21
rect 43 19 44 21
rect 50 21 52 28
rect 58 21 62 22
rect 50 19 62 21
rect 40 18 44 19
rect 58 18 62 19
rect 76 21 80 22
rect 89 21 91 29
rect 102 28 106 29
rect 113 22 115 69
rect 125 69 127 71
rect 129 69 130 71
rect 125 68 130 69
rect 125 42 127 68
rect 122 41 127 42
rect 122 39 123 41
rect 125 39 127 41
rect 137 41 139 79
rect 148 79 149 81
rect 151 79 152 81
rect 148 71 152 79
rect 148 69 149 71
rect 151 69 152 71
rect 148 61 152 69
rect 148 59 149 61
rect 151 59 152 61
rect 148 58 152 59
rect 158 81 164 82
rect 158 79 161 81
rect 163 79 164 81
rect 158 78 164 79
rect 172 81 176 88
rect 172 79 173 81
rect 175 79 176 81
rect 158 72 162 78
rect 158 71 164 72
rect 158 69 161 71
rect 163 69 164 71
rect 158 68 164 69
rect 172 71 176 79
rect 172 69 173 71
rect 175 69 176 71
rect 158 62 162 68
rect 158 61 164 62
rect 158 59 161 61
rect 163 59 164 61
rect 158 58 164 59
rect 172 61 176 69
rect 172 59 173 61
rect 175 59 176 61
rect 172 58 176 59
rect 146 51 150 52
rect 158 51 162 58
rect 146 49 147 51
rect 149 49 163 51
rect 146 48 150 49
rect 146 41 150 42
rect 137 39 147 41
rect 149 39 150 41
rect 122 38 126 39
rect 76 19 77 21
rect 79 19 91 21
rect 98 21 102 22
rect 112 21 116 22
rect 98 19 99 21
rect 101 19 113 21
rect 115 19 116 21
rect 76 18 80 19
rect 98 18 102 19
rect 112 18 116 19
rect 124 21 128 22
rect 137 21 139 39
rect 146 38 150 39
rect 146 31 150 32
rect 158 31 162 49
rect 146 29 147 31
rect 149 29 163 31
rect 146 28 150 29
rect 158 22 162 29
rect 124 19 125 21
rect 127 19 139 21
rect 148 21 152 22
rect 148 19 149 21
rect 151 19 152 21
rect 124 18 128 19
rect 148 12 152 19
rect 158 21 164 22
rect 158 19 161 21
rect 163 19 164 21
rect 158 18 164 19
rect 172 21 176 22
rect 172 19 173 21
rect 175 19 176 21
rect 172 12 176 19
rect -2 11 182 12
rect -2 9 17 11
rect 19 9 53 11
rect 55 9 101 11
rect 103 9 149 11
rect 151 9 173 11
rect 175 9 182 11
rect -2 7 182 9
rect -2 5 29 7
rect 31 5 41 7
rect 43 5 65 7
rect 67 5 77 7
rect 79 5 125 7
rect 127 5 137 7
rect 139 5 182 7
rect -2 0 182 5
<< ptie >>
rect 27 7 45 9
rect 63 7 81 9
rect 27 5 29 7
rect 31 5 41 7
rect 43 5 45 7
rect 27 3 45 5
rect 63 5 65 7
rect 67 5 77 7
rect 79 5 81 7
rect 123 7 141 9
rect 123 5 125 7
rect 127 5 137 7
rect 139 5 141 7
rect 63 3 81 5
rect 123 3 141 5
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 47 15 49 25
rect 59 15 61 25
rect 71 15 73 25
rect 83 15 85 25
rect 119 15 121 25
rect 131 15 133 25
rect 143 15 145 25
rect 95 5 97 15
rect 107 5 109 15
rect 155 5 157 25
rect 167 5 169 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 47 75 49 95
rect 59 75 61 95
rect 71 65 73 85
rect 83 65 85 85
rect 95 75 97 95
rect 107 75 109 95
rect 119 75 121 95
rect 131 75 133 95
rect 143 75 145 95
rect 155 55 157 95
rect 167 55 169 95
<< polyct1 >>
rect 49 69 51 71
rect 15 59 17 61
rect 99 69 101 71
rect 39 59 41 61
rect 59 59 61 61
rect 69 59 71 61
rect 103 59 105 61
rect 127 69 129 71
rect 5 49 7 51
rect 69 49 71 51
rect 15 29 17 31
rect 31 39 33 41
rect 79 39 81 41
rect 123 39 125 41
rect 49 29 51 31
rect 59 29 61 31
rect 69 29 71 31
rect 103 29 105 31
rect 99 19 101 21
rect 147 49 149 51
rect 147 39 149 41
rect 147 29 149 31
<< ndifct1 >>
rect 5 19 7 21
rect 29 19 31 21
rect 41 19 43 21
rect 77 19 79 21
rect 113 19 115 21
rect 125 19 127 21
rect 149 19 151 21
rect 17 9 19 11
rect 53 9 55 11
rect 101 9 103 11
rect 149 9 151 11
rect 161 19 163 21
rect 173 19 175 21
rect 173 9 175 11
<< ptiect1 >>
rect 29 5 31 7
rect 41 5 43 7
rect 65 5 67 7
rect 77 5 79 7
rect 125 5 127 7
rect 137 5 139 7
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 5 69 7 71
rect 41 79 43 81
rect 53 89 55 91
rect 29 69 31 71
rect 77 69 79 71
rect 101 89 103 91
rect 113 79 115 81
rect 125 79 127 81
rect 149 89 151 91
rect 149 79 151 81
rect 149 69 151 71
rect 149 59 151 61
rect 161 79 163 81
rect 161 69 163 71
rect 161 59 163 61
rect 173 89 175 91
rect 173 79 175 81
rect 173 69 175 71
rect 173 59 175 61
<< labels >>
rlabel alu1 20 50 20 50 6 ck
rlabel alu1 60 20 60 20 6 i
rlabel alu1 50 50 50 50 6 i
rlabel alu1 60 80 60 80 6 i
rlabel alu1 90 6 90 6 6 vss
rlabel alu1 90 94 90 94 6 vdd
rlabel alu1 160 50 160 50 6 q
<< end >>
