magic
tech scmos
timestamp 1199202262
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 33 31 35
rect 9 31 19 33
rect 21 31 27 33
rect 29 31 31 33
rect 9 29 31 31
rect 9 26 11 29
rect 19 26 21 29
rect 9 2 11 6
rect 19 2 21 6
<< ndif >>
rect 2 17 9 26
rect 2 15 4 17
rect 6 15 9 17
rect 2 10 9 15
rect 2 8 4 10
rect 6 8 9 10
rect 2 6 9 8
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 11 15 14 17
rect 16 15 19 17
rect 11 6 19 15
rect 21 24 29 26
rect 21 22 24 24
rect 26 22 29 24
rect 21 17 29 22
rect 21 15 24 17
rect 26 15 29 17
rect 21 13 29 15
rect 21 6 27 13
<< pdif >>
rect 4 51 9 65
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 63 19 65
rect 11 61 14 63
rect 16 61 19 63
rect 11 55 19 61
rect 11 53 14 55
rect 16 53 19 55
rect 11 38 19 53
rect 21 49 29 65
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 63 38 65
rect 31 61 34 63
rect 36 61 38 63
rect 31 55 38 61
rect 31 53 34 55
rect 36 53 38 55
rect 31 38 38 53
<< alu1 >>
rect -2 64 42 72
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 23 49 27 51
rect 23 47 24 49
rect 26 47 27 49
rect 23 42 27 47
rect 2 40 4 42
rect 6 40 24 42
rect 26 40 27 42
rect 2 38 27 40
rect 2 26 6 38
rect 34 34 38 43
rect 17 33 38 34
rect 17 31 19 33
rect 21 31 27 33
rect 29 31 38 33
rect 17 30 38 31
rect 2 24 17 26
rect 2 22 14 24
rect 16 22 17 24
rect 13 17 17 22
rect 13 15 14 17
rect 16 15 17 17
rect 13 13 17 15
rect 34 21 38 30
rect -2 7 42 8
rect -2 5 33 7
rect 35 5 42 7
rect -2 0 42 5
<< ptie >>
rect 31 7 37 9
rect 31 5 33 7
rect 35 5 37 7
rect 31 3 37 5
<< nmos >>
rect 9 6 11 26
rect 19 6 21 26
<< pmos >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
<< polyct1 >>
rect 19 31 21 33
rect 27 31 29 33
<< ndifct0 >>
rect 4 15 6 17
rect 4 8 6 10
rect 24 22 26 24
rect 24 15 26 17
<< ndifct1 >>
rect 14 22 16 24
rect 14 15 16 17
<< ptiect1 >>
rect 33 5 35 7
<< pdifct0 >>
rect 14 61 16 63
rect 14 53 16 55
rect 34 61 36 63
rect 34 53 36 55
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 24 47 26 49
rect 24 40 26 42
<< alu0 >>
rect 13 63 17 64
rect 13 61 14 63
rect 16 61 17 63
rect 13 55 17 61
rect 13 53 14 55
rect 16 53 17 55
rect 13 51 17 53
rect 33 63 37 64
rect 33 61 34 63
rect 36 61 37 63
rect 33 55 37 61
rect 33 53 34 55
rect 36 53 37 55
rect 33 51 37 53
rect 2 17 8 18
rect 2 15 4 17
rect 6 15 8 17
rect 2 10 8 15
rect 22 24 28 25
rect 22 22 24 24
rect 26 22 28 24
rect 22 17 28 22
rect 22 15 24 17
rect 26 15 28 17
rect 2 8 4 10
rect 6 8 8 10
rect 22 8 28 15
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel polyct1 20 32 20 32 6 a
rlabel alu1 20 40 20 40 6 z
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 36 32 36 32 6 a
<< end >>
