magic
tech scmos
timestamp 1199973020
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -5 40 101 97
<< pwell >>
rect -5 -9 101 40
<< poly >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 81 75 83
rect 66 79 71 81
rect 73 79 75 81
rect 66 77 75 79
rect 53 74 55 77
rect 73 74 75 77
rect 85 81 94 83
rect 85 79 87 81
rect 89 79 94 81
rect 85 77 94 79
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 41 14 43
rect 2 39 7 41
rect 9 39 14 41
rect 2 37 14 39
rect 18 41 30 43
rect 18 39 23 41
rect 25 39 30 41
rect 18 37 30 39
rect 34 41 46 43
rect 34 39 39 41
rect 41 39 46 41
rect 34 37 46 39
rect 50 41 62 43
rect 50 39 55 41
rect 57 39 62 41
rect 50 37 62 39
rect 66 41 78 43
rect 66 39 68 41
rect 70 39 78 41
rect 66 37 78 39
rect 82 37 94 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 5 62 11
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndif >>
rect 2 25 9 34
rect 2 23 4 25
rect 6 23 9 25
rect 2 18 9 23
rect 2 16 4 18
rect 6 16 9 18
rect 2 14 9 16
rect 11 28 21 34
rect 11 26 15 28
rect 17 26 21 28
rect 11 21 21 26
rect 11 19 15 21
rect 17 19 21 21
rect 11 14 21 19
rect 23 18 30 34
rect 23 16 26 18
rect 28 16 30 18
rect 23 14 30 16
rect 34 18 41 34
rect 34 16 36 18
rect 38 16 41 18
rect 34 14 41 16
rect 43 29 53 34
rect 43 27 47 29
rect 49 27 53 29
rect 43 21 53 27
rect 43 19 47 21
rect 49 19 53 21
rect 43 14 53 19
rect 55 18 62 34
rect 55 16 58 18
rect 60 16 62 18
rect 55 14 62 16
rect 66 18 73 34
rect 66 16 68 18
rect 70 16 73 18
rect 66 14 73 16
rect 75 29 85 34
rect 75 27 79 29
rect 81 27 85 29
rect 75 21 85 27
rect 75 19 79 21
rect 81 19 85 21
rect 75 14 85 19
rect 87 25 94 34
rect 87 23 90 25
rect 92 23 94 25
rect 87 18 94 23
rect 87 16 90 18
rect 92 16 94 18
rect 87 14 94 16
rect 13 2 19 14
rect 45 2 51 14
rect 77 2 83 14
<< pdif >>
rect 13 74 19 86
rect 45 74 51 86
rect 77 74 83 86
rect 2 72 9 74
rect 2 70 4 72
rect 6 70 9 72
rect 2 65 9 70
rect 2 63 4 65
rect 6 63 9 65
rect 2 46 9 63
rect 11 61 21 74
rect 11 59 15 61
rect 17 59 21 61
rect 11 54 21 59
rect 11 52 15 54
rect 17 52 21 54
rect 11 46 21 52
rect 23 72 30 74
rect 23 70 26 72
rect 28 70 30 72
rect 23 65 30 70
rect 23 63 26 65
rect 28 63 30 65
rect 23 46 30 63
rect 34 72 41 74
rect 34 70 36 72
rect 38 70 41 72
rect 34 65 41 70
rect 34 63 36 65
rect 38 63 41 65
rect 34 46 41 63
rect 43 61 53 74
rect 43 59 47 61
rect 49 59 53 61
rect 43 53 53 59
rect 43 51 47 53
rect 49 51 53 53
rect 43 46 53 51
rect 55 72 62 74
rect 55 70 58 72
rect 60 70 62 72
rect 55 65 62 70
rect 55 63 58 65
rect 60 63 62 65
rect 55 46 62 63
rect 66 72 73 74
rect 66 70 68 72
rect 70 70 73 72
rect 66 65 73 70
rect 66 63 68 65
rect 70 63 73 65
rect 66 46 73 63
rect 75 61 85 74
rect 75 59 79 61
rect 81 59 85 61
rect 75 53 85 59
rect 75 51 79 53
rect 81 51 85 53
rect 75 46 85 51
rect 87 71 94 74
rect 87 69 90 71
rect 92 69 94 71
rect 87 64 94 69
rect 87 62 90 64
rect 92 62 94 64
rect 87 46 94 62
<< alu1 >>
rect -2 89 98 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 73 87 87 89
rect 89 87 91 89
rect 93 87 98 89
rect -2 86 98 87
rect 3 81 7 86
rect 3 79 4 81
rect 6 79 7 81
rect 3 72 7 79
rect 3 70 4 72
rect 6 70 7 72
rect 3 65 7 70
rect 3 63 4 65
rect 6 63 7 65
rect 25 81 29 86
rect 25 79 26 81
rect 28 79 29 81
rect 25 72 29 79
rect 25 70 26 72
rect 28 70 29 72
rect 25 65 29 70
rect 25 63 26 65
rect 28 63 29 65
rect 3 61 7 63
rect 14 61 18 63
rect 25 61 29 63
rect 35 81 39 86
rect 35 79 36 81
rect 38 79 39 81
rect 35 72 39 79
rect 35 70 36 72
rect 38 70 39 72
rect 35 65 39 70
rect 35 63 36 65
rect 38 63 39 65
rect 57 81 61 86
rect 57 79 58 81
rect 60 79 61 81
rect 57 73 61 79
rect 57 72 93 73
rect 57 70 58 72
rect 60 70 68 72
rect 70 71 93 72
rect 70 70 90 71
rect 57 69 90 70
rect 92 69 93 71
rect 57 65 61 69
rect 57 63 58 65
rect 60 63 61 65
rect 35 61 39 63
rect 46 61 50 63
rect 57 61 61 63
rect 67 65 71 69
rect 67 63 68 65
rect 70 63 71 65
rect 89 64 93 69
rect 67 61 71 63
rect 78 61 82 63
rect 14 59 15 61
rect 17 59 18 61
rect 6 41 10 55
rect 14 54 18 59
rect 46 59 47 61
rect 49 59 50 61
rect 46 54 50 59
rect 78 59 79 61
rect 81 59 82 61
rect 89 62 90 64
rect 92 62 93 64
rect 89 60 93 62
rect 78 54 82 59
rect 14 52 15 54
rect 17 53 82 54
rect 17 52 47 53
rect 14 51 47 52
rect 49 51 79 53
rect 81 51 82 53
rect 14 50 82 51
rect 6 39 7 41
rect 9 39 10 41
rect 6 38 10 39
rect 22 41 26 43
rect 22 39 23 41
rect 25 39 26 41
rect 22 38 26 39
rect 38 41 42 43
rect 38 39 39 41
rect 41 39 42 41
rect 38 38 42 39
rect 54 41 58 43
rect 54 39 55 41
rect 57 39 58 41
rect 54 38 58 39
rect 67 41 71 43
rect 67 39 68 41
rect 70 39 71 41
rect 67 38 71 39
rect 6 34 71 38
rect 6 33 10 34
rect 78 30 82 50
rect 14 29 82 30
rect 14 28 47 29
rect 3 25 7 27
rect 3 23 4 25
rect 6 23 7 25
rect 3 18 7 23
rect 3 16 4 18
rect 6 16 7 18
rect 14 26 15 28
rect 17 27 47 28
rect 49 27 79 29
rect 81 27 82 29
rect 17 26 82 27
rect 14 21 18 26
rect 14 19 15 21
rect 17 19 18 21
rect 46 21 50 26
rect 14 17 18 19
rect 25 18 29 20
rect 3 9 7 16
rect 3 7 4 9
rect 6 7 7 9
rect 3 2 7 7
rect 25 16 26 18
rect 28 16 29 18
rect 25 9 29 16
rect 25 7 26 9
rect 28 7 29 9
rect 25 2 29 7
rect 35 18 39 20
rect 35 16 36 18
rect 38 16 39 18
rect 46 19 47 21
rect 49 19 50 21
rect 78 21 82 26
rect 46 17 50 19
rect 57 18 61 20
rect 35 9 39 16
rect 35 7 36 9
rect 38 7 39 9
rect 35 2 39 7
rect 57 16 58 18
rect 60 16 61 18
rect 57 9 61 16
rect 57 7 58 9
rect 60 7 61 9
rect 57 2 61 7
rect 67 18 71 20
rect 67 16 68 18
rect 70 16 71 18
rect 78 19 79 21
rect 81 19 82 21
rect 78 17 82 19
rect 89 25 93 27
rect 89 23 90 25
rect 92 23 93 25
rect 89 18 93 23
rect 67 9 71 16
rect 67 7 68 9
rect 70 7 71 9
rect 67 2 71 7
rect 89 16 90 18
rect 92 16 93 18
rect 89 9 93 16
rect 89 7 90 9
rect 92 7 93 9
rect 89 2 93 7
rect -2 1 98 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 73 -1 87 1
rect 89 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< alu2 >>
rect -2 89 98 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 71 89
rect 73 87 87 89
rect 89 87 98 89
rect -2 81 98 87
rect -2 79 4 81
rect 6 79 26 81
rect 28 79 36 81
rect 38 79 58 81
rect 60 79 98 81
rect -2 76 98 79
rect -2 9 98 12
rect -2 7 4 9
rect 6 7 26 9
rect 28 7 36 9
rect 38 7 58 9
rect 60 7 68 9
rect 70 7 90 9
rect 92 7 98 9
rect -2 1 98 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 71 1
rect 73 -1 87 1
rect 89 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 71 3
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 57 -3 71 -1
rect 89 1 96 3
rect 89 -1 91 1
rect 93 -1 96 1
rect 89 -3 96 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 71 91
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 57 85 71 87
rect 89 89 96 91
rect 89 87 91 89
rect 93 87 96 89
rect 89 85 96 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polyct0 >>
rect 71 79 73 81
rect 87 79 89 81
<< polyct1 >>
rect 7 39 9 41
rect 23 39 25 41
rect 39 39 41 41
rect 55 39 57 41
rect 68 39 70 41
<< ndifct1 >>
rect 4 23 6 25
rect 4 16 6 18
rect 15 26 17 28
rect 15 19 17 21
rect 26 16 28 18
rect 36 16 38 18
rect 47 27 49 29
rect 47 19 49 21
rect 58 16 60 18
rect 68 16 70 18
rect 79 27 81 29
rect 79 19 81 21
rect 90 23 92 25
rect 90 16 92 18
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
rect 67 87 69 89
rect 91 87 93 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 91 -1 93 1
<< pdifct1 >>
rect 4 70 6 72
rect 4 63 6 65
rect 15 59 17 61
rect 15 52 17 54
rect 26 70 28 72
rect 26 63 28 65
rect 36 70 38 72
rect 36 63 38 65
rect 47 59 49 61
rect 47 51 49 53
rect 58 70 60 72
rect 58 63 60 65
rect 68 70 70 72
rect 68 63 70 65
rect 79 59 81 61
rect 79 51 81 53
rect 90 69 92 71
rect 90 62 92 64
<< alu0 >>
rect 69 81 91 82
rect 69 79 71 81
rect 73 79 87 81
rect 89 79 91 81
rect 69 78 91 79
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 71 87 73 89
rect 87 87 89 89
rect 4 79 6 81
rect 26 79 28 81
rect 36 79 38 81
rect 58 79 60 81
rect 4 7 6 9
rect 26 7 28 9
rect 36 7 38 9
rect 58 7 60 9
rect 68 7 70 9
rect 90 7 92 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
rect 71 -1 73 1
rect 87 -1 89 1
<< labels >>
rlabel alu1 8 44 8 44 6 a
rlabel ndifct1 16 20 16 20 6 z
rlabel alu1 24 28 24 28 6 z
rlabel alu1 32 28 32 28 6 z
rlabel alu1 24 36 24 36 6 a
rlabel alu1 32 36 32 36 6 a
rlabel alu1 16 36 16 36 6 a
rlabel alu1 24 52 24 52 6 z
rlabel alu1 32 52 32 52 6 z
rlabel pdifct1 16 60 16 60 6 z
rlabel alu1 40 28 40 28 6 z
rlabel alu1 56 28 56 28 6 z
rlabel alu1 48 24 48 24 6 z
rlabel alu1 48 36 48 36 6 a
rlabel alu1 56 36 56 36 6 a
rlabel alu1 40 36 40 36 6 a
rlabel alu1 56 52 56 52 6 z
rlabel alu1 48 56 48 56 6 z
rlabel alu1 40 52 40 52 6 z
rlabel alu1 64 28 64 28 6 z
rlabel alu1 72 28 72 28 6 z
rlabel alu1 64 36 64 36 6 a
rlabel alu1 64 52 64 52 6 z
rlabel alu1 72 52 72 52 6 z
rlabel alu1 80 40 80 40 6 z
rlabel alu2 16 6 16 6 6 vss
rlabel alu2 48 6 48 6 6 vss
rlabel alu2 48 82 48 82 6 vdd
<< end >>
