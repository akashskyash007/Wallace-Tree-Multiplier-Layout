magic
tech scmos
timestamp 1199202291
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 9 35 11 38
rect 19 35 21 38
rect 9 33 21 35
rect 9 31 17 33
rect 19 31 21 33
rect 9 29 21 31
rect 9 26 11 29
rect 19 26 21 29
rect 9 2 11 7
rect 19 2 21 7
<< ndif >>
rect 2 18 9 26
rect 2 16 4 18
rect 6 16 9 18
rect 2 11 9 16
rect 2 9 4 11
rect 6 9 9 11
rect 2 7 9 9
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 11 15 14 17
rect 16 15 19 17
rect 11 7 19 15
rect 21 18 29 26
rect 21 16 24 18
rect 26 16 29 18
rect 21 11 29 16
rect 21 9 24 11
rect 26 9 29 11
rect 21 7 29 9
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
<< alu1 >>
rect -2 64 34 72
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 50 17 55
rect 2 48 14 50
rect 16 48 17 50
rect 2 46 17 48
rect 2 26 6 46
rect 26 34 30 43
rect 15 33 30 34
rect 15 31 17 33
rect 19 31 30 33
rect 15 30 30 31
rect 2 24 23 26
rect 2 22 14 24
rect 16 22 23 24
rect 13 17 17 22
rect 13 15 14 17
rect 16 15 17 17
rect 13 13 17 15
rect -2 0 34 8
<< nmos >>
rect 9 7 11 26
rect 19 7 21 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
<< polyct1 >>
rect 17 31 19 33
<< ndifct0 >>
rect 4 16 6 18
rect 4 9 6 11
rect 24 16 26 18
rect 24 9 26 11
<< ndifct1 >>
rect 14 22 16 24
rect 14 15 16 17
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 24 62 26 64
rect 24 55 26 57
<< pdifct1 >>
rect 14 55 16 57
rect 14 48 16 50
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 22 57 28 62
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 2 18 8 19
rect 2 16 4 18
rect 6 16 8 18
rect 2 11 8 16
rect 22 18 28 19
rect 22 16 24 18
rect 26 16 28 18
rect 2 9 4 11
rect 6 9 8 11
rect 2 8 8 9
rect 22 11 28 16
rect 22 9 24 11
rect 26 9 28 11
rect 22 8 28 9
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 32 20 32 6 a
rlabel alu1 20 24 20 24 6 z
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 40 28 40 6 a
<< end >>
