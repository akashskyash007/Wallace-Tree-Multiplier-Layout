magic
tech scmos
timestamp 1199203555
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 69 31 74
rect 36 72 64 74
rect 36 69 38 72
rect 55 64 57 68
rect 62 64 64 72
rect 74 70 76 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 29 34 31 42
rect 36 38 38 42
rect 55 39 57 42
rect 51 37 57 39
rect 51 35 53 37
rect 55 35 57 37
rect 51 34 57 35
rect 10 24 12 33
rect 19 29 21 33
rect 29 32 57 34
rect 62 38 64 42
rect 74 39 76 42
rect 62 36 70 38
rect 62 34 66 36
rect 68 34 70 36
rect 62 32 70 34
rect 74 37 81 39
rect 74 35 77 37
rect 79 35 81 37
rect 74 33 81 35
rect 17 27 21 29
rect 37 28 39 32
rect 62 29 64 32
rect 74 29 76 33
rect 17 24 19 27
rect 27 24 29 28
rect 37 12 39 16
rect 62 12 64 16
rect 10 6 12 11
rect 17 6 19 11
rect 27 8 29 11
rect 74 8 76 16
rect 27 6 76 8
<< ndif >>
rect 32 24 37 28
rect 2 11 10 24
rect 12 11 17 24
rect 19 21 27 24
rect 19 19 22 21
rect 24 19 27 21
rect 19 11 27 19
rect 29 22 37 24
rect 29 20 32 22
rect 34 20 37 22
rect 29 16 37 20
rect 39 20 46 28
rect 39 18 42 20
rect 44 18 46 20
rect 39 16 46 18
rect 55 27 62 29
rect 55 25 57 27
rect 59 25 62 27
rect 55 20 62 25
rect 55 18 57 20
rect 59 18 62 20
rect 55 16 62 18
rect 64 20 74 29
rect 64 18 69 20
rect 71 18 74 20
rect 64 16 74 18
rect 76 22 81 29
rect 76 20 83 22
rect 76 18 79 20
rect 81 18 83 20
rect 76 16 83 18
rect 29 11 34 16
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
<< pdif >>
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 42 9 58
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 69 26 70
rect 21 53 29 69
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 42 36 69
rect 38 67 46 69
rect 38 65 41 67
rect 43 65 46 67
rect 38 54 46 65
rect 66 68 74 70
rect 66 66 69 68
rect 71 66 74 68
rect 66 64 74 66
rect 38 42 44 54
rect 50 48 55 64
rect 48 46 55 48
rect 48 44 50 46
rect 52 44 55 46
rect 48 42 55 44
rect 57 42 62 64
rect 64 42 74 64
rect 76 63 81 70
rect 76 61 83 63
rect 76 59 79 61
rect 81 59 83 61
rect 76 57 83 59
rect 76 42 81 57
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 2 53 18 54
rect 2 51 14 53
rect 16 51 18 53
rect 2 50 18 51
rect 2 22 6 50
rect 58 39 62 55
rect 66 49 78 55
rect 50 37 62 39
rect 50 35 53 37
rect 55 35 62 37
rect 50 33 62 35
rect 66 36 70 39
rect 68 34 70 36
rect 74 38 78 49
rect 74 37 81 38
rect 74 35 77 37
rect 79 35 81 37
rect 74 34 81 35
rect 66 30 70 34
rect 66 25 79 30
rect 2 21 26 22
rect 2 19 22 21
rect 24 19 26 21
rect 2 18 26 19
rect -2 11 98 12
rect -2 9 4 11
rect 6 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 10 11 12 24
rect 17 11 19 24
rect 27 11 29 24
rect 37 16 39 28
rect 62 16 64 29
rect 74 16 76 29
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 69
rect 36 42 38 69
rect 55 42 57 64
rect 62 42 64 64
rect 74 42 76 70
<< polyct0 >>
rect 11 35 13 37
rect 21 35 23 37
<< polyct1 >>
rect 53 35 55 37
rect 66 34 68 36
rect 77 35 79 37
<< ndifct0 >>
rect 32 20 34 22
rect 42 18 44 20
rect 57 25 59 27
rect 57 18 59 20
rect 69 18 71 20
rect 79 18 81 20
<< ndifct1 >>
rect 22 19 24 21
rect 4 9 6 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 60 6 62
rect 24 51 26 53
rect 24 44 26 46
rect 41 65 43 67
rect 69 66 71 68
rect 50 44 52 46
rect 79 59 81 61
<< pdifct1 >>
rect 14 51 16 53
<< alu0 >>
rect 40 67 44 68
rect 40 65 41 67
rect 43 65 44 67
rect 67 66 69 68
rect 71 66 73 68
rect 67 65 73 66
rect 40 63 44 65
rect 2 62 36 63
rect 2 60 4 62
rect 6 60 36 62
rect 2 59 36 60
rect 50 61 89 62
rect 50 59 79 61
rect 81 59 89 61
rect 32 58 89 59
rect 32 55 54 58
rect 23 53 27 55
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 10 44 24 46
rect 26 44 27 46
rect 10 42 27 44
rect 10 37 14 42
rect 32 38 36 55
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 19 37 36 38
rect 19 35 21 37
rect 23 35 36 37
rect 19 34 36 35
rect 42 46 54 47
rect 42 44 50 46
rect 52 44 54 46
rect 42 43 54 44
rect 10 29 35 30
rect 42 29 46 43
rect 65 32 66 38
rect 10 27 61 29
rect 10 26 57 27
rect 31 25 57 26
rect 59 25 61 27
rect 31 22 35 25
rect 31 20 32 22
rect 34 20 35 22
rect 31 18 35 20
rect 40 20 46 21
rect 40 18 42 20
rect 44 18 46 20
rect 40 12 46 18
rect 55 20 61 25
rect 85 21 89 58
rect 55 18 57 20
rect 59 18 61 20
rect 55 17 61 18
rect 67 20 73 21
rect 67 18 69 20
rect 71 18 73 20
rect 67 12 73 18
rect 77 20 89 21
rect 77 18 79 20
rect 81 18 89 20
rect 77 17 89 18
<< labels >>
rlabel polyct0 12 36 12 36 6 an
rlabel alu0 33 24 33 24 6 an
rlabel alu0 27 36 27 36 6 bn
rlabel alu0 25 48 25 48 6 an
rlabel alu0 19 61 19 61 6 bn
rlabel alu0 58 23 58 23 6 an
rlabel alu0 48 45 48 45 6 an
rlabel alu0 83 19 83 19 6 bn
rlabel alu0 69 60 69 60 6 bn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 52 36 52 36 6 a2
rlabel alu1 68 32 68 32 6 a1
rlabel alu1 60 44 60 44 6 a2
rlabel alu1 68 52 68 52 6 b
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 76 28 76 28 6 a1
rlabel alu1 76 48 76 48 6 b
<< end >>
