magic
tech scmos
timestamp 1199203078
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 64 11 69
rect 21 60 23 65
rect 9 37 11 52
rect 44 58 46 63
rect 54 58 56 63
rect 61 58 63 63
rect 21 47 23 50
rect 15 45 23 47
rect 44 46 46 50
rect 15 43 17 45
rect 19 44 23 45
rect 40 44 46 46
rect 19 43 21 44
rect 15 41 21 43
rect 9 35 15 37
rect 9 33 11 35
rect 13 33 15 35
rect 9 31 15 33
rect 9 28 11 31
rect 19 29 21 41
rect 40 39 42 44
rect 54 39 56 42
rect 25 37 42 39
rect 25 35 27 37
rect 29 35 31 37
rect 25 33 31 35
rect 40 30 42 37
rect 49 37 56 39
rect 49 35 51 37
rect 53 35 56 37
rect 49 33 56 35
rect 61 39 63 42
rect 61 37 67 39
rect 61 35 63 37
rect 65 35 67 37
rect 61 33 67 35
rect 50 30 52 33
rect 19 26 22 29
rect 20 23 22 26
rect 61 23 63 33
rect 9 17 11 22
rect 40 18 42 23
rect 50 18 52 23
rect 20 12 22 17
rect 61 11 63 16
<< ndif >>
rect 2 26 9 28
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 11 23 17 28
rect 33 28 40 30
rect 33 26 35 28
rect 37 26 40 28
rect 33 23 40 26
rect 42 28 50 30
rect 42 26 45 28
rect 47 26 50 28
rect 42 23 50 26
rect 52 23 59 30
rect 11 22 20 23
rect 13 21 20 22
rect 13 19 15 21
rect 17 19 20 21
rect 13 17 20 19
rect 22 21 29 23
rect 22 19 25 21
rect 27 19 29 21
rect 22 17 29 19
rect 54 20 61 23
rect 54 18 56 20
rect 58 18 61 20
rect 54 16 61 18
rect 63 21 70 23
rect 63 19 66 21
rect 68 19 70 21
rect 63 16 70 19
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 64 19 69
rect 35 71 42 73
rect 35 69 38 71
rect 40 69 42 71
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 52 9 58
rect 11 60 19 64
rect 11 52 21 60
rect 13 50 21 52
rect 23 56 28 60
rect 35 58 42 69
rect 23 54 31 56
rect 23 52 27 54
rect 29 52 31 54
rect 23 50 31 52
rect 35 50 44 58
rect 46 54 54 58
rect 46 52 49 54
rect 51 52 54 54
rect 46 50 54 52
rect 49 42 54 50
rect 56 42 61 58
rect 63 56 70 58
rect 63 54 66 56
rect 68 54 70 56
rect 63 42 70 54
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 71 74 79
rect -2 69 15 71
rect 17 69 38 71
rect 40 69 74 71
rect -2 68 74 69
rect 10 46 14 55
rect 10 45 23 46
rect 10 43 17 45
rect 19 43 23 45
rect 10 42 23 43
rect 10 35 23 38
rect 10 33 11 35
rect 13 34 23 35
rect 13 33 14 34
rect 10 25 14 33
rect 34 54 54 55
rect 34 52 49 54
rect 51 52 54 54
rect 34 49 54 52
rect 34 28 38 49
rect 66 39 70 47
rect 58 37 70 39
rect 58 35 63 37
rect 65 35 70 37
rect 58 33 70 35
rect 34 26 35 28
rect 37 26 38 28
rect 34 17 38 26
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 9 22 11 28
rect 40 23 42 30
rect 50 23 52 30
rect 20 17 22 23
rect 61 16 63 23
<< pmos >>
rect 9 52 11 64
rect 21 50 23 60
rect 44 50 46 58
rect 54 42 56 58
rect 61 42 63 58
<< polyct0 >>
rect 27 35 29 37
rect 51 35 53 37
<< polyct1 >>
rect 17 43 19 45
rect 11 33 13 35
rect 63 35 65 37
<< ndifct0 >>
rect 4 24 6 26
rect 45 26 47 28
rect 15 19 17 21
rect 25 19 27 21
rect 56 18 58 20
rect 66 19 68 21
<< ndifct1 >>
rect 35 26 37 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 60 6 62
rect 27 52 29 54
rect 66 54 68 56
<< pdifct1 >>
rect 15 69 17 71
rect 38 69 40 71
rect 49 52 51 54
<< alu0 >>
rect 2 62 62 63
rect 2 60 4 62
rect 6 60 62 62
rect 2 59 62 60
rect 2 28 6 59
rect 26 54 30 56
rect 26 52 27 54
rect 29 52 30 54
rect 26 37 30 52
rect 26 35 27 37
rect 29 35 30 37
rect 2 26 7 28
rect 2 24 4 26
rect 6 24 7 26
rect 26 30 30 35
rect 24 26 30 30
rect 58 46 62 59
rect 65 56 69 68
rect 65 54 66 56
rect 68 54 69 56
rect 65 52 69 54
rect 50 42 62 46
rect 50 37 54 42
rect 50 35 51 37
rect 53 35 54 37
rect 50 33 54 35
rect 2 22 7 24
rect 13 21 19 22
rect 13 19 15 21
rect 17 19 19 21
rect 13 12 19 19
rect 24 21 28 26
rect 24 19 25 21
rect 27 19 28 21
rect 24 17 28 19
rect 43 28 69 29
rect 43 26 45 28
rect 47 26 69 28
rect 43 25 69 26
rect 65 21 69 25
rect 54 20 60 21
rect 54 18 56 20
rect 58 18 60 20
rect 54 12 60 18
rect 65 19 66 21
rect 68 19 69 21
rect 65 17 69 19
<< labels >>
rlabel alu0 4 42 4 42 6 a2n
rlabel alu0 26 23 26 23 6 bn
rlabel alu0 28 41 28 41 6 bn
rlabel alu0 67 23 67 23 6 n1
rlabel alu0 56 27 56 27 6 n1
rlabel alu0 52 39 52 39 6 a2n
rlabel alu0 32 61 32 61 6 a2n
rlabel alu1 12 28 12 28 6 a2
rlabel alu1 12 52 12 52 6 b
rlabel alu1 20 36 20 36 6 a2
rlabel alu1 20 44 20 44 6 b
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 36 36 36 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 36 60 36 6 a1
rlabel alu1 68 40 68 40 6 a1
<< end >>
