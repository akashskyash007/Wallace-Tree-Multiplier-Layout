magic
tech scmos
timestamp 1199202668
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 14 54 16 59
rect 24 54 26 59
rect 35 54 37 59
rect 45 54 47 59
rect 14 35 16 38
rect 24 35 26 38
rect 35 35 37 38
rect 45 35 47 38
rect 9 33 26 35
rect 9 31 11 33
rect 13 31 26 33
rect 9 29 26 31
rect 24 26 26 29
rect 31 33 47 35
rect 31 31 43 33
rect 45 31 47 33
rect 31 29 47 31
rect 31 26 33 29
rect 24 8 26 13
rect 31 8 33 13
<< ndif >>
rect 17 24 24 26
rect 17 22 19 24
rect 21 22 24 24
rect 17 17 24 22
rect 17 15 19 17
rect 21 15 24 17
rect 17 13 24 15
rect 26 13 31 26
rect 33 24 41 26
rect 33 22 36 24
rect 38 22 41 24
rect 33 17 41 22
rect 33 15 36 17
rect 38 15 41 17
rect 33 13 41 15
<< pdif >>
rect 6 52 14 54
rect 6 50 9 52
rect 11 50 14 52
rect 6 38 14 50
rect 16 49 24 54
rect 16 47 19 49
rect 21 47 24 49
rect 16 42 24 47
rect 16 40 19 42
rect 21 40 24 42
rect 16 38 24 40
rect 26 52 35 54
rect 26 50 29 52
rect 31 50 35 52
rect 26 38 35 50
rect 37 49 45 54
rect 37 47 40 49
rect 42 47 45 49
rect 37 42 45 47
rect 37 40 40 42
rect 42 40 45 42
rect 37 38 45 40
rect 47 52 54 54
rect 47 50 50 52
rect 52 50 54 52
rect 47 45 54 50
rect 47 43 50 45
rect 52 43 54 45
rect 47 38 54 43
<< alu1 >>
rect -2 67 58 72
rect -2 65 41 67
rect 43 65 49 67
rect 51 65 58 67
rect -2 64 58 65
rect 18 49 22 51
rect 18 47 19 49
rect 21 47 22 49
rect 39 49 43 51
rect 2 35 6 43
rect 18 42 22 47
rect 39 47 40 49
rect 42 47 43 49
rect 39 42 43 47
rect 18 40 19 42
rect 21 40 40 42
rect 42 40 43 42
rect 18 38 43 40
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 18 24 22 38
rect 41 33 54 34
rect 41 31 43 33
rect 45 31 54 33
rect 41 30 54 31
rect 18 22 19 24
rect 21 22 22 24
rect 18 17 22 22
rect 18 15 19 17
rect 21 15 22 17
rect 18 13 22 15
rect 50 21 54 30
rect -2 7 58 8
rect -2 5 5 7
rect 7 5 49 7
rect 51 5 58 7
rect -2 0 58 5
<< ptie >>
rect 3 7 9 24
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 47 7 53 24
rect 47 5 49 7
rect 51 5 53 7
rect 47 3 53 5
<< ntie >>
rect 39 67 53 69
rect 39 65 41 67
rect 43 65 49 67
rect 51 65 53 67
rect 39 63 53 65
<< nmos >>
rect 24 13 26 26
rect 31 13 33 26
<< pmos >>
rect 14 38 16 54
rect 24 38 26 54
rect 35 38 37 54
rect 45 38 47 54
<< polyct1 >>
rect 11 31 13 33
rect 43 31 45 33
<< ndifct0 >>
rect 36 22 38 24
rect 36 15 38 17
<< ndifct1 >>
rect 19 22 21 24
rect 19 15 21 17
<< ntiect1 >>
rect 41 65 43 67
rect 49 65 51 67
<< ptiect1 >>
rect 5 5 7 7
rect 49 5 51 7
<< pdifct0 >>
rect 9 50 11 52
rect 29 50 31 52
rect 50 50 52 52
rect 50 43 52 45
<< pdifct1 >>
rect 19 47 21 49
rect 19 40 21 42
rect 40 47 42 49
rect 40 40 42 42
<< alu0 >>
rect 8 52 12 64
rect 8 50 9 52
rect 11 50 12 52
rect 28 52 32 64
rect 8 48 12 50
rect 28 50 29 52
rect 31 50 32 52
rect 49 52 53 64
rect 28 48 32 50
rect 49 50 50 52
rect 52 50 53 52
rect 49 45 53 50
rect 49 43 50 45
rect 52 43 53 45
rect 49 41 53 43
rect 35 24 39 26
rect 35 22 36 24
rect 38 22 39 24
rect 35 17 39 22
rect 35 15 36 17
rect 38 15 39 17
rect 35 8 39 15
<< labels >>
rlabel alu1 4 36 4 36 6 b
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 20 32 20 32 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 40 36 40 6 z
rlabel alu1 28 40 28 40 6 z
rlabel alu1 28 68 28 68 6 vdd
rlabel polyct1 44 32 44 32 6 a
rlabel alu1 52 24 52 24 6 a
<< end >>
