magic
tech scmos
timestamp 1199202683
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 50 56 52 61
rect 60 56 62 61
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 50 39 52 42
rect 60 39 62 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 19 33 31 35
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 37 52 39
rect 56 37 62 39
rect 36 35 43 37
rect 45 35 47 37
rect 36 33 47 35
rect 56 35 58 37
rect 60 35 62 37
rect 56 33 62 35
rect 36 30 38 33
rect 12 12 14 17
rect 19 12 21 17
rect 29 12 31 17
rect 36 12 38 17
<< ndif >>
rect 3 17 12 30
rect 14 17 19 30
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 17 29 19
rect 31 17 36 30
rect 38 17 47 30
rect 3 11 10 17
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
rect 40 11 47 17
rect 40 9 42 11
rect 44 9 47 11
rect 40 7 47 9
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 42 9 62
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 53 19 59
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 42 29 62
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 64 48 66
rect 41 62 44 64
rect 46 62 48 64
rect 41 56 48 62
rect 41 42 50 56
rect 52 53 60 56
rect 52 51 55 53
rect 57 51 60 53
rect 52 42 60 51
rect 62 54 70 56
rect 62 52 65 54
rect 67 52 70 54
rect 62 46 70 52
rect 62 44 65 46
rect 67 44 70 46
rect 62 42 70 44
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 2 53 59 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 51 55 53
rect 57 51 59 53
rect 2 50 59 51
rect 2 22 6 50
rect 25 42 57 46
rect 10 37 21 39
rect 10 35 11 37
rect 13 35 21 37
rect 10 33 21 35
rect 25 37 31 42
rect 53 38 57 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 17 30 21 33
rect 41 30 47 35
rect 53 37 63 38
rect 53 35 58 37
rect 60 35 63 37
rect 53 34 63 35
rect 17 26 47 30
rect 2 21 31 22
rect 2 19 24 21
rect 26 19 31 21
rect 2 18 31 19
rect -2 11 74 12
rect -2 9 6 11
rect 8 9 42 11
rect 44 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 12 17 14 30
rect 19 17 21 30
rect 29 17 31 30
rect 36 17 38 30
<< pmos >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
rect 50 42 52 56
rect 60 42 62 56
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 43 35 45 37
rect 58 35 60 37
<< ndifct1 >>
rect 24 19 26 21
rect 6 9 8 11
rect 42 9 44 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 62 6 64
rect 14 59 16 61
rect 24 62 26 64
rect 44 62 46 64
rect 65 52 67 54
rect 65 44 67 46
<< pdifct1 >>
rect 14 51 16 53
rect 34 59 36 61
rect 34 51 36 53
rect 55 51 57 53
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 23 64 27 68
rect 3 60 7 62
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 23 62 24 64
rect 26 62 27 64
rect 43 64 47 68
rect 23 60 27 62
rect 13 54 17 59
rect 43 62 44 64
rect 46 62 47 64
rect 43 60 47 62
rect 64 54 68 68
rect 64 52 65 54
rect 67 52 68 54
rect 64 46 68 52
rect 64 44 65 46
rect 67 44 68 46
rect 64 42 68 44
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel alu1 28 28 28 28 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 32 44 32 6 a
rlabel alu1 44 44 44 44 6 b
rlabel alu1 52 44 52 44 6 b
rlabel alu1 36 44 36 44 6 b
rlabel alu1 36 56 36 56 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 36 60 36 6 b
<< end >>
