magic
tech scmos
timestamp 1199203177
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 22 66 24 70
rect 29 66 31 70
rect 36 66 38 70
rect 46 66 48 70
rect 53 66 55 70
rect 60 66 62 70
rect 9 57 11 61
rect 9 35 11 38
rect 22 37 24 40
rect 19 35 25 37
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 21 35
rect 23 33 25 35
rect 19 31 25 33
rect 29 31 31 40
rect 36 37 38 40
rect 46 37 48 40
rect 36 35 48 37
rect 40 33 42 35
rect 44 33 46 35
rect 40 31 46 33
rect 53 31 55 40
rect 60 37 62 40
rect 60 35 70 37
rect 64 33 66 35
rect 68 33 70 35
rect 64 31 70 33
rect 9 26 11 29
rect 19 26 21 31
rect 29 29 35 31
rect 29 27 31 29
rect 33 27 35 29
rect 29 25 35 27
rect 40 22 42 31
rect 50 29 56 31
rect 50 27 52 29
rect 54 27 56 29
rect 50 25 56 27
rect 50 22 52 25
rect 9 5 11 10
rect 19 5 21 10
rect 40 2 42 6
rect 50 2 52 6
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 10 9 13
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 11 15 14 17
rect 16 15 19 17
rect 11 10 19 15
rect 21 22 26 26
rect 21 10 40 22
rect 23 7 40 10
rect 23 5 25 7
rect 27 5 34 7
rect 36 6 40 7
rect 42 16 50 22
rect 42 14 45 16
rect 47 14 50 16
rect 42 6 50 14
rect 52 17 59 22
rect 52 15 55 17
rect 57 15 59 17
rect 52 10 59 15
rect 52 8 55 10
rect 57 8 59 10
rect 52 6 59 8
rect 36 5 38 6
rect 23 3 38 5
<< pdif >>
rect 13 64 22 66
rect 13 62 16 64
rect 18 62 22 64
rect 13 57 22 62
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 48 9 53
rect 2 46 4 48
rect 6 46 9 48
rect 2 44 9 46
rect 4 38 9 44
rect 11 40 22 57
rect 24 40 29 66
rect 31 40 36 66
rect 38 57 46 66
rect 38 55 41 57
rect 43 55 46 57
rect 38 40 46 55
rect 48 40 53 66
rect 55 40 60 66
rect 62 64 70 66
rect 62 62 65 64
rect 67 62 70 64
rect 62 57 70 62
rect 62 55 65 57
rect 67 55 70 57
rect 62 40 70 55
rect 11 38 16 40
<< alu1 >>
rect -2 67 74 72
rect -2 65 5 67
rect 7 65 74 67
rect -2 64 74 65
rect 2 57 47 58
rect 2 55 41 57
rect 43 55 47 57
rect 2 53 4 55
rect 6 54 47 55
rect 2 48 6 53
rect 2 46 4 48
rect 2 25 6 46
rect 10 46 23 50
rect 31 46 70 50
rect 10 33 14 46
rect 31 42 35 46
rect 10 31 11 33
rect 13 31 14 33
rect 10 29 14 31
rect 18 38 35 42
rect 41 38 55 42
rect 18 35 24 38
rect 18 33 21 35
rect 23 33 24 35
rect 18 29 24 33
rect 41 35 47 38
rect 41 33 42 35
rect 44 33 47 35
rect 30 29 34 31
rect 41 30 47 33
rect 65 35 70 46
rect 65 33 66 35
rect 68 33 70 35
rect 65 31 70 33
rect 30 27 31 29
rect 33 27 34 29
rect 30 26 34 27
rect 2 24 8 25
rect 2 22 4 24
rect 6 22 8 24
rect 2 17 8 22
rect 2 15 4 17
rect 6 15 8 17
rect 2 13 8 15
rect 30 22 70 26
rect 66 13 70 22
rect -2 7 74 8
rect -2 5 25 7
rect 27 5 34 7
rect 36 5 65 7
rect 67 5 74 7
rect -2 0 74 5
<< ptie >>
rect 63 7 69 24
rect 63 5 65 7
rect 67 5 69 7
rect 63 3 69 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 10 11 26
rect 19 10 21 26
rect 40 6 42 22
rect 50 6 52 22
<< pmos >>
rect 9 38 11 57
rect 22 40 24 66
rect 29 40 31 66
rect 36 40 38 66
rect 46 40 48 66
rect 53 40 55 66
rect 60 40 62 66
<< polyct0 >>
rect 52 27 54 29
<< polyct1 >>
rect 11 31 13 33
rect 21 33 23 35
rect 42 33 44 35
rect 66 33 68 35
rect 31 27 33 29
<< ndifct0 >>
rect 14 22 16 24
rect 14 15 16 17
rect 45 14 47 16
rect 55 15 57 17
rect 55 8 57 10
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
rect 25 5 27 7
rect 34 5 36 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 65 5 67 7
<< pdifct0 >>
rect 16 62 18 64
rect 65 62 67 64
rect 65 55 67 57
<< pdifct1 >>
rect 4 53 6 55
rect 4 46 6 48
rect 41 55 43 57
<< alu0 >>
rect 14 62 16 64
rect 18 62 20 64
rect 14 61 20 62
rect 63 62 65 64
rect 67 62 69 64
rect 63 57 69 62
rect 63 55 65 57
rect 67 55 69 57
rect 63 54 69 55
rect 6 44 7 54
rect 51 29 55 31
rect 51 27 52 29
rect 54 27 55 29
rect 51 26 55 27
rect 13 24 17 26
rect 13 22 14 24
rect 16 22 17 24
rect 13 17 17 22
rect 53 17 59 18
rect 13 15 14 17
rect 16 16 49 17
rect 16 15 45 16
rect 13 14 45 15
rect 47 14 49 16
rect 13 13 49 14
rect 53 15 55 17
rect 57 15 59 17
rect 53 10 59 15
rect 53 8 55 10
rect 57 8 59 10
<< labels >>
rlabel alu0 15 19 15 19 6 n3
rlabel alu0 31 15 31 15 6 n3
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 32 20 32 6 a1
rlabel alu1 12 36 12 36 6 b
rlabel alu1 20 48 20 48 6 b
rlabel alu1 20 56 20 56 6 z
rlabel alu1 12 56 12 56 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 36 24 36 24 6 a2
rlabel alu1 28 40 28 40 6 a1
rlabel alu1 36 48 36 48 6 a1
rlabel alu1 36 56 36 56 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 44 24 44 24 6 a2
rlabel alu1 52 24 52 24 6 a2
rlabel alu1 44 36 44 36 6 a3
rlabel alu1 52 40 52 40 6 a3
rlabel alu1 44 48 44 48 6 a1
rlabel alu1 52 48 52 48 6 a1
rlabel alu1 44 56 44 56 6 z
rlabel alu1 68 16 68 16 6 a2
rlabel alu1 60 24 60 24 6 a2
rlabel alu1 68 40 68 40 6 a1
rlabel alu1 60 48 60 48 6 a1
<< end >>
