magic
tech scmos
timestamp 1199203180
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 22 70 24 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 70 48 74
rect 53 70 55 74
rect 60 70 62 74
rect 9 61 11 65
rect 9 39 11 42
rect 22 41 24 44
rect 19 39 25 41
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 21 39
rect 23 37 25 39
rect 19 35 25 37
rect 29 35 31 44
rect 36 41 38 44
rect 46 41 48 44
rect 36 39 48 41
rect 40 37 42 39
rect 44 37 46 39
rect 40 35 46 37
rect 53 35 55 44
rect 60 41 62 44
rect 60 39 70 41
rect 64 37 66 39
rect 68 37 70 39
rect 64 35 70 37
rect 9 30 11 33
rect 19 30 21 35
rect 29 33 35 35
rect 29 31 31 33
rect 33 31 35 33
rect 29 29 35 31
rect 40 26 42 35
rect 50 33 56 35
rect 50 31 52 33
rect 54 31 56 33
rect 50 29 56 31
rect 50 26 52 29
rect 9 9 11 14
rect 19 9 21 14
rect 40 6 42 10
rect 50 6 52 10
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 14 9 17
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 14 19 19
rect 21 26 26 30
rect 21 14 40 26
rect 23 11 40 14
rect 23 9 25 11
rect 27 9 34 11
rect 36 10 40 11
rect 42 20 50 26
rect 42 18 45 20
rect 47 18 50 20
rect 42 10 50 18
rect 52 21 59 26
rect 52 19 55 21
rect 57 19 59 21
rect 52 14 59 19
rect 52 12 55 14
rect 57 12 59 14
rect 52 10 59 12
rect 36 9 38 10
rect 23 7 38 9
<< pdif >>
rect 13 68 22 70
rect 13 66 16 68
rect 18 66 22 68
rect 13 61 22 66
rect 2 59 9 61
rect 2 57 4 59
rect 6 57 9 59
rect 2 52 9 57
rect 2 50 4 52
rect 6 50 9 52
rect 2 48 9 50
rect 4 42 9 48
rect 11 44 22 61
rect 24 44 29 70
rect 31 44 36 70
rect 38 61 46 70
rect 38 59 41 61
rect 43 59 46 61
rect 38 44 46 59
rect 48 44 53 70
rect 55 44 60 70
rect 62 68 70 70
rect 62 66 65 68
rect 67 66 70 68
rect 62 61 70 66
rect 62 59 65 61
rect 67 59 70 61
rect 62 44 70 59
rect 11 42 16 44
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 61 47 62
rect 2 59 41 61
rect 43 59 47 61
rect 2 57 4 59
rect 6 58 47 59
rect 2 52 6 57
rect 2 50 4 52
rect 2 29 6 50
rect 10 50 23 54
rect 31 50 70 54
rect 10 37 14 50
rect 31 46 35 50
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 18 42 35 46
rect 41 42 55 46
rect 18 39 24 42
rect 18 37 21 39
rect 23 37 24 39
rect 18 33 24 37
rect 41 39 47 42
rect 41 37 42 39
rect 44 37 47 39
rect 30 33 34 35
rect 41 34 47 37
rect 65 39 70 50
rect 65 37 66 39
rect 68 37 70 39
rect 65 35 70 37
rect 30 31 31 33
rect 33 31 34 33
rect 30 30 34 31
rect 2 28 8 29
rect 2 26 4 28
rect 6 26 8 28
rect 2 21 8 26
rect 2 19 4 21
rect 6 19 8 21
rect 2 17 8 19
rect 30 26 70 30
rect 66 17 70 26
rect -2 11 74 12
rect -2 9 25 11
rect 27 9 34 11
rect 36 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 9 14 11 30
rect 19 14 21 30
rect 40 10 42 26
rect 50 10 52 26
<< pmos >>
rect 9 42 11 61
rect 22 44 24 70
rect 29 44 31 70
rect 36 44 38 70
rect 46 44 48 70
rect 53 44 55 70
rect 60 44 62 70
<< polyct0 >>
rect 52 31 54 33
<< polyct1 >>
rect 11 35 13 37
rect 21 37 23 39
rect 42 37 44 39
rect 66 37 68 39
rect 31 31 33 33
<< ndifct0 >>
rect 14 26 16 28
rect 14 19 16 21
rect 45 18 47 20
rect 55 19 57 21
rect 55 12 57 14
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
rect 25 9 27 11
rect 34 9 36 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 16 66 18 68
rect 65 66 67 68
rect 65 59 67 61
<< pdifct1 >>
rect 4 57 6 59
rect 4 50 6 52
rect 41 59 43 61
<< alu0 >>
rect 14 66 16 68
rect 18 66 20 68
rect 14 65 20 66
rect 63 66 65 68
rect 67 66 69 68
rect 63 61 69 66
rect 63 59 65 61
rect 67 59 69 61
rect 63 58 69 59
rect 6 48 7 58
rect 51 33 55 35
rect 51 31 52 33
rect 54 31 55 33
rect 51 30 55 31
rect 13 28 17 30
rect 13 26 14 28
rect 16 26 17 28
rect 13 21 17 26
rect 53 21 59 22
rect 13 19 14 21
rect 16 20 49 21
rect 16 19 45 20
rect 13 18 45 19
rect 47 18 49 20
rect 13 17 49 18
rect 53 19 55 21
rect 57 19 59 21
rect 53 14 59 19
rect 53 12 55 14
rect 57 12 59 14
<< labels >>
rlabel alu0 15 23 15 23 6 n3
rlabel alu0 31 19 31 19 6 n3
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 20 36 20 36 6 a1
rlabel alu1 20 52 20 52 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 28 44 28 44 6 a1
rlabel alu1 36 52 36 52 6 a1
rlabel alu1 28 60 28 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 52 28 52 28 6 a2
rlabel alu1 44 40 44 40 6 a3
rlabel alu1 52 44 52 44 6 a3
rlabel alu1 52 52 52 52 6 a1
rlabel alu1 44 52 44 52 6 a1
rlabel alu1 44 60 44 60 6 z
rlabel alu1 60 28 60 28 6 a2
rlabel alu1 68 20 68 20 6 a2
rlabel alu1 68 44 68 44 6 a1
rlabel alu1 60 52 60 52 6 a1
<< end >>
