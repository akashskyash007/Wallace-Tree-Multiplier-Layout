magic
tech scmos
timestamp 1199202168
<< ab >>
rect 0 0 200 80
<< nwell >>
rect -5 36 205 88
<< pwell >>
rect -5 -8 205 36
<< poly >>
rect 21 70 23 74
rect 31 70 33 74
rect 41 70 43 74
rect 51 70 53 74
rect 61 70 63 74
rect 71 70 73 74
rect 81 70 83 74
rect 91 70 93 74
rect 101 70 103 74
rect 108 70 110 74
rect 121 70 123 74
rect 128 70 130 74
rect 138 70 140 74
rect 145 70 147 74
rect 157 70 159 74
rect 167 70 169 74
rect 177 70 179 74
rect 10 50 12 55
rect 10 39 12 42
rect 21 39 23 42
rect 31 39 33 42
rect 10 37 33 39
rect 10 35 12 37
rect 14 35 19 37
rect 21 35 23 37
rect 10 33 23 35
rect 21 30 23 33
rect 31 30 33 37
rect 41 37 43 42
rect 51 37 53 42
rect 61 37 63 42
rect 41 35 63 37
rect 41 30 43 35
rect 51 30 53 35
rect 61 30 63 35
rect 71 39 73 42
rect 81 39 83 42
rect 91 39 93 42
rect 101 39 103 42
rect 71 37 93 39
rect 71 35 73 37
rect 75 35 83 37
rect 71 33 83 35
rect 71 30 73 33
rect 81 30 83 33
rect 91 30 93 37
rect 97 37 103 39
rect 97 35 99 37
rect 101 35 103 37
rect 97 33 103 35
rect 101 30 103 33
rect 108 39 110 42
rect 121 39 123 42
rect 108 37 123 39
rect 108 35 115 37
rect 117 35 123 37
rect 108 33 123 35
rect 108 30 110 33
rect 121 30 123 33
rect 128 39 130 42
rect 138 39 140 42
rect 128 37 140 39
rect 128 35 130 37
rect 132 35 140 37
rect 128 33 140 35
rect 128 30 130 33
rect 138 30 140 33
rect 145 39 147 42
rect 157 39 159 42
rect 167 39 169 42
rect 177 39 179 42
rect 145 37 179 39
rect 145 35 147 37
rect 149 35 160 37
rect 145 33 160 35
rect 145 30 147 33
rect 158 30 160 33
rect 168 30 170 37
rect 21 9 23 14
rect 31 9 33 14
rect 41 11 43 16
rect 51 11 53 16
rect 61 8 63 16
rect 71 12 73 16
rect 81 12 83 16
rect 91 12 93 16
rect 101 8 103 16
rect 108 11 110 16
rect 121 11 123 16
rect 128 11 130 16
rect 138 11 140 16
rect 145 11 147 16
rect 61 6 103 8
rect 158 6 160 10
rect 168 6 170 10
<< ndif >>
rect 14 27 21 30
rect 14 25 16 27
rect 18 25 21 27
rect 14 20 21 25
rect 14 18 16 20
rect 18 18 21 20
rect 14 14 21 18
rect 23 28 31 30
rect 23 26 26 28
rect 28 26 31 28
rect 23 21 31 26
rect 23 19 26 21
rect 28 19 31 21
rect 23 14 31 19
rect 33 27 41 30
rect 33 25 36 27
rect 38 25 41 27
rect 33 20 41 25
rect 33 18 36 20
rect 38 18 41 20
rect 33 16 41 18
rect 43 28 51 30
rect 43 26 46 28
rect 48 26 51 28
rect 43 21 51 26
rect 43 19 46 21
rect 48 19 51 21
rect 43 16 51 19
rect 53 20 61 30
rect 53 18 56 20
rect 58 18 61 20
rect 53 16 61 18
rect 63 28 71 30
rect 63 26 66 28
rect 68 26 71 28
rect 63 21 71 26
rect 63 19 66 21
rect 68 19 71 21
rect 63 16 71 19
rect 73 28 81 30
rect 73 26 76 28
rect 78 26 81 28
rect 73 16 81 26
rect 83 21 91 30
rect 83 19 86 21
rect 88 19 91 21
rect 83 16 91 19
rect 93 28 101 30
rect 93 26 96 28
rect 98 26 101 28
rect 93 16 101 26
rect 103 16 108 30
rect 110 16 121 30
rect 123 16 128 30
rect 130 28 138 30
rect 130 26 133 28
rect 135 26 138 28
rect 130 16 138 26
rect 140 16 145 30
rect 147 16 158 30
rect 33 14 39 16
rect 112 11 119 16
rect 149 14 158 16
rect 149 12 151 14
rect 153 12 158 14
rect 112 9 114 11
rect 116 9 119 11
rect 149 10 158 12
rect 160 28 168 30
rect 160 26 163 28
rect 165 26 168 28
rect 160 21 168 26
rect 160 19 163 21
rect 165 19 168 21
rect 160 10 168 19
rect 170 22 178 30
rect 170 20 173 22
rect 175 20 178 22
rect 170 14 178 20
rect 170 12 173 14
rect 175 12 178 14
rect 170 10 178 12
rect 112 7 119 9
<< pdif >>
rect 14 68 21 70
rect 14 66 16 68
rect 18 66 21 68
rect 14 61 21 66
rect 14 59 16 61
rect 18 59 21 61
rect 14 54 21 59
rect 14 52 16 54
rect 18 52 21 54
rect 14 50 21 52
rect 5 48 10 50
rect 3 46 10 48
rect 3 44 5 46
rect 7 44 10 46
rect 3 42 10 44
rect 12 42 21 50
rect 23 53 31 70
rect 23 51 26 53
rect 28 51 31 53
rect 23 46 31 51
rect 23 44 26 46
rect 28 44 31 46
rect 23 42 31 44
rect 33 68 41 70
rect 33 66 36 68
rect 38 66 41 68
rect 33 61 41 66
rect 33 59 36 61
rect 38 59 41 61
rect 33 54 41 59
rect 33 52 36 54
rect 38 52 41 54
rect 33 42 41 52
rect 43 54 51 70
rect 43 52 46 54
rect 48 52 51 54
rect 43 47 51 52
rect 43 45 46 47
rect 48 45 51 47
rect 43 42 51 45
rect 53 68 61 70
rect 53 66 56 68
rect 58 66 61 68
rect 53 61 61 66
rect 53 59 56 61
rect 58 59 61 61
rect 53 54 61 59
rect 53 52 56 54
rect 58 52 61 54
rect 53 42 61 52
rect 63 61 71 70
rect 63 59 66 61
rect 68 59 71 61
rect 63 54 71 59
rect 63 52 66 54
rect 68 52 71 54
rect 63 47 71 52
rect 63 45 66 47
rect 68 45 71 47
rect 63 42 71 45
rect 73 53 81 70
rect 73 51 76 53
rect 78 51 81 53
rect 73 46 81 51
rect 73 44 76 46
rect 78 44 81 46
rect 73 42 81 44
rect 83 61 91 70
rect 83 59 86 61
rect 88 59 91 61
rect 83 54 91 59
rect 83 52 86 54
rect 88 52 91 54
rect 83 42 91 52
rect 93 53 101 70
rect 93 51 96 53
rect 98 51 101 53
rect 93 46 101 51
rect 93 44 96 46
rect 98 44 101 46
rect 93 42 101 44
rect 103 42 108 70
rect 110 68 121 70
rect 110 66 114 68
rect 116 66 121 68
rect 110 42 121 66
rect 123 42 128 70
rect 130 53 138 70
rect 130 51 133 53
rect 135 51 138 53
rect 130 42 138 51
rect 140 42 145 70
rect 147 68 157 70
rect 147 66 151 68
rect 153 66 157 68
rect 147 42 157 66
rect 159 61 167 70
rect 159 59 162 61
rect 164 59 167 61
rect 159 54 167 59
rect 159 52 162 54
rect 164 52 167 54
rect 159 42 167 52
rect 169 68 177 70
rect 169 66 172 68
rect 174 66 177 68
rect 169 61 177 66
rect 169 59 172 61
rect 174 59 177 61
rect 169 42 177 59
rect 179 55 184 70
rect 179 53 186 55
rect 179 51 182 53
rect 184 51 186 53
rect 179 46 186 51
rect 179 44 182 46
rect 184 44 186 46
rect 179 42 186 44
<< alu1 >>
rect -2 81 202 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 202 81
rect -2 68 202 79
rect 74 53 79 55
rect 74 51 76 53
rect 78 51 79 53
rect 74 46 79 51
rect 94 53 158 54
rect 94 51 96 53
rect 98 51 133 53
rect 135 51 158 53
rect 94 50 158 51
rect 94 46 99 50
rect 74 44 76 46
rect 78 44 96 46
rect 98 44 99 46
rect 2 37 22 39
rect 2 35 12 37
rect 14 35 19 37
rect 21 35 22 37
rect 2 33 22 35
rect 74 42 99 44
rect 113 42 150 46
rect 2 25 6 33
rect 82 29 86 42
rect 97 37 109 38
rect 97 35 99 37
rect 101 35 109 37
rect 97 34 109 35
rect 113 37 119 42
rect 113 35 115 37
rect 117 35 119 37
rect 113 34 119 35
rect 123 37 135 38
rect 123 35 130 37
rect 132 35 135 37
rect 123 34 135 35
rect 146 37 150 42
rect 146 35 147 37
rect 149 35 150 37
rect 105 30 109 34
rect 123 30 127 34
rect 146 33 150 35
rect 74 28 100 29
rect 74 26 76 28
rect 78 26 96 28
rect 98 26 100 28
rect 105 26 127 30
rect 154 29 158 50
rect 131 28 158 29
rect 131 26 133 28
rect 135 26 158 28
rect 74 25 100 26
rect 131 25 158 26
rect -2 11 202 12
rect -2 9 114 11
rect 116 9 202 11
rect -2 1 202 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 202 1
rect -2 -2 202 -1
<< ptie >>
rect 0 1 200 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 200 1
rect 0 -3 200 -1
<< ntie >>
rect 0 81 200 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 200 81
rect 0 77 200 79
<< nmos >>
rect 21 14 23 30
rect 31 14 33 30
rect 41 16 43 30
rect 51 16 53 30
rect 61 16 63 30
rect 71 16 73 30
rect 81 16 83 30
rect 91 16 93 30
rect 101 16 103 30
rect 108 16 110 30
rect 121 16 123 30
rect 128 16 130 30
rect 138 16 140 30
rect 145 16 147 30
rect 158 10 160 30
rect 168 10 170 30
<< pmos >>
rect 10 42 12 50
rect 21 42 23 70
rect 31 42 33 70
rect 41 42 43 70
rect 51 42 53 70
rect 61 42 63 70
rect 71 42 73 70
rect 81 42 83 70
rect 91 42 93 70
rect 101 42 103 70
rect 108 42 110 70
rect 121 42 123 70
rect 128 42 130 70
rect 138 42 140 70
rect 145 42 147 70
rect 157 42 159 70
rect 167 42 169 70
rect 177 42 179 70
<< polyct0 >>
rect 73 35 75 37
<< polyct1 >>
rect 12 35 14 37
rect 19 35 21 37
rect 99 35 101 37
rect 115 35 117 37
rect 130 35 132 37
rect 147 35 149 37
<< ndifct0 >>
rect 16 25 18 27
rect 16 18 18 20
rect 26 26 28 28
rect 26 19 28 21
rect 36 25 38 27
rect 36 18 38 20
rect 46 26 48 28
rect 46 19 48 21
rect 56 18 58 20
rect 66 26 68 28
rect 66 19 68 21
rect 86 19 88 21
rect 151 12 153 14
rect 163 26 165 28
rect 163 19 165 21
rect 173 20 175 22
rect 173 12 175 14
<< ndifct1 >>
rect 76 26 78 28
rect 96 26 98 28
rect 133 26 135 28
rect 114 9 116 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
rect 171 79 173 81
rect 179 79 181 81
rect 187 79 189 81
rect 195 79 197 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
rect 171 -1 173 1
rect 179 -1 181 1
rect 187 -1 189 1
rect 195 -1 197 1
<< pdifct0 >>
rect 16 66 18 68
rect 16 59 18 61
rect 16 52 18 54
rect 5 44 7 46
rect 26 51 28 53
rect 26 44 28 46
rect 36 66 38 68
rect 36 59 38 61
rect 36 52 38 54
rect 46 52 48 54
rect 46 45 48 47
rect 56 66 58 68
rect 56 59 58 61
rect 56 52 58 54
rect 66 59 68 61
rect 66 52 68 54
rect 66 45 68 47
rect 86 59 88 61
rect 86 52 88 54
rect 114 66 116 68
rect 151 66 153 68
rect 162 59 164 61
rect 162 52 164 54
rect 172 66 174 68
rect 172 59 174 61
rect 182 51 184 53
rect 182 44 184 46
<< pdifct1 >>
rect 76 51 78 53
rect 76 44 78 46
rect 96 51 98 53
rect 96 44 98 46
rect 133 51 135 53
<< alu0 >>
rect 4 59 8 68
rect 15 66 16 68
rect 18 66 19 68
rect 15 61 19 66
rect 15 59 16 61
rect 18 59 19 61
rect 15 54 19 59
rect 35 66 36 68
rect 38 66 39 68
rect 35 61 39 66
rect 35 59 36 61
rect 38 59 39 61
rect 15 52 16 54
rect 18 52 19 54
rect 15 50 19 52
rect 25 53 29 55
rect 25 51 26 53
rect 28 51 29 53
rect 25 47 29 51
rect 35 54 39 59
rect 55 66 56 68
rect 58 66 59 68
rect 55 61 59 66
rect 112 66 114 68
rect 116 66 118 68
rect 112 65 118 66
rect 149 66 151 68
rect 153 66 155 68
rect 149 65 155 66
rect 170 66 172 68
rect 174 66 176 68
rect 55 59 56 61
rect 58 59 59 61
rect 35 52 36 54
rect 38 52 39 54
rect 35 50 39 52
rect 45 54 49 56
rect 45 52 46 54
rect 48 52 49 54
rect 3 46 29 47
rect 3 44 5 46
rect 7 44 26 46
rect 28 44 29 46
rect 3 43 29 44
rect 45 47 49 52
rect 55 54 59 59
rect 55 52 56 54
rect 58 52 59 54
rect 55 50 59 52
rect 64 61 166 62
rect 64 59 66 61
rect 68 59 86 61
rect 88 59 162 61
rect 164 59 166 61
rect 64 58 166 59
rect 170 61 176 66
rect 170 59 172 61
rect 174 59 176 61
rect 189 59 193 68
rect 170 58 176 59
rect 64 54 69 58
rect 64 52 66 54
rect 68 52 69 54
rect 64 47 69 52
rect 45 45 46 47
rect 48 45 66 47
rect 68 45 69 47
rect 45 43 69 45
rect 85 54 89 58
rect 161 54 166 58
rect 85 52 86 54
rect 88 52 89 54
rect 85 50 89 52
rect 161 52 162 54
rect 164 53 186 54
rect 164 52 182 53
rect 161 51 182 52
rect 184 51 186 53
rect 161 50 186 51
rect 25 38 29 43
rect 25 37 77 38
rect 25 35 73 37
rect 75 35 77 37
rect 25 34 77 35
rect 15 27 19 29
rect 15 25 16 27
rect 18 25 19 27
rect 4 12 8 21
rect 15 20 19 25
rect 15 18 16 20
rect 18 18 19 20
rect 15 12 19 18
rect 25 28 29 34
rect 25 26 26 28
rect 28 26 29 28
rect 25 21 29 26
rect 25 19 26 21
rect 28 19 29 21
rect 25 17 29 19
rect 35 27 39 29
rect 35 25 36 27
rect 38 25 39 27
rect 35 20 39 25
rect 35 18 36 20
rect 38 18 39 20
rect 35 12 39 18
rect 45 28 69 30
rect 45 26 46 28
rect 48 26 66 28
rect 68 26 69 28
rect 45 21 49 26
rect 64 22 69 26
rect 180 46 186 50
rect 180 44 182 46
rect 184 44 186 46
rect 180 43 186 44
rect 162 28 167 30
rect 162 26 163 28
rect 165 26 167 28
rect 162 22 167 26
rect 45 19 46 21
rect 48 19 49 21
rect 45 17 49 19
rect 55 20 59 22
rect 55 18 56 20
rect 58 18 59 20
rect 64 21 167 22
rect 64 19 66 21
rect 68 19 86 21
rect 88 19 163 21
rect 165 19 167 21
rect 64 18 167 19
rect 172 22 176 24
rect 172 20 173 22
rect 175 20 176 22
rect 55 12 59 18
rect 149 14 155 15
rect 149 12 151 14
rect 153 12 155 14
rect 172 14 176 20
rect 172 12 173 14
rect 175 12 176 14
rect 186 12 190 21
<< labels >>
rlabel alu0 47 23 47 23 6 n3
rlabel alu0 66 24 66 24 6 n3
rlabel alu0 66 52 66 52 6 n1
rlabel alu0 47 49 47 49 6 n1
rlabel alu0 87 56 87 56 6 n1
rlabel alu0 115 20 115 20 6 n3
rlabel alu0 164 24 164 24 6 n3
rlabel alu0 183 48 183 48 6 n1
rlabel alu0 163 56 163 56 6 n1
rlabel alu0 173 52 173 52 6 n1
rlabel alu1 4 32 4 32 6 c
rlabel alu1 12 36 12 36 6 c
rlabel polyct1 20 36 20 36 6 c
rlabel alu1 76 52 76 52 6 z
rlabel alu1 100 6 100 6 6 vss
rlabel alu1 108 28 108 28 6 b
rlabel alu1 116 28 116 28 6 b
rlabel alu1 116 40 116 40 6 a
rlabel alu1 92 44 92 44 6 z
rlabel polyct1 100 36 100 36 6 b
rlabel alu1 84 36 84 36 6 z
rlabel alu1 116 52 116 52 6 z
rlabel alu1 100 52 100 52 6 z
rlabel alu1 108 52 108 52 6 z
rlabel alu1 100 74 100 74 6 vdd
rlabel alu1 124 28 124 28 6 b
rlabel alu1 124 44 124 44 6 a
rlabel polyct1 148 36 148 36 6 a
rlabel alu1 132 36 132 36 6 b
rlabel alu1 132 44 132 44 6 a
rlabel alu1 140 44 140 44 6 a
rlabel alu1 156 36 156 36 6 z
rlabel alu1 140 52 140 52 6 z
rlabel alu1 148 52 148 52 6 z
rlabel alu1 132 52 132 52 6 z
rlabel alu1 124 52 124 52 6 z
<< end >>
