magic
tech scmos
timestamp 1199980631
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -8 40 104 97
<< pwell >>
rect -8 -9 104 40
<< poly >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 69 84 78 86
rect 69 82 74 84
rect 76 82 78 84
rect 69 80 78 82
rect 82 84 91 86
rect 82 82 84 84
rect 86 82 91 84
rect 82 80 91 82
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 66 46 75 48
rect 66 44 71 46
rect 73 44 75 46
rect 66 42 75 44
rect 79 46 94 48
rect 79 44 87 46
rect 89 44 94 46
rect 79 42 94 44
rect 2 36 17 38
rect 2 34 7 36
rect 9 34 17 36
rect 2 32 17 34
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 66 36 81 38
rect 66 34 71 36
rect 73 34 81 36
rect 66 32 81 34
rect 85 36 94 38
rect 85 34 87 36
rect 89 34 94 36
rect 85 32 94 34
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 2 14 8
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
rect 69 2 78 8
rect 82 2 91 8
<< ndif >>
rect 2 23 9 29
rect 2 21 4 23
rect 6 21 9 23
rect 2 16 9 21
rect 2 14 4 16
rect 6 14 9 16
rect 2 11 9 14
rect 11 25 21 29
rect 11 23 15 25
rect 17 23 21 25
rect 11 17 21 23
rect 11 15 15 17
rect 17 15 21 17
rect 11 11 21 15
rect 23 15 30 29
rect 23 13 26 15
rect 28 13 30 15
rect 23 11 30 13
rect 34 15 41 29
rect 34 13 36 15
rect 38 13 41 15
rect 34 11 41 13
rect 43 25 53 29
rect 43 23 47 25
rect 49 23 53 25
rect 43 17 53 23
rect 43 15 47 17
rect 49 15 53 17
rect 43 11 53 15
rect 55 15 62 29
rect 55 13 58 15
rect 60 13 62 15
rect 55 11 62 13
rect 66 15 73 29
rect 66 13 68 15
rect 70 13 73 15
rect 66 11 73 13
rect 75 11 85 29
rect 87 23 94 29
rect 87 21 90 23
rect 92 21 94 23
rect 87 16 94 21
rect 87 14 90 16
rect 92 14 94 16
rect 87 11 94 14
<< pdif >>
rect 2 74 9 77
rect 2 72 4 74
rect 6 72 9 74
rect 2 67 9 72
rect 2 65 4 67
rect 6 65 9 67
rect 2 51 9 65
rect 11 65 21 77
rect 11 63 15 65
rect 17 63 21 65
rect 11 57 21 63
rect 11 55 15 57
rect 17 55 21 57
rect 11 51 21 55
rect 23 74 30 77
rect 23 72 26 74
rect 28 72 30 74
rect 23 67 30 72
rect 23 65 26 67
rect 28 65 30 67
rect 23 51 30 65
rect 34 74 41 77
rect 34 72 36 74
rect 38 72 41 74
rect 34 67 41 72
rect 34 65 36 67
rect 38 65 41 67
rect 34 51 41 65
rect 43 65 53 77
rect 43 63 47 65
rect 49 63 53 65
rect 43 57 53 63
rect 43 55 47 57
rect 49 55 53 57
rect 43 51 53 55
rect 55 74 62 77
rect 55 72 58 74
rect 60 72 62 74
rect 55 67 62 72
rect 55 65 58 67
rect 60 65 62 67
rect 55 51 62 65
rect 66 74 73 77
rect 66 72 68 74
rect 70 72 73 74
rect 66 67 73 72
rect 66 65 68 67
rect 70 65 73 67
rect 66 51 73 65
rect 75 65 85 77
rect 75 63 79 65
rect 81 63 85 65
rect 75 51 85 63
rect 87 74 94 77
rect 87 72 90 74
rect 92 72 94 74
rect 87 67 94 72
rect 87 65 90 67
rect 92 65 94 67
rect 87 51 94 65
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 83 7 85
rect -2 81 7 83
rect 3 74 7 81
rect 30 83 31 85
rect 33 83 34 85
rect 30 76 34 83
rect 62 85 66 90
rect 62 83 63 85
rect 65 83 66 85
rect 62 76 66 83
rect 94 85 98 90
rect 90 83 95 85
rect 97 83 98 85
rect 90 81 98 83
rect 90 76 94 81
rect 3 72 4 74
rect 6 72 7 74
rect 3 67 7 72
rect 25 74 39 76
rect 25 72 26 74
rect 28 72 36 74
rect 38 72 39 74
rect 25 67 29 72
rect 3 65 4 67
rect 6 65 7 67
rect 3 63 7 65
rect 13 65 18 67
rect 13 63 15 65
rect 17 63 18 65
rect 25 65 26 67
rect 28 65 29 67
rect 25 63 29 65
rect 35 67 39 72
rect 57 74 71 76
rect 57 72 58 74
rect 60 72 68 74
rect 70 72 71 74
rect 57 67 61 72
rect 35 65 36 67
rect 38 65 39 67
rect 35 63 39 65
rect 46 65 50 67
rect 46 63 47 65
rect 49 63 50 65
rect 57 65 58 67
rect 60 65 61 67
rect 57 63 61 65
rect 67 67 71 72
rect 89 74 94 76
rect 89 72 90 74
rect 92 72 94 74
rect 89 67 94 72
rect 67 65 68 67
rect 70 65 71 67
rect 67 63 71 65
rect 78 65 82 67
rect 78 63 79 65
rect 81 63 82 65
rect 89 65 90 67
rect 92 65 94 67
rect 89 63 94 65
rect 13 58 18 63
rect 46 58 50 63
rect 78 58 82 63
rect 13 57 82 58
rect 13 55 15 57
rect 17 55 47 57
rect 49 55 82 57
rect 13 54 82 55
rect 5 46 11 48
rect 5 44 7 46
rect 9 44 11 46
rect 5 42 11 44
rect 21 46 27 50
rect 21 44 23 46
rect 25 44 27 46
rect 21 42 27 44
rect 38 46 42 48
rect 38 44 39 46
rect 41 44 42 46
rect 38 42 42 44
rect 54 46 58 48
rect 54 44 55 46
rect 57 44 58 46
rect 54 42 58 44
rect 70 46 74 48
rect 70 44 71 46
rect 73 44 74 46
rect 70 42 74 44
rect 5 38 74 42
rect 5 36 11 38
rect 5 34 7 36
rect 9 34 11 36
rect 5 30 11 34
rect 21 36 27 38
rect 21 34 23 36
rect 25 34 27 36
rect 21 33 27 34
rect 38 36 42 38
rect 38 34 39 36
rect 41 34 42 36
rect 38 32 42 34
rect 54 36 58 38
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 70 36 74 38
rect 70 34 71 36
rect 73 34 74 36
rect 70 32 74 34
rect 78 26 82 54
rect 13 25 82 26
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 16 7 21
rect 3 14 4 16
rect 6 14 7 16
rect 3 7 7 14
rect 13 23 15 25
rect 17 23 47 25
rect 49 23 82 25
rect 13 22 82 23
rect 13 17 18 22
rect 13 15 15 17
rect 17 15 18 17
rect 46 17 50 22
rect 13 13 18 15
rect 24 15 40 16
rect 24 13 26 15
rect 28 13 36 15
rect 38 13 40 15
rect 46 15 47 17
rect 49 15 50 17
rect 46 13 50 15
rect 56 15 72 16
rect 56 13 58 15
rect 60 13 68 15
rect 70 13 72 15
rect 78 13 82 22
rect 89 23 93 25
rect 89 21 90 23
rect 92 21 93 23
rect 89 16 93 21
rect 89 14 90 16
rect 92 14 93 16
rect 24 12 40 13
rect 56 12 72 13
rect -2 5 7 7
rect -2 3 -1 5
rect 1 3 7 5
rect 30 5 34 12
rect 30 3 31 5
rect 33 3 34 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 5 66 12
rect 62 3 63 5
rect 65 3 66 5
rect 89 7 93 14
rect 89 5 98 7
rect 89 3 95 5
rect 97 3 98 5
rect 62 -2 66 3
rect 94 -2 98 3
<< alu2 >>
rect -2 85 98 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 95 85
rect 97 83 98 85
rect -2 80 98 83
rect -2 5 98 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 95 5
rect 97 3 98 5
rect -2 -2 98 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
rect 93 5 99 7
rect 93 3 95 5
rect 97 3 99 5
rect 93 0 99 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
rect 93 85 99 88
rect 93 83 95 85
rect 97 83 99 85
rect 93 81 99 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polyct0 >>
rect 74 82 76 84
rect 84 82 86 84
rect 87 44 89 46
rect 87 34 89 36
<< polyct1 >>
rect 7 44 9 46
rect 23 44 25 46
rect 39 44 41 46
rect 55 44 57 46
rect 71 44 73 46
rect 7 34 9 36
rect 23 34 25 36
rect 39 34 41 36
rect 55 34 57 36
rect 71 34 73 36
<< ndifct1 >>
rect 4 21 6 23
rect 4 14 6 16
rect 15 23 17 25
rect 15 15 17 17
rect 26 13 28 15
rect 36 13 38 15
rect 47 23 49 25
rect 47 15 49 17
rect 58 13 60 15
rect 68 13 70 15
rect 90 21 92 23
rect 90 14 92 16
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< pdifct1 >>
rect 4 72 6 74
rect 4 65 6 67
rect 15 63 17 65
rect 15 55 17 57
rect 26 72 28 74
rect 26 65 28 67
rect 36 72 38 74
rect 36 65 38 67
rect 47 63 49 65
rect 47 55 49 57
rect 58 72 60 74
rect 58 65 60 67
rect 68 72 70 74
rect 68 65 70 67
rect 79 63 81 65
rect 90 72 92 74
rect 90 65 92 67
<< alu0 >>
rect 73 84 87 86
rect 73 82 74 84
rect 76 82 84 84
rect 86 82 87 84
rect 73 80 87 82
rect 86 46 90 48
rect 86 44 87 46
rect 89 44 90 46
rect 86 36 90 44
rect 86 34 87 36
rect 89 34 90 36
rect 86 32 90 34
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< labels >>
rlabel alu1 8 36 8 36 6 a
rlabel alu1 16 20 16 20 6 z
rlabel alu1 32 24 32 24 6 z
rlabel alu1 24 24 24 24 6 z
rlabel alu1 16 40 16 40 6 a
rlabel alu1 32 40 32 40 6 a
rlabel alu1 24 44 24 44 6 a
rlabel alu1 24 56 24 56 6 z
rlabel alu1 32 56 32 56 6 z
rlabel alu1 16 60 16 60 6 z
rlabel alu1 40 24 40 24 6 z
rlabel alu1 56 24 56 24 6 z
rlabel alu1 40 40 40 40 6 a
rlabel alu1 56 40 56 40 6 a
rlabel alu1 48 40 48 40 6 a
rlabel alu1 56 56 56 56 6 z
rlabel alu1 40 56 40 56 6 z
rlabel alu1 72 24 72 24 6 z
rlabel alu1 64 24 64 24 6 z
rlabel alu1 72 40 72 40 6 a
rlabel alu1 64 40 64 40 6 a
rlabel alu1 64 56 64 56 6 z
rlabel alu1 72 56 72 56 6 z
rlabel alu1 80 40 80 40 6 z
rlabel alu2 48 4 48 4 6 vss
rlabel alu2 48 84 48 84 6 vdd
<< end >>
