magic
tech scmos
timestamp 1199201893
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 9 47 11 50
rect 9 45 15 47
rect 9 43 11 45
rect 13 43 15 45
rect 9 41 15 43
rect 19 37 21 50
rect 29 44 31 50
rect 14 35 21 37
rect 25 42 31 44
rect 39 47 41 50
rect 39 45 47 47
rect 39 43 43 45
rect 45 43 47 45
rect 14 31 16 35
rect 25 31 27 42
rect 39 41 47 43
rect 39 37 41 41
rect 9 29 16 31
rect 9 27 11 29
rect 13 27 16 29
rect 9 25 16 27
rect 14 22 16 25
rect 21 29 27 31
rect 21 27 23 29
rect 25 27 27 29
rect 21 25 27 27
rect 31 35 41 37
rect 21 22 23 25
rect 31 22 33 35
rect 38 29 47 31
rect 38 27 43 29
rect 45 27 47 29
rect 38 25 47 27
rect 38 22 40 25
rect 14 10 16 15
rect 21 10 23 15
rect 31 10 33 15
rect 38 10 40 15
<< ndif >>
rect 5 15 14 22
rect 16 15 21 22
rect 23 20 31 22
rect 23 18 26 20
rect 28 18 31 20
rect 23 15 31 18
rect 33 15 38 22
rect 40 19 48 22
rect 40 17 44 19
rect 46 17 48 19
rect 40 15 48 17
rect 5 11 12 15
rect 5 9 8 11
rect 10 9 12 11
rect 5 7 12 9
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 50 9 62
rect 11 62 19 66
rect 11 60 14 62
rect 16 60 19 62
rect 11 50 19 60
rect 21 54 29 66
rect 21 52 24 54
rect 26 52 29 54
rect 21 50 29 52
rect 31 62 39 66
rect 31 60 34 62
rect 36 60 39 62
rect 31 50 39 60
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 50 49 62
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 22 54 28 55
rect 2 52 24 54
rect 26 52 28 54
rect 2 50 28 52
rect 33 50 47 54
rect 2 21 6 50
rect 11 45 34 46
rect 13 43 34 45
rect 11 42 34 43
rect 41 45 47 50
rect 41 43 43 45
rect 45 43 47 45
rect 41 42 47 43
rect 30 38 34 42
rect 10 34 23 38
rect 30 34 46 38
rect 10 29 14 34
rect 10 27 11 29
rect 13 27 14 29
rect 10 25 14 27
rect 21 29 38 30
rect 21 27 23 29
rect 25 27 38 29
rect 21 26 38 27
rect 2 20 30 21
rect 2 18 26 20
rect 28 18 30 20
rect 2 17 30 18
rect 34 17 38 26
rect 42 29 46 34
rect 42 27 43 29
rect 45 27 46 29
rect 42 25 46 27
rect -2 11 58 12
rect -2 9 8 11
rect 10 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 14 15 16 22
rect 21 15 23 22
rect 31 15 33 22
rect 38 15 40 22
<< pmos >>
rect 9 50 11 66
rect 19 50 21 66
rect 29 50 31 66
rect 39 50 41 66
<< polyct1 >>
rect 11 43 13 45
rect 43 43 45 45
rect 11 27 13 29
rect 23 27 25 29
rect 43 27 45 29
<< ndifct0 >>
rect 44 17 46 19
<< ndifct1 >>
rect 26 18 28 20
rect 8 9 10 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 62 6 64
rect 14 60 16 62
rect 34 60 36 62
rect 44 62 46 64
<< pdifct1 >>
rect 24 52 26 54
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 43 64 47 68
rect 3 60 7 62
rect 12 62 38 63
rect 12 60 14 62
rect 16 60 34 62
rect 36 60 38 62
rect 43 62 44 64
rect 46 62 47 64
rect 43 60 47 62
rect 12 59 38 60
rect 10 46 14 47
rect 10 42 11 46
rect 10 41 30 42
rect 43 19 47 21
rect 43 17 44 19
rect 46 17 47 19
rect 43 12 47 17
<< labels >>
rlabel alu0 25 61 25 61 6 n3
rlabel alu1 4 32 4 32 6 z
rlabel polyct1 12 28 12 28 6 b1
rlabel alu1 20 36 20 36 6 b1
rlabel alu1 20 44 20 44 6 a1
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 20 36 20 6 b2
rlabel alu1 28 28 28 28 6 b2
rlabel alu1 36 36 36 36 6 a1
rlabel alu1 28 44 28 44 6 a1
rlabel alu1 36 52 36 52 6 a2
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 28 44 28 6 a1
rlabel alu1 44 48 44 48 6 a2
<< end >>
