magic
tech scmos
timestamp 1199202794
<< ab >>
rect 0 0 136 72
<< nwell >>
rect -5 32 141 77
<< pwell >>
rect -5 -5 141 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 99 66 101 70
rect 109 66 111 70
rect 119 57 121 61
rect 9 35 11 44
rect 19 43 21 46
rect 19 41 25 43
rect 19 39 21 41
rect 23 39 25 41
rect 19 37 25 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 32 15 33
rect 13 31 17 32
rect 9 29 17 31
rect 15 26 17 29
rect 22 26 24 37
rect 29 35 31 46
rect 39 35 41 46
rect 49 43 51 46
rect 45 41 51 43
rect 45 39 47 41
rect 49 39 51 41
rect 45 37 51 39
rect 29 33 41 35
rect 29 31 37 33
rect 39 31 41 33
rect 29 29 41 31
rect 29 26 31 29
rect 39 26 41 29
rect 46 26 48 37
rect 59 31 61 46
rect 69 31 71 46
rect 79 43 81 46
rect 79 41 85 43
rect 79 39 81 41
rect 83 39 85 41
rect 79 37 85 39
rect 53 29 77 31
rect 53 26 55 29
rect 62 25 68 29
rect 75 26 77 29
rect 82 26 84 37
rect 89 35 91 46
rect 99 35 101 46
rect 109 42 111 46
rect 105 40 111 42
rect 105 38 107 40
rect 109 38 111 40
rect 105 36 111 38
rect 89 33 101 35
rect 89 31 92 33
rect 94 31 101 33
rect 89 29 101 31
rect 89 26 91 29
rect 99 26 101 29
rect 106 26 108 36
rect 119 35 121 39
rect 119 33 127 35
rect 119 31 123 33
rect 125 31 127 33
rect 113 29 127 31
rect 113 26 115 29
rect 62 23 64 25
rect 66 23 68 25
rect 62 21 68 23
rect 15 2 17 6
rect 22 2 24 6
rect 29 2 31 6
rect 39 2 41 6
rect 46 2 48 6
rect 53 2 55 6
rect 75 2 77 6
rect 82 2 84 6
rect 89 2 91 6
rect 99 2 101 6
rect 106 2 108 6
rect 113 2 115 6
<< ndif >>
rect 7 10 15 26
rect 7 8 10 10
rect 12 8 15 10
rect 7 6 15 8
rect 17 6 22 26
rect 24 6 29 26
rect 31 17 39 26
rect 31 15 34 17
rect 36 15 39 17
rect 31 6 39 15
rect 41 6 46 26
rect 48 6 53 26
rect 55 18 60 26
rect 70 18 75 26
rect 55 10 75 18
rect 55 8 58 10
rect 60 8 70 10
rect 72 8 75 10
rect 55 6 75 8
rect 77 6 82 26
rect 84 6 89 26
rect 91 17 99 26
rect 91 15 94 17
rect 96 15 99 17
rect 91 6 99 15
rect 101 6 106 26
rect 108 6 113 26
rect 115 17 123 26
rect 115 15 118 17
rect 120 15 123 17
rect 115 10 123 15
rect 115 8 118 10
rect 120 8 123 10
rect 115 6 123 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 44 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 46 19 48
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 46 29 55
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 50 39 55
rect 31 48 34 50
rect 36 48 39 50
rect 31 46 39 48
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 46 49 55
rect 51 57 59 66
rect 51 55 54 57
rect 56 55 59 57
rect 51 50 59 55
rect 51 48 54 50
rect 56 48 59 50
rect 51 46 59 48
rect 61 64 69 66
rect 61 62 64 64
rect 66 62 69 64
rect 61 57 69 62
rect 61 55 64 57
rect 66 55 69 57
rect 61 46 69 55
rect 71 57 79 66
rect 71 55 74 57
rect 76 55 79 57
rect 71 50 79 55
rect 71 48 74 50
rect 76 48 79 50
rect 71 46 79 48
rect 81 64 89 66
rect 81 62 84 64
rect 86 62 89 64
rect 81 57 89 62
rect 81 55 84 57
rect 86 55 89 57
rect 81 46 89 55
rect 91 57 99 66
rect 91 55 94 57
rect 96 55 99 57
rect 91 50 99 55
rect 91 48 94 50
rect 96 48 99 50
rect 91 46 99 48
rect 101 64 109 66
rect 101 62 104 64
rect 106 62 109 64
rect 101 57 109 62
rect 101 55 104 57
rect 106 55 109 57
rect 101 46 109 55
rect 111 57 116 66
rect 111 53 119 57
rect 111 51 114 53
rect 116 51 119 53
rect 111 46 119 51
rect 11 44 16 46
rect 114 39 119 46
rect 121 55 129 57
rect 121 53 125 55
rect 127 53 129 55
rect 121 48 129 53
rect 121 46 125 48
rect 127 46 129 48
rect 121 39 129 46
<< alu1 >>
rect -2 67 138 72
rect -2 65 126 67
rect 128 65 138 67
rect -2 64 138 65
rect 33 57 38 59
rect 33 55 34 57
rect 36 55 38 57
rect 33 50 38 55
rect 73 57 78 59
rect 73 55 74 57
rect 76 55 78 57
rect 73 50 78 55
rect 113 53 119 59
rect 113 51 114 53
rect 116 51 119 53
rect 113 50 119 51
rect 2 48 14 50
rect 16 48 34 50
rect 36 48 54 50
rect 56 48 74 50
rect 76 48 94 50
rect 96 48 119 50
rect 2 46 119 48
rect 2 18 6 46
rect 19 41 119 42
rect 19 39 21 41
rect 23 39 47 41
rect 49 39 81 41
rect 83 40 119 41
rect 83 39 107 40
rect 19 38 107 39
rect 109 38 119 40
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 33 33 96 34
rect 33 31 37 33
rect 39 31 92 33
rect 94 31 96 33
rect 33 30 96 31
rect 105 30 111 38
rect 121 33 127 34
rect 121 31 123 33
rect 125 31 127 33
rect 121 26 127 31
rect 10 25 127 26
rect 10 23 64 25
rect 66 23 127 25
rect 10 22 127 23
rect 2 17 103 18
rect 2 15 34 17
rect 36 15 94 17
rect 96 15 103 17
rect 2 14 103 15
rect -2 7 138 8
rect -2 5 129 7
rect 131 5 138 7
rect -2 0 138 5
<< ptie >>
rect 127 7 133 24
rect 127 5 129 7
rect 131 5 133 7
rect 127 3 133 5
<< ntie >>
rect 121 67 133 69
rect 121 65 126 67
rect 128 65 133 67
rect 121 63 133 65
<< nmos >>
rect 15 6 17 26
rect 22 6 24 26
rect 29 6 31 26
rect 39 6 41 26
rect 46 6 48 26
rect 53 6 55 26
rect 75 6 77 26
rect 82 6 84 26
rect 89 6 91 26
rect 99 6 101 26
rect 106 6 108 26
rect 113 6 115 26
<< pmos >>
rect 9 44 11 66
rect 19 46 21 66
rect 29 46 31 66
rect 39 46 41 66
rect 49 46 51 66
rect 59 46 61 66
rect 69 46 71 66
rect 79 46 81 66
rect 89 46 91 66
rect 99 46 101 66
rect 109 46 111 66
rect 119 39 121 57
<< polyct1 >>
rect 21 39 23 41
rect 11 31 13 33
rect 47 39 49 41
rect 37 31 39 33
rect 81 39 83 41
rect 107 38 109 40
rect 92 31 94 33
rect 123 31 125 33
rect 64 23 66 25
<< ndifct0 >>
rect 10 8 12 10
rect 58 8 60 10
rect 70 8 72 10
rect 118 15 120 17
rect 118 8 120 10
<< ndifct1 >>
rect 34 15 36 17
rect 94 15 96 17
<< ntiect1 >>
rect 126 65 128 67
<< ptiect1 >>
rect 129 5 131 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 55 16 57
rect 24 62 26 64
rect 24 55 26 57
rect 44 62 46 64
rect 44 55 46 57
rect 54 55 56 57
rect 64 62 66 64
rect 64 55 66 57
rect 84 62 86 64
rect 84 55 86 57
rect 94 55 96 57
rect 104 62 106 64
rect 104 55 106 57
rect 125 53 127 55
rect 125 46 127 48
<< pdifct1 >>
rect 14 48 16 50
rect 34 55 36 57
rect 34 48 36 50
rect 54 48 56 50
rect 74 55 76 57
rect 74 48 76 50
rect 94 48 96 50
rect 114 51 116 53
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 50 17 55
rect 22 57 28 62
rect 42 62 44 64
rect 46 62 48 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 42 57 48 62
rect 62 62 64 64
rect 66 62 68 64
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 53 57 57 59
rect 53 55 54 57
rect 56 55 57 57
rect 53 50 57 55
rect 62 57 68 62
rect 82 62 84 64
rect 86 62 88 64
rect 62 55 64 57
rect 66 55 68 57
rect 62 54 68 55
rect 82 57 88 62
rect 102 62 104 64
rect 106 62 108 64
rect 82 55 84 57
rect 86 55 88 57
rect 82 54 88 55
rect 93 57 97 59
rect 93 55 94 57
rect 96 55 97 57
rect 93 50 97 55
rect 102 57 108 62
rect 102 55 104 57
rect 106 55 108 57
rect 102 54 108 55
rect 123 55 129 64
rect 123 53 125 55
rect 127 53 129 55
rect 123 48 129 53
rect 123 46 125 48
rect 127 46 129 48
rect 123 45 129 46
rect 116 17 122 18
rect 116 15 118 17
rect 120 15 122 17
rect 8 10 14 11
rect 8 8 10 10
rect 12 8 14 10
rect 56 10 62 11
rect 56 8 58 10
rect 60 8 62 10
rect 68 10 74 11
rect 68 8 70 10
rect 72 8 74 10
rect 116 10 122 15
rect 116 8 118 10
rect 120 8 122 10
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 24 20 24 6 a
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 28 24 28 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 36 24 36 24 6 a
rlabel alu1 36 32 36 32 6 c
rlabel alu1 44 32 44 32 6 c
rlabel alu1 28 40 28 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 68 4 68 4 6 vss
rlabel alu1 60 16 60 16 6 z
rlabel alu1 68 16 68 16 6 z
rlabel alu1 76 16 76 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 52 24 52 24 6 a
rlabel alu1 68 24 68 24 6 a
rlabel alu1 76 24 76 24 6 a
rlabel alu1 60 24 60 24 6 a
rlabel alu1 60 32 60 32 6 c
rlabel alu1 68 32 68 32 6 c
rlabel alu1 76 32 76 32 6 c
rlabel alu1 52 32 52 32 6 c
rlabel alu1 52 40 52 40 6 b
rlabel alu1 68 40 68 40 6 b
rlabel alu1 76 40 76 40 6 b
rlabel alu1 60 40 60 40 6 b
rlabel alu1 52 48 52 48 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 68 68 68 68 6 vdd
rlabel alu1 92 16 92 16 6 z
rlabel alu1 100 16 100 16 6 z
rlabel alu1 84 16 84 16 6 z
rlabel alu1 84 24 84 24 6 a
rlabel alu1 92 24 92 24 6 a
rlabel alu1 108 24 108 24 6 a
rlabel alu1 100 24 100 24 6 a
rlabel alu1 92 32 92 32 6 c
rlabel alu1 84 32 84 32 6 c
rlabel alu1 84 40 84 40 6 b
rlabel alu1 92 40 92 40 6 b
rlabel alu1 108 36 108 36 6 b
rlabel alu1 100 40 100 40 6 b
rlabel alu1 84 48 84 48 6 z
rlabel alu1 92 48 92 48 6 z
rlabel alu1 108 48 108 48 6 z
rlabel alu1 100 48 100 48 6 z
rlabel alu1 116 24 116 24 6 a
rlabel alu1 124 28 124 28 6 a
rlabel alu1 116 40 116 40 6 b
rlabel alu1 116 52 116 52 6 z
<< end >>
