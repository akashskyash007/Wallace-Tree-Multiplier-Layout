magic
tech scmos
timestamp 1199543659
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -5 48 105 105
<< pwell >>
rect -5 -5 105 48
<< poly >>
rect 35 94 37 98
rect 47 94 49 98
rect 57 94 59 98
rect 81 94 83 98
rect 11 84 13 88
rect 23 85 25 89
rect 11 43 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 21 51 25 53
rect 33 51 37 53
rect 21 43 23 51
rect 33 43 35 51
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 35 43
rect 27 39 29 41
rect 31 39 35 41
rect 47 43 49 55
rect 57 43 59 55
rect 81 53 83 56
rect 75 51 83 53
rect 75 49 77 51
rect 79 49 83 51
rect 75 47 83 49
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 27 37 35 39
rect 11 34 13 37
rect 21 34 23 37
rect 33 34 35 37
rect 45 37 53 39
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 45 34 47 37
rect 57 34 59 37
rect 81 35 83 47
rect 33 18 35 22
rect 45 18 47 22
rect 11 12 13 16
rect 21 13 23 17
rect 57 18 59 22
rect 81 11 83 15
<< ndif >>
rect 3 16 11 34
rect 13 17 21 34
rect 23 22 33 34
rect 35 22 45 34
rect 47 22 57 34
rect 59 22 67 34
rect 23 21 31 22
rect 23 19 27 21
rect 29 19 31 21
rect 23 17 31 19
rect 37 21 43 22
rect 37 19 39 21
rect 41 19 43 21
rect 37 17 43 19
rect 13 16 18 17
rect 3 11 9 16
rect 49 11 55 22
rect 61 21 67 22
rect 61 19 63 21
rect 65 19 67 21
rect 61 17 67 19
rect 73 31 81 35
rect 73 29 75 31
rect 77 29 81 31
rect 73 21 81 29
rect 73 19 75 21
rect 77 19 81 21
rect 73 15 81 19
rect 83 31 91 35
rect 83 29 87 31
rect 89 29 91 31
rect 83 21 91 29
rect 83 19 87 21
rect 89 19 91 21
rect 83 15 91 19
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 28 85 35 94
rect 15 84 23 85
rect 3 81 11 84
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 56 23 84
rect 25 81 35 85
rect 25 79 29 81
rect 31 79 35 81
rect 25 56 35 79
rect 37 71 47 94
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 13 55 18 56
rect 42 55 47 56
rect 49 55 57 94
rect 59 81 67 94
rect 59 79 63 81
rect 65 79 67 81
rect 59 55 67 79
rect 73 91 81 94
rect 73 89 75 91
rect 77 89 81 91
rect 73 81 81 89
rect 73 79 75 81
rect 77 79 81 81
rect 73 56 81 79
rect 83 81 91 94
rect 83 79 87 81
rect 89 79 91 81
rect 83 71 91 79
rect 83 69 87 71
rect 89 69 91 71
rect 83 61 91 69
rect 83 59 87 61
rect 89 59 91 61
rect 83 56 91 59
<< alu1 >>
rect -2 91 102 100
rect -2 89 17 91
rect 19 89 75 91
rect 77 89 102 91
rect -2 88 102 89
rect 3 81 67 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 79 63 81
rect 65 79 67 81
rect 3 78 67 79
rect 74 81 78 88
rect 88 82 92 83
rect 74 79 75 81
rect 77 79 78 81
rect 74 77 78 79
rect 85 81 92 82
rect 85 79 87 81
rect 89 79 92 81
rect 85 78 92 79
rect 8 41 12 73
rect 8 39 9 41
rect 11 39 12 41
rect 8 17 12 39
rect 18 41 22 73
rect 18 39 19 41
rect 21 39 22 41
rect 18 27 22 39
rect 28 41 32 73
rect 88 72 92 78
rect 28 39 29 41
rect 31 39 32 41
rect 28 37 32 39
rect 38 71 80 72
rect 38 69 41 71
rect 43 69 80 71
rect 38 68 80 69
rect 85 71 92 72
rect 85 69 87 71
rect 89 69 92 71
rect 85 68 92 69
rect 38 32 42 68
rect 28 28 42 32
rect 48 41 52 63
rect 48 39 49 41
rect 51 39 52 41
rect 28 22 32 28
rect 48 27 52 39
rect 58 41 62 63
rect 76 51 80 68
rect 88 62 92 68
rect 85 61 92 62
rect 85 59 87 61
rect 89 59 92 61
rect 85 58 92 59
rect 76 49 77 51
rect 79 49 80 51
rect 76 47 80 49
rect 58 39 59 41
rect 61 39 62 41
rect 58 27 62 39
rect 74 31 78 33
rect 88 32 92 58
rect 74 29 75 31
rect 77 29 78 31
rect 25 21 32 22
rect 25 19 27 21
rect 29 19 32 21
rect 25 18 32 19
rect 37 21 67 22
rect 37 19 39 21
rect 41 19 63 21
rect 65 19 67 21
rect 37 18 67 19
rect 74 21 78 29
rect 85 31 92 32
rect 85 29 87 31
rect 89 29 92 31
rect 85 28 92 29
rect 88 22 92 28
rect 74 19 75 21
rect 77 19 78 21
rect 74 12 78 19
rect 85 21 92 22
rect 85 19 87 21
rect 89 19 92 21
rect 85 18 92 19
rect 88 17 92 18
rect -2 11 102 12
rect -2 9 5 11
rect 7 9 51 11
rect 53 9 102 11
rect -2 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 102 9
rect -2 5 85 7
rect 87 5 93 7
rect 95 5 102 7
rect -2 0 102 5
<< ptie >>
rect 21 9 43 11
rect 21 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 43 9
rect 83 7 97 9
rect 21 5 43 7
rect 83 5 85 7
rect 87 5 93 7
rect 95 5 97 7
rect 83 3 97 5
<< nmos >>
rect 11 16 13 34
rect 21 17 23 34
rect 33 22 35 34
rect 45 22 47 34
rect 57 22 59 34
rect 81 15 83 35
<< pmos >>
rect 11 55 13 84
rect 23 56 25 85
rect 35 56 37 94
rect 47 55 49 94
rect 57 55 59 94
rect 81 56 83 94
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 77 49 79 51
rect 49 39 51 41
rect 59 39 61 41
<< ndifct1 >>
rect 27 19 29 21
rect 39 19 41 21
rect 63 19 65 21
rect 75 29 77 31
rect 75 19 77 21
rect 87 29 89 31
rect 87 19 89 21
rect 5 9 7 11
rect 51 9 53 11
<< ptiect1 >>
rect 23 7 25 9
rect 31 7 33 9
rect 39 7 41 9
rect 85 5 87 7
rect 93 5 95 7
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 29 79 31 81
rect 41 69 43 71
rect 63 79 65 81
rect 75 89 77 91
rect 75 79 77 81
rect 87 79 89 81
rect 87 69 89 71
rect 87 59 89 61
<< labels >>
rlabel alu1 10 45 10 45 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 30 55 30 55 6 i4
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 60 45 60 45 6 i3
rlabel alu1 50 94 50 94 6 vdd
rlabel alu1 90 50 90 50 6 q
<< end >>
