magic
tech scmos
timestamp 1199202744
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 59 11 65
rect 19 59 21 65
rect 31 57 33 61
rect 41 57 43 61
rect 9 35 11 40
rect 19 37 21 40
rect 31 37 33 40
rect 19 35 33 37
rect 41 35 43 40
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 27 35
rect 29 33 31 35
rect 19 31 31 33
rect 41 33 47 35
rect 41 31 43 33
rect 45 31 47 33
rect 12 26 14 29
rect 19 26 21 31
rect 29 26 31 31
rect 36 29 47 31
rect 36 26 38 29
rect 12 4 14 9
rect 19 4 21 9
rect 29 8 31 13
rect 36 8 38 13
<< ndif >>
rect 3 9 12 26
rect 14 9 19 26
rect 21 17 29 26
rect 21 15 24 17
rect 26 15 29 17
rect 21 13 29 15
rect 31 13 36 26
rect 38 17 46 26
rect 38 15 41 17
rect 43 15 46 17
rect 38 13 46 15
rect 21 9 26 13
rect 3 7 10 9
rect 3 5 6 7
rect 8 5 10 7
rect 3 3 10 5
<< pdif >>
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 40 9 48
rect 11 51 19 59
rect 11 49 14 51
rect 16 49 19 51
rect 11 44 19 49
rect 11 42 14 44
rect 16 42 19 44
rect 11 40 19 42
rect 21 57 29 59
rect 21 55 25 57
rect 27 55 31 57
rect 21 40 31 55
rect 33 55 41 57
rect 33 53 36 55
rect 38 53 41 55
rect 33 48 41 53
rect 33 46 36 48
rect 38 46 41 48
rect 33 40 41 46
rect 43 55 50 57
rect 43 53 46 55
rect 48 53 50 55
rect 43 48 50 53
rect 43 46 46 48
rect 48 46 50 48
rect 43 40 50 46
<< alu1 >>
rect -2 67 58 72
rect -2 65 35 67
rect 37 65 45 67
rect 47 65 58 67
rect -2 64 58 65
rect 34 55 40 59
rect 13 51 17 54
rect 13 49 14 51
rect 16 50 17 51
rect 34 53 36 55
rect 38 53 40 55
rect 34 50 40 53
rect 16 49 40 50
rect 13 48 40 49
rect 13 46 36 48
rect 38 46 40 48
rect 13 44 17 46
rect 13 43 14 44
rect 2 42 14 43
rect 16 42 17 44
rect 2 39 17 42
rect 2 18 6 39
rect 25 38 39 42
rect 25 35 31 38
rect 10 33 18 35
rect 10 31 11 33
rect 13 31 18 33
rect 10 29 18 31
rect 25 33 27 35
rect 29 33 31 35
rect 25 30 31 33
rect 41 33 47 34
rect 41 31 43 33
rect 45 31 47 33
rect 14 26 18 29
rect 41 26 47 31
rect 14 22 47 26
rect 2 17 31 18
rect 2 15 24 17
rect 26 15 31 17
rect 2 14 31 15
rect -2 7 58 8
rect -2 5 6 7
rect 8 5 46 7
rect 48 5 58 7
rect -2 0 58 5
<< ptie >>
rect 44 7 50 9
rect 44 5 46 7
rect 48 5 50 7
rect 44 3 50 5
<< ntie >>
rect 33 67 49 69
rect 33 65 35 67
rect 37 65 45 67
rect 47 65 49 67
rect 33 63 49 65
<< nmos >>
rect 12 9 14 26
rect 19 9 21 26
rect 29 13 31 26
rect 36 13 38 26
<< pmos >>
rect 9 40 11 59
rect 19 40 21 59
rect 31 40 33 57
rect 41 40 43 57
<< polyct1 >>
rect 11 31 13 33
rect 27 33 29 35
rect 43 31 45 33
<< ndifct0 >>
rect 41 15 43 17
<< ndifct1 >>
rect 24 15 26 17
rect 6 5 8 7
<< ntiect1 >>
rect 35 65 37 67
rect 45 65 47 67
<< ptiect1 >>
rect 46 5 48 7
<< pdifct0 >>
rect 4 55 6 57
rect 4 48 6 50
rect 25 55 27 57
rect 46 53 48 55
rect 46 46 48 48
<< pdifct1 >>
rect 14 49 16 51
rect 14 42 16 44
rect 36 53 38 55
rect 36 46 38 48
<< alu0 >>
rect 2 57 8 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 50 8 55
rect 23 57 29 64
rect 23 55 25 57
rect 27 55 29 57
rect 23 54 29 55
rect 2 48 4 50
rect 6 48 8 50
rect 2 47 8 48
rect 34 45 40 46
rect 44 55 50 64
rect 44 53 46 55
rect 48 53 50 55
rect 44 48 50 53
rect 44 46 46 48
rect 48 46 50 48
rect 44 45 50 46
rect 39 17 45 18
rect 39 15 41 17
rect 43 15 45 17
rect 39 8 45 15
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 20 24 20 24 6 a
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 16 28 16 6 z
rlabel alu1 28 24 28 24 6 a
rlabel alu1 36 24 36 24 6 a
rlabel alu1 36 40 36 40 6 b
rlabel alu1 28 36 28 36 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 28 44 28 6 a
<< end >>
