magic
tech scmos
timestamp 1199201652
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 65 31 70
rect 39 62 41 66
rect 9 42 11 45
rect 19 42 21 45
rect 9 40 21 42
rect 9 38 17 40
rect 19 38 21 40
rect 29 39 31 45
rect 9 36 21 38
rect 25 37 31 39
rect 9 30 11 36
rect 25 35 27 37
rect 29 35 31 37
rect 39 39 41 42
rect 39 37 47 39
rect 39 35 43 37
rect 45 35 47 37
rect 25 33 31 35
rect 35 33 47 35
rect 28 30 30 33
rect 35 30 37 33
rect 9 6 11 10
rect 28 8 30 13
rect 35 8 37 13
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 21 28 30
rect 11 19 15 21
rect 17 19 28 21
rect 11 14 28 19
rect 11 12 15 14
rect 17 13 28 14
rect 30 13 35 30
rect 37 23 42 30
rect 37 21 44 23
rect 37 19 40 21
rect 42 19 44 21
rect 37 17 44 19
rect 37 13 42 17
rect 17 12 26 13
rect 11 10 26 12
<< pdif >>
rect 2 63 9 65
rect 2 61 4 63
rect 6 61 9 63
rect 2 45 9 61
rect 11 61 19 65
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 45 19 52
rect 21 63 29 65
rect 21 61 24 63
rect 26 61 29 63
rect 21 45 29 61
rect 31 62 36 65
rect 31 60 39 62
rect 31 58 34 60
rect 36 58 39 60
rect 31 53 39 58
rect 31 51 34 53
rect 36 51 39 53
rect 31 45 39 51
rect 34 42 39 45
rect 41 60 48 62
rect 41 58 44 60
rect 46 58 48 60
rect 41 53 48 58
rect 41 51 44 53
rect 46 51 48 53
rect 41 42 48 51
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 55 17 59
rect 2 54 17 55
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 30 6 50
rect 33 42 47 46
rect 25 37 37 38
rect 25 35 27 37
rect 29 35 37 37
rect 25 34 37 35
rect 41 37 47 42
rect 41 35 43 37
rect 45 35 47 37
rect 41 34 47 35
rect 33 30 37 34
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 33 26 47 30
rect 2 21 7 26
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 10 11 30
rect 28 13 30 30
rect 35 13 37 30
<< pmos >>
rect 9 45 11 65
rect 19 45 21 65
rect 29 45 31 65
rect 39 42 41 62
<< polyct0 >>
rect 17 38 19 40
<< polyct1 >>
rect 27 35 29 37
rect 43 35 45 37
<< ndifct0 >>
rect 15 19 17 21
rect 15 12 17 14
rect 40 19 42 21
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 61 6 63
rect 24 61 26 63
rect 34 58 36 60
rect 34 51 36 53
rect 44 58 46 60
rect 44 51 46 53
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 3 63 7 68
rect 23 63 27 68
rect 3 61 4 63
rect 6 61 7 63
rect 3 59 7 61
rect 23 61 24 63
rect 26 61 27 63
rect 23 59 27 61
rect 33 60 38 62
rect 33 58 34 60
rect 36 58 38 60
rect 33 54 38 58
rect 23 53 38 54
rect 23 51 34 53
rect 36 51 38 53
rect 23 50 38 51
rect 42 60 48 68
rect 42 58 44 60
rect 46 58 48 60
rect 42 53 48 58
rect 42 51 44 53
rect 46 51 48 53
rect 42 50 48 51
rect 23 46 27 50
rect 16 42 27 46
rect 16 40 20 42
rect 16 38 17 40
rect 19 38 20 40
rect 16 30 20 38
rect 16 26 28 30
rect 24 22 28 26
rect 13 21 19 22
rect 13 19 15 21
rect 17 19 19 21
rect 13 14 19 19
rect 24 21 44 22
rect 24 19 40 21
rect 42 19 44 21
rect 24 18 44 19
rect 13 12 15 14
rect 17 12 19 14
<< labels >>
rlabel alu0 18 36 18 36 6 zn
rlabel alu0 30 52 30 52 6 zn
rlabel alu0 35 56 35 56 6 zn
rlabel alu0 34 20 34 20 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel polyct1 28 36 28 36 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 40 44 40 6 b
<< end >>
