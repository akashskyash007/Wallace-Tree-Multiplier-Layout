magic
tech scmos
timestamp 1199544097
<< ab >>
rect 0 0 280 100
<< nwell >>
rect -5 48 285 105
<< pwell >>
rect -5 -5 285 48
<< poly >>
rect 27 94 29 98
rect 39 94 41 98
rect 51 94 53 98
rect 59 94 61 98
rect 71 94 73 98
rect 83 94 85 98
rect 91 94 93 98
rect 15 70 17 74
rect 15 53 17 56
rect 7 51 17 53
rect 7 49 9 51
rect 11 49 17 51
rect 7 47 17 49
rect 15 37 17 47
rect 27 53 29 75
rect 39 73 41 76
rect 33 71 41 73
rect 33 69 35 71
rect 37 69 41 71
rect 33 67 41 69
rect 195 94 197 98
rect 207 94 209 98
rect 219 94 221 98
rect 231 94 233 98
rect 243 94 245 98
rect 255 94 257 98
rect 267 94 269 98
rect 121 85 123 89
rect 147 85 149 89
rect 159 85 161 89
rect 171 85 173 89
rect 183 85 185 89
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 15 25 17 29
rect 27 23 29 47
rect 39 41 41 67
rect 51 63 53 75
rect 47 61 53 63
rect 47 59 49 61
rect 51 59 53 61
rect 47 57 53 59
rect 47 51 53 53
rect 59 51 61 75
rect 71 73 73 76
rect 83 73 85 76
rect 47 49 49 51
rect 51 49 61 51
rect 47 47 53 49
rect 39 39 53 41
rect 33 31 41 33
rect 33 29 35 31
rect 37 29 41 31
rect 33 27 41 29
rect 39 23 41 27
rect 51 23 53 39
rect 59 23 61 49
rect 69 71 73 73
rect 79 71 85 73
rect 69 33 71 71
rect 79 53 81 71
rect 91 63 93 76
rect 103 69 105 73
rect 85 61 93 63
rect 85 59 87 61
rect 89 59 93 61
rect 85 57 93 59
rect 75 51 81 53
rect 103 51 105 55
rect 121 53 123 65
rect 147 63 149 66
rect 159 63 161 66
rect 171 63 173 66
rect 195 73 197 76
rect 195 71 203 73
rect 195 69 199 71
rect 201 69 203 71
rect 195 67 203 69
rect 141 61 149 63
rect 157 61 163 63
rect 75 49 77 51
rect 79 49 105 51
rect 75 47 81 49
rect 79 39 81 47
rect 65 31 71 33
rect 65 29 67 31
rect 69 29 71 31
rect 65 27 71 29
rect 75 37 81 39
rect 85 41 93 43
rect 85 39 87 41
rect 89 39 93 41
rect 85 37 93 39
rect 103 37 105 49
rect 117 51 123 53
rect 117 49 119 51
rect 121 49 123 51
rect 117 47 123 49
rect 129 51 135 53
rect 141 51 143 61
rect 157 59 159 61
rect 161 59 163 61
rect 157 57 163 59
rect 169 61 175 63
rect 169 59 171 61
rect 173 59 175 61
rect 169 57 175 59
rect 167 51 173 53
rect 183 51 185 65
rect 207 63 209 75
rect 201 61 209 63
rect 201 59 203 61
rect 205 59 209 61
rect 201 57 209 59
rect 219 51 221 75
rect 231 73 233 76
rect 225 71 233 73
rect 225 69 227 71
rect 229 69 233 71
rect 225 67 233 69
rect 243 53 245 75
rect 243 51 251 53
rect 129 49 131 51
rect 133 49 169 51
rect 171 49 233 51
rect 129 47 135 49
rect 75 23 77 37
rect 81 31 87 33
rect 81 29 83 31
rect 85 29 87 31
rect 81 27 87 29
rect 71 21 77 23
rect 71 18 73 21
rect 83 19 85 27
rect 91 19 93 37
rect 103 25 105 29
rect 121 25 123 47
rect 141 29 143 49
rect 167 47 173 49
rect 147 41 153 43
rect 177 41 185 43
rect 219 41 227 43
rect 147 39 149 41
rect 151 39 179 41
rect 181 39 223 41
rect 225 39 227 41
rect 147 37 153 39
rect 177 37 185 39
rect 157 31 163 33
rect 157 29 159 31
rect 161 29 163 31
rect 141 27 149 29
rect 157 27 163 29
rect 169 31 175 33
rect 169 29 171 31
rect 173 29 175 31
rect 169 27 175 29
rect 27 7 29 11
rect 39 7 41 11
rect 51 7 53 11
rect 59 7 61 11
rect 147 24 149 27
rect 159 24 161 27
rect 171 24 173 27
rect 183 25 185 37
rect 219 37 227 39
rect 201 31 209 33
rect 201 29 203 31
rect 205 29 209 31
rect 201 27 209 29
rect 121 11 123 15
rect 147 11 149 15
rect 159 11 161 15
rect 171 11 173 15
rect 183 11 185 15
rect 195 21 203 23
rect 195 19 199 21
rect 201 19 203 21
rect 195 17 203 19
rect 195 14 197 17
rect 207 15 209 27
rect 219 25 221 37
rect 231 25 233 49
rect 243 49 247 51
rect 249 49 251 51
rect 243 47 251 49
rect 255 43 257 55
rect 267 43 269 55
rect 245 41 269 43
rect 245 39 247 41
rect 249 39 269 41
rect 245 37 269 39
rect 243 31 251 33
rect 243 29 247 31
rect 249 29 251 31
rect 243 27 251 29
rect 243 24 245 27
rect 255 25 257 37
rect 267 25 269 37
rect 71 2 73 6
rect 83 3 85 7
rect 91 3 93 7
rect 219 11 221 15
rect 231 11 233 15
rect 243 11 245 15
rect 195 2 197 6
rect 207 2 209 6
rect 255 2 257 6
rect 267 2 269 6
<< ndif >>
rect 7 29 15 37
rect 17 33 25 37
rect 17 31 21 33
rect 23 31 25 33
rect 17 29 25 31
rect 7 21 13 29
rect 43 31 49 33
rect 43 29 45 31
rect 47 29 49 31
rect 43 23 49 29
rect 7 19 9 21
rect 11 19 13 21
rect 7 17 13 19
rect 19 21 27 23
rect 19 19 21 21
rect 23 19 27 21
rect 19 11 27 19
rect 29 11 39 23
rect 41 11 51 23
rect 53 11 59 23
rect 61 21 69 23
rect 61 19 65 21
rect 67 19 69 21
rect 61 18 69 19
rect 95 35 103 37
rect 95 33 97 35
rect 99 33 103 35
rect 95 29 103 33
rect 105 29 117 37
rect 107 25 117 29
rect 95 21 101 23
rect 95 19 97 21
rect 99 19 101 21
rect 78 18 83 19
rect 61 11 71 18
rect 63 6 71 11
rect 73 11 83 18
rect 73 9 77 11
rect 79 9 83 11
rect 73 7 83 9
rect 85 7 91 19
rect 93 9 101 19
rect 107 15 121 25
rect 123 21 133 25
rect 178 24 183 25
rect 123 19 129 21
rect 131 19 133 21
rect 123 15 133 19
rect 139 21 147 24
rect 139 19 141 21
rect 143 19 147 21
rect 139 15 147 19
rect 149 15 159 24
rect 161 15 171 24
rect 173 21 183 24
rect 173 19 177 21
rect 179 19 183 21
rect 173 15 183 19
rect 185 15 193 25
rect 107 11 117 15
rect 151 11 157 15
rect 187 14 193 15
rect 211 21 219 25
rect 211 19 213 21
rect 215 19 219 21
rect 211 15 219 19
rect 221 21 231 25
rect 221 19 225 21
rect 227 19 231 21
rect 221 15 231 19
rect 233 24 238 25
rect 250 24 255 25
rect 233 15 243 24
rect 245 21 255 24
rect 245 19 249 21
rect 251 19 255 21
rect 245 15 255 19
rect 202 14 207 15
rect 107 9 109 11
rect 111 9 117 11
rect 151 9 153 11
rect 155 9 157 11
rect 93 7 98 9
rect 107 7 117 9
rect 151 7 157 9
rect 73 6 80 7
rect 187 6 195 14
rect 197 11 207 14
rect 197 9 201 11
rect 203 9 207 11
rect 197 6 207 9
rect 209 6 217 15
rect 247 11 255 15
rect 247 9 249 11
rect 251 9 255 11
rect 247 6 255 9
rect 257 21 267 25
rect 257 19 261 21
rect 263 19 267 21
rect 257 6 267 19
rect 269 21 277 25
rect 269 19 273 21
rect 275 19 277 21
rect 269 11 277 19
rect 269 9 273 11
rect 275 9 277 11
rect 269 6 277 9
<< pdif >>
rect 7 81 13 83
rect 7 79 9 81
rect 11 79 13 81
rect 7 70 13 79
rect 19 81 27 94
rect 19 79 21 81
rect 23 79 27 81
rect 19 75 27 79
rect 29 76 39 94
rect 41 76 51 94
rect 29 75 34 76
rect 7 56 15 70
rect 17 61 25 70
rect 17 59 21 61
rect 23 59 25 61
rect 17 56 25 59
rect 43 75 51 76
rect 53 75 59 94
rect 61 81 71 94
rect 61 79 65 81
rect 67 79 71 81
rect 61 76 71 79
rect 73 91 83 94
rect 73 89 77 91
rect 79 89 83 91
rect 73 76 83 89
rect 85 76 91 94
rect 93 81 101 94
rect 93 79 97 81
rect 99 79 101 81
rect 93 76 101 79
rect 107 91 117 93
rect 151 93 157 95
rect 151 91 153 93
rect 155 91 157 93
rect 107 89 109 91
rect 111 89 117 91
rect 107 85 117 89
rect 151 85 157 91
rect 187 85 195 94
rect 61 75 66 76
rect 43 71 49 75
rect 43 69 45 71
rect 47 69 49 71
rect 43 67 49 69
rect 107 69 121 85
rect 95 61 103 69
rect 95 59 97 61
rect 99 59 103 61
rect 95 55 103 59
rect 105 65 121 69
rect 123 71 133 85
rect 123 69 129 71
rect 131 69 133 71
rect 123 65 133 69
rect 139 71 147 85
rect 139 69 141 71
rect 143 69 147 71
rect 139 66 147 69
rect 149 66 159 85
rect 161 66 171 85
rect 173 71 183 85
rect 173 69 177 71
rect 179 69 183 71
rect 173 66 183 69
rect 105 55 117 65
rect 178 65 183 66
rect 185 76 195 85
rect 197 91 207 94
rect 197 89 201 91
rect 203 89 207 91
rect 197 76 207 89
rect 185 65 193 76
rect 202 75 207 76
rect 209 81 219 94
rect 209 79 213 81
rect 215 79 219 81
rect 209 75 219 79
rect 221 81 231 94
rect 221 79 225 81
rect 227 79 231 81
rect 221 76 231 79
rect 233 76 243 94
rect 221 75 226 76
rect 238 75 243 76
rect 245 91 255 94
rect 245 89 249 91
rect 251 89 255 91
rect 245 81 255 89
rect 245 79 249 81
rect 251 79 255 81
rect 245 75 255 79
rect 247 71 255 75
rect 247 69 249 71
rect 251 69 255 71
rect 247 61 255 69
rect 247 59 249 61
rect 251 59 255 61
rect 247 55 255 59
rect 257 81 267 94
rect 257 79 261 81
rect 263 79 267 81
rect 257 71 267 79
rect 257 69 261 71
rect 263 69 267 71
rect 257 61 267 69
rect 257 59 261 61
rect 263 59 267 61
rect 257 55 267 59
rect 269 91 277 94
rect 269 89 273 91
rect 275 89 277 91
rect 269 81 277 89
rect 269 79 273 81
rect 275 79 277 81
rect 269 71 277 79
rect 269 69 273 71
rect 275 69 277 71
rect 269 61 277 69
rect 269 59 273 61
rect 275 59 277 61
rect 269 55 277 59
<< alu1 >>
rect -2 95 282 100
rect -2 93 127 95
rect 129 93 141 95
rect 143 93 165 95
rect 167 93 177 95
rect 179 93 282 95
rect -2 91 153 93
rect 155 91 282 93
rect -2 89 77 91
rect 79 89 109 91
rect 111 89 201 91
rect 203 89 249 91
rect 251 89 273 91
rect 275 89 282 91
rect -2 88 282 89
rect 8 81 12 88
rect 96 82 100 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 77 12 79
rect 19 81 69 82
rect 19 79 21 81
rect 23 79 65 81
rect 67 79 69 81
rect 19 78 69 79
rect 96 81 162 82
rect 96 79 97 81
rect 99 79 162 81
rect 96 78 162 79
rect 8 72 12 73
rect 96 72 100 78
rect 8 71 39 72
rect 8 69 35 71
rect 37 69 39 71
rect 8 68 39 69
rect 43 71 112 72
rect 43 69 45 71
rect 47 69 112 71
rect 43 68 112 69
rect 8 51 12 68
rect 8 49 9 51
rect 11 49 12 51
rect 8 27 12 49
rect 18 61 53 62
rect 18 59 21 61
rect 23 59 49 61
rect 51 59 53 61
rect 18 58 53 59
rect 18 34 22 58
rect 28 51 32 53
rect 28 49 29 51
rect 31 49 32 51
rect 28 41 32 49
rect 39 51 53 52
rect 39 49 49 51
rect 51 49 53 51
rect 39 48 53 49
rect 58 42 62 68
rect 54 38 62 42
rect 68 52 72 63
rect 86 62 90 63
rect 77 61 90 62
rect 77 59 87 61
rect 89 59 90 61
rect 77 58 90 59
rect 95 61 102 62
rect 95 59 97 61
rect 99 59 102 61
rect 95 58 102 59
rect 86 52 90 58
rect 68 51 81 52
rect 68 49 77 51
rect 79 49 81 51
rect 68 48 81 49
rect 86 48 93 52
rect 18 33 25 34
rect 18 31 21 33
rect 23 32 25 33
rect 54 32 58 38
rect 68 37 72 48
rect 86 42 90 48
rect 77 41 90 42
rect 77 39 87 41
rect 89 39 90 41
rect 77 38 90 39
rect 86 37 90 38
rect 98 37 102 58
rect 96 35 102 37
rect 96 33 97 35
rect 99 33 102 35
rect 96 32 102 33
rect 23 31 39 32
rect 18 30 35 31
rect 20 29 35 30
rect 37 29 39 31
rect 20 28 39 29
rect 43 31 58 32
rect 43 29 45 31
rect 47 29 58 31
rect 43 28 58 29
rect 65 31 100 32
rect 65 29 67 31
rect 69 29 83 31
rect 85 29 100 31
rect 65 28 100 29
rect 8 21 12 23
rect 108 22 112 68
rect 8 19 9 21
rect 11 19 12 21
rect 8 12 12 19
rect 19 21 69 22
rect 19 19 21 21
rect 23 19 65 21
rect 67 19 69 21
rect 19 18 69 19
rect 95 21 112 22
rect 95 19 97 21
rect 99 19 112 21
rect 95 18 112 19
rect 118 51 122 73
rect 118 49 119 51
rect 121 49 122 51
rect 118 17 122 49
rect 128 71 132 73
rect 128 69 129 71
rect 131 69 132 71
rect 128 52 132 69
rect 139 71 145 72
rect 139 69 141 71
rect 143 69 152 71
rect 139 68 152 69
rect 140 67 152 68
rect 128 51 135 52
rect 128 49 131 51
rect 133 49 135 51
rect 128 48 135 49
rect 128 21 132 48
rect 148 41 152 67
rect 148 39 149 41
rect 151 39 152 41
rect 148 23 152 39
rect 158 61 162 78
rect 212 81 216 83
rect 212 79 213 81
rect 215 79 216 81
rect 212 72 216 79
rect 223 81 240 82
rect 223 79 225 81
rect 227 79 240 81
rect 223 78 240 79
rect 175 71 192 72
rect 175 69 177 71
rect 179 69 192 71
rect 175 68 192 69
rect 197 71 216 72
rect 197 69 199 71
rect 201 69 216 71
rect 197 68 216 69
rect 188 62 192 68
rect 158 59 159 61
rect 161 59 162 61
rect 158 31 162 59
rect 169 61 182 62
rect 169 59 171 61
rect 173 59 182 61
rect 169 58 182 59
rect 158 29 159 31
rect 161 29 162 31
rect 158 27 162 29
rect 168 51 172 53
rect 168 49 169 51
rect 171 49 172 51
rect 168 32 172 49
rect 178 41 182 58
rect 178 39 179 41
rect 181 39 182 41
rect 178 37 182 39
rect 188 61 207 62
rect 188 59 203 61
rect 205 59 207 61
rect 188 58 207 59
rect 188 32 192 58
rect 168 31 175 32
rect 168 29 171 31
rect 173 29 175 31
rect 168 28 175 29
rect 188 31 207 32
rect 188 29 203 31
rect 205 29 207 31
rect 188 28 207 29
rect 140 22 152 23
rect 188 22 192 28
rect 212 22 216 68
rect 224 71 231 72
rect 224 69 227 71
rect 229 69 231 71
rect 224 68 231 69
rect 224 42 228 68
rect 221 41 228 42
rect 221 39 223 41
rect 225 39 228 41
rect 221 38 228 39
rect 236 42 240 78
rect 248 81 252 88
rect 248 79 249 81
rect 251 79 252 81
rect 248 71 252 79
rect 248 69 249 71
rect 251 69 252 71
rect 248 61 252 69
rect 248 59 249 61
rect 251 59 252 61
rect 248 57 252 59
rect 258 82 262 83
rect 258 81 265 82
rect 258 79 261 81
rect 263 79 265 81
rect 258 78 265 79
rect 272 81 276 88
rect 272 79 273 81
rect 275 79 276 81
rect 258 72 262 78
rect 258 71 265 72
rect 258 69 261 71
rect 263 69 265 71
rect 258 68 265 69
rect 272 71 276 79
rect 272 69 273 71
rect 275 69 276 71
rect 258 62 262 68
rect 258 61 265 62
rect 258 59 261 61
rect 263 59 265 61
rect 258 58 265 59
rect 272 61 276 69
rect 272 59 273 61
rect 275 59 276 61
rect 258 52 262 58
rect 272 57 276 59
rect 245 51 263 52
rect 245 49 247 51
rect 249 49 263 51
rect 245 48 263 49
rect 236 41 251 42
rect 236 39 247 41
rect 249 39 251 41
rect 236 38 251 39
rect 236 22 240 38
rect 258 32 262 48
rect 245 31 263 32
rect 245 29 247 31
rect 249 29 263 31
rect 245 28 263 29
rect 128 19 129 21
rect 131 19 132 21
rect 128 17 132 19
rect 139 21 152 22
rect 139 19 141 21
rect 143 19 152 21
rect 175 21 192 22
rect 175 19 177 21
rect 179 19 192 21
rect 139 18 145 19
rect 175 18 192 19
rect 197 21 216 22
rect 197 19 199 21
rect 201 19 213 21
rect 215 19 216 21
rect 197 18 216 19
rect 223 21 240 22
rect 223 19 225 21
rect 227 19 240 21
rect 223 18 240 19
rect 248 21 252 23
rect 248 19 249 21
rect 251 19 252 21
rect 212 17 216 18
rect 248 12 252 19
rect 258 22 262 28
rect 258 21 265 22
rect 258 19 261 21
rect 263 19 265 21
rect 258 18 265 19
rect 272 21 276 23
rect 272 19 273 21
rect 275 19 276 21
rect 258 17 262 18
rect 272 12 276 19
rect -2 11 282 12
rect -2 9 77 11
rect 79 9 109 11
rect 111 9 153 11
rect 155 9 201 11
rect 203 9 249 11
rect 251 9 273 11
rect 275 9 282 11
rect -2 7 282 9
rect -2 5 127 7
rect 129 5 141 7
rect 143 5 165 7
rect 167 5 177 7
rect 179 5 225 7
rect 227 5 237 7
rect 239 5 282 7
rect -2 0 282 5
<< ptie >>
rect 125 7 145 9
rect 163 7 181 9
rect 125 5 127 7
rect 129 5 141 7
rect 143 5 145 7
rect 125 3 145 5
rect 163 5 165 7
rect 167 5 177 7
rect 179 5 181 7
rect 223 7 241 9
rect 163 3 181 5
rect 223 5 225 7
rect 227 5 237 7
rect 239 5 241 7
rect 223 3 241 5
<< ntie >>
rect 125 95 145 97
rect 163 95 181 97
rect 125 93 127 95
rect 129 93 141 95
rect 143 93 145 95
rect 125 91 145 93
rect 163 93 165 95
rect 167 93 177 95
rect 179 93 181 95
rect 163 91 181 93
<< nmos >>
rect 15 29 17 37
rect 27 11 29 23
rect 39 11 41 23
rect 51 11 53 23
rect 59 11 61 23
rect 103 29 105 37
rect 71 6 73 18
rect 83 7 85 19
rect 91 7 93 19
rect 121 15 123 25
rect 147 15 149 24
rect 159 15 161 24
rect 171 15 173 24
rect 183 15 185 25
rect 219 15 221 25
rect 231 15 233 25
rect 243 15 245 24
rect 195 6 197 14
rect 207 6 209 15
rect 255 6 257 25
rect 267 6 269 25
<< pmos >>
rect 27 75 29 94
rect 39 76 41 94
rect 15 56 17 70
rect 51 75 53 94
rect 59 75 61 94
rect 71 76 73 94
rect 83 76 85 94
rect 91 76 93 94
rect 103 55 105 69
rect 121 65 123 85
rect 147 66 149 85
rect 159 66 161 85
rect 171 66 173 85
rect 183 65 185 85
rect 195 76 197 94
rect 207 75 209 94
rect 219 75 221 94
rect 231 76 233 94
rect 243 75 245 94
rect 255 55 257 94
rect 267 55 269 94
<< polyct1 >>
rect 9 49 11 51
rect 35 69 37 71
rect 29 49 31 51
rect 49 59 51 61
rect 49 49 51 51
rect 35 29 37 31
rect 87 59 89 61
rect 199 69 201 71
rect 77 49 79 51
rect 67 29 69 31
rect 87 39 89 41
rect 119 49 121 51
rect 159 59 161 61
rect 171 59 173 61
rect 203 59 205 61
rect 227 69 229 71
rect 131 49 133 51
rect 169 49 171 51
rect 83 29 85 31
rect 149 39 151 41
rect 179 39 181 41
rect 223 39 225 41
rect 159 29 161 31
rect 171 29 173 31
rect 203 29 205 31
rect 199 19 201 21
rect 247 49 249 51
rect 247 39 249 41
rect 247 29 249 31
<< ndifct1 >>
rect 21 31 23 33
rect 45 29 47 31
rect 9 19 11 21
rect 21 19 23 21
rect 65 19 67 21
rect 97 33 99 35
rect 97 19 99 21
rect 77 9 79 11
rect 129 19 131 21
rect 141 19 143 21
rect 177 19 179 21
rect 213 19 215 21
rect 225 19 227 21
rect 249 19 251 21
rect 109 9 111 11
rect 153 9 155 11
rect 201 9 203 11
rect 249 9 251 11
rect 261 19 263 21
rect 273 19 275 21
rect 273 9 275 11
<< ntiect1 >>
rect 127 93 129 95
rect 141 93 143 95
rect 165 93 167 95
rect 177 93 179 95
<< ptiect1 >>
rect 127 5 129 7
rect 141 5 143 7
rect 165 5 167 7
rect 177 5 179 7
rect 225 5 227 7
rect 237 5 239 7
<< pdifct1 >>
rect 9 79 11 81
rect 21 79 23 81
rect 21 59 23 61
rect 65 79 67 81
rect 77 89 79 91
rect 97 79 99 81
rect 153 91 155 93
rect 109 89 111 91
rect 45 69 47 71
rect 97 59 99 61
rect 129 69 131 71
rect 141 69 143 71
rect 177 69 179 71
rect 201 89 203 91
rect 213 79 215 81
rect 225 79 227 81
rect 249 89 251 91
rect 249 79 251 81
rect 249 69 251 71
rect 249 59 251 61
rect 261 79 263 81
rect 261 69 263 71
rect 261 59 263 61
rect 273 89 275 91
rect 273 79 275 81
rect 273 69 275 71
rect 273 59 275 61
<< labels >>
rlabel polyct1 50 50 50 50 6 i1
rlabel polyct1 10 50 10 50 6 cmd1
rlabel polyct1 30 50 30 50 6 i2
rlabel alu1 80 40 80 40 6 i0
rlabel alu1 90 50 90 50 6 i0
rlabel alu1 70 50 70 50 6 cmd0
rlabel alu1 80 60 80 60 6 i0
rlabel alu1 140 6 140 6 6 vss
rlabel alu1 120 45 120 45 6 ck
rlabel alu1 140 94 140 94 6 vdd
rlabel alu1 250 30 250 30 6 q
rlabel alu1 260 50 260 50 6 q
rlabel alu1 250 50 250 50 6 q
<< end >>
