magic
tech scmos
timestamp 1199469704
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 15 94 17 98
rect 23 94 25 98
rect 35 94 37 98
rect 43 94 45 98
rect 57 80 59 85
rect 15 53 17 56
rect 8 51 17 53
rect 8 49 10 51
rect 12 50 17 51
rect 12 49 19 50
rect 8 47 19 49
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 11 31 13 37
rect 17 37 19 47
rect 23 43 25 56
rect 35 53 37 56
rect 29 51 37 53
rect 29 49 31 51
rect 33 49 37 51
rect 29 47 37 49
rect 23 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 43 41 45 56
rect 57 53 59 56
rect 51 51 59 53
rect 51 49 53 51
rect 55 49 59 51
rect 51 47 59 49
rect 43 39 52 41
rect 43 37 48 39
rect 50 37 52 39
rect 17 34 21 37
rect 19 31 21 34
rect 31 31 33 37
rect 39 35 52 37
rect 39 31 41 35
rect 57 31 59 47
rect 57 14 59 19
rect 11 9 13 14
rect 19 9 21 14
rect 31 9 33 14
rect 39 9 41 14
<< ndif >>
rect 3 14 11 31
rect 13 14 19 31
rect 21 21 31 31
rect 21 19 25 21
rect 27 19 31 21
rect 21 14 31 19
rect 33 14 39 31
rect 41 29 57 31
rect 41 27 49 29
rect 51 27 57 29
rect 41 21 57 27
rect 41 19 49 21
rect 51 19 57 21
rect 59 29 67 31
rect 59 27 63 29
rect 65 27 67 29
rect 59 25 67 27
rect 59 19 64 25
rect 41 14 55 19
rect 3 10 9 14
rect 3 8 5 10
rect 7 8 9 10
rect 3 6 9 8
<< pdif >>
rect 6 91 15 94
rect 6 89 9 91
rect 11 89 15 91
rect 6 81 15 89
rect 6 79 9 81
rect 11 79 15 81
rect 6 56 15 79
rect 17 56 23 94
rect 25 61 35 94
rect 25 59 29 61
rect 31 59 35 61
rect 25 56 35 59
rect 37 56 43 94
rect 45 91 55 94
rect 45 89 49 91
rect 51 89 55 91
rect 45 81 55 89
rect 45 79 49 81
rect 51 80 55 81
rect 51 79 57 80
rect 45 56 57 79
rect 59 70 64 80
rect 59 68 67 70
rect 59 66 63 68
rect 65 66 67 68
rect 59 60 67 66
rect 59 58 63 60
rect 65 58 67 60
rect 59 56 67 58
<< alu1 >>
rect -2 95 72 100
rect -2 93 63 95
rect 65 93 72 95
rect -2 91 72 93
rect -2 89 9 91
rect 11 89 49 91
rect 51 89 72 91
rect -2 88 72 89
rect 8 81 12 88
rect 8 79 9 81
rect 11 79 12 81
rect 8 77 12 79
rect 48 81 52 88
rect 48 79 49 81
rect 51 79 52 81
rect 48 77 52 79
rect 7 68 53 72
rect 7 51 13 68
rect 7 49 10 51
rect 12 49 13 51
rect 7 47 13 49
rect 18 53 22 63
rect 28 61 42 63
rect 28 59 29 61
rect 31 59 42 61
rect 28 57 42 59
rect 18 51 34 53
rect 18 49 31 51
rect 33 49 34 51
rect 18 47 34 49
rect 18 43 22 47
rect 7 41 22 43
rect 7 39 9 41
rect 11 39 22 41
rect 7 37 22 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 32 33 39
rect 7 28 33 32
rect 7 18 13 28
rect 38 22 42 57
rect 47 53 53 68
rect 62 68 66 70
rect 62 66 63 68
rect 65 66 66 68
rect 62 60 66 66
rect 62 58 63 60
rect 65 58 66 60
rect 47 51 57 53
rect 47 49 53 51
rect 55 49 57 51
rect 47 47 57 49
rect 62 40 66 58
rect 46 39 66 40
rect 46 37 48 39
rect 50 37 66 39
rect 46 36 66 37
rect 23 21 42 22
rect 23 19 25 21
rect 27 19 42 21
rect 23 17 42 19
rect 48 29 52 31
rect 48 27 49 29
rect 51 27 52 29
rect 48 21 52 27
rect 62 29 66 36
rect 62 27 63 29
rect 65 27 66 29
rect 62 25 66 27
rect 48 19 49 21
rect 51 19 52 21
rect 48 12 52 19
rect -2 10 72 12
rect -2 8 5 10
rect 7 8 72 10
rect -2 7 72 8
rect -2 5 63 7
rect 65 5 72 7
rect -2 0 72 5
<< ptie >>
rect 61 7 67 9
rect 61 5 63 7
rect 65 5 67 7
rect 61 3 67 5
<< ntie >>
rect 61 95 67 97
rect 61 93 63 95
rect 65 93 67 95
rect 61 91 67 93
<< nmos >>
rect 11 14 13 31
rect 19 14 21 31
rect 31 14 33 31
rect 39 14 41 31
rect 57 19 59 31
<< pmos >>
rect 15 56 17 94
rect 23 56 25 94
rect 35 56 37 94
rect 43 56 45 94
rect 57 56 59 80
<< polyct1 >>
rect 10 49 12 51
rect 9 39 11 41
rect 31 49 33 51
rect 29 39 31 41
rect 53 49 55 51
rect 48 37 50 39
<< ndifct1 >>
rect 25 19 27 21
rect 49 27 51 29
rect 49 19 51 21
rect 63 27 65 29
rect 5 8 7 10
<< ntiect1 >>
rect 63 93 65 95
<< ptiect1 >>
rect 63 5 65 7
<< pdifct1 >>
rect 9 89 11 91
rect 9 79 11 81
rect 29 59 31 61
rect 49 89 51 91
rect 49 79 51 81
rect 63 66 65 68
rect 63 58 65 60
<< labels >>
rlabel ndifct1 64 28 64 28 6 sn
rlabel polyct1 49 38 49 38 6 sn
rlabel pdifct1 64 59 64 59 6 sn
rlabel pdifct1 64 67 64 67 6 sn
rlabel alu1 10 25 10 25 6 a0
rlabel polyct1 10 40 10 40 6 a1
rlabel alu1 10 60 10 60 6 s
rlabel alu1 30 20 30 20 6 z
rlabel alu1 20 30 20 30 6 a0
rlabel alu1 30 35 30 35 6 a0
rlabel alu1 30 50 30 50 6 a1
rlabel alu1 20 50 20 50 6 a1
rlabel alu1 20 70 20 70 6 s
rlabel alu1 30 70 30 70 6 s
rlabel pdifct1 30 60 30 60 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 40 40 40 6 z
rlabel alu1 40 70 40 70 6 s
rlabel alu1 50 60 50 60 6 s
rlabel alu1 35 94 35 94 6 vdd
<< end >>
