magic
tech scmos
timestamp 1199543798
<< ab >>
rect 0 0 30 100
<< nwell >>
rect -2 48 32 104
<< pwell >>
rect -2 -4 32 48
<< poly >>
rect 13 75 15 78
rect 13 53 15 55
rect 7 51 15 53
rect 7 49 9 51
rect 11 49 15 51
rect 7 47 15 49
<< pdif >>
rect 3 71 13 75
rect 3 69 7 71
rect 9 69 13 71
rect 3 61 13 69
rect 3 59 7 61
rect 9 59 13 61
rect 3 55 13 59
rect 15 71 23 75
rect 15 69 19 71
rect 21 69 23 71
rect 15 61 23 69
rect 15 59 19 61
rect 21 59 23 61
rect 15 55 23 59
<< alu1 >>
rect -2 91 32 100
rect -2 89 7 91
rect 9 89 19 91
rect 21 89 32 91
rect -2 88 32 89
rect 6 71 10 88
rect 6 69 7 71
rect 9 69 10 71
rect 6 61 10 69
rect 6 59 7 61
rect 9 59 10 61
rect 6 58 10 59
rect 18 71 22 82
rect 18 69 19 71
rect 21 69 22 71
rect 18 61 22 69
rect 18 59 19 61
rect 21 59 22 61
rect 8 51 12 52
rect 8 49 9 51
rect 11 49 12 51
rect 8 31 12 49
rect 8 29 9 31
rect 11 29 12 31
rect 8 21 12 29
rect 8 19 9 21
rect 11 19 12 21
rect 8 12 12 19
rect 18 18 22 59
rect -2 11 32 12
rect -2 9 9 11
rect 11 9 19 11
rect 21 9 32 11
rect -2 0 32 9
<< ptie >>
rect 7 31 13 33
rect 7 29 9 31
rect 11 29 13 31
rect 7 21 13 29
rect 7 19 9 21
rect 11 19 13 21
rect 7 13 13 19
rect 7 11 23 13
rect 7 9 9 11
rect 11 9 19 11
rect 21 9 23 11
rect 7 7 23 9
<< ntie >>
rect 5 91 23 93
rect 5 89 7 91
rect 9 89 19 91
rect 21 89 23 91
rect 5 87 23 89
<< pmos >>
rect 13 55 15 75
<< polyct1 >>
rect 9 49 11 51
<< ntiect1 >>
rect 7 89 9 91
rect 19 89 21 91
<< ptiect1 >>
rect 9 29 11 31
rect 9 19 11 21
rect 9 9 11 11
rect 19 9 21 11
<< pdifct1 >>
rect 7 69 9 71
rect 7 59 9 61
rect 19 69 21 71
rect 19 59 21 61
<< labels >>
rlabel alu1 15 6 15 6 6 vss
rlabel alu1 20 50 20 50 6 q
rlabel alu1 15 94 15 94 6 vdd
<< end >>
