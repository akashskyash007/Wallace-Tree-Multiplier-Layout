magic
tech scmos
timestamp 1199980689
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -8 40 104 97
<< pwell >>
rect -8 -9 104 40
<< poly >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 69 84 78 86
rect 69 82 74 84
rect 76 82 78 84
rect 69 80 78 82
rect 82 84 91 86
rect 82 82 84 84
rect 86 82 91 84
rect 82 80 91 82
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 49 46
rect 51 44 62 46
rect 47 42 62 44
rect 66 46 75 48
rect 66 44 71 46
rect 73 44 75 46
rect 66 42 75 44
rect 79 42 94 48
rect 2 32 17 38
rect 21 32 30 38
rect 34 36 49 38
rect 34 34 36 36
rect 38 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 66 36 81 38
rect 66 34 71 36
rect 73 34 81 36
rect 66 32 81 34
rect 85 32 94 38
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 6 27 8
rect 18 4 23 6
rect 25 4 27 6
rect 18 2 27 4
rect 37 2 46 8
rect 50 2 59 8
rect 69 2 78 8
rect 82 6 91 8
rect 82 4 84 6
rect 86 4 91 6
rect 82 2 91 4
<< ndif >>
rect 2 11 9 29
rect 11 11 21 29
rect 23 11 30 29
rect 34 24 41 29
rect 34 22 36 24
rect 38 22 41 24
rect 34 17 41 22
rect 34 15 36 17
rect 38 15 41 17
rect 34 11 41 15
rect 43 16 53 29
rect 43 14 47 16
rect 49 14 53 16
rect 43 11 53 14
rect 55 25 62 29
rect 55 23 58 25
rect 60 23 62 25
rect 55 18 62 23
rect 55 16 58 18
rect 60 16 62 18
rect 55 11 62 16
rect 66 25 73 29
rect 66 23 68 25
rect 70 23 73 25
rect 66 18 73 23
rect 66 16 68 18
rect 70 16 73 18
rect 66 11 73 16
rect 75 16 85 29
rect 75 14 79 16
rect 81 14 85 16
rect 75 11 85 14
rect 87 11 94 29
<< pdif >>
rect 2 74 9 77
rect 2 72 4 74
rect 6 72 9 74
rect 2 67 9 72
rect 2 65 4 67
rect 6 65 9 67
rect 2 51 9 65
rect 11 65 21 77
rect 11 63 15 65
rect 17 63 21 65
rect 11 58 21 63
rect 11 56 15 58
rect 17 56 21 58
rect 11 51 21 56
rect 23 74 30 77
rect 23 72 26 74
rect 28 72 30 74
rect 23 67 30 72
rect 23 65 26 67
rect 28 65 30 67
rect 23 51 30 65
rect 34 65 41 77
rect 34 63 36 65
rect 38 63 41 65
rect 34 58 41 63
rect 34 56 36 58
rect 38 56 41 58
rect 34 51 41 56
rect 43 73 53 77
rect 43 71 47 73
rect 49 71 53 73
rect 43 66 53 71
rect 43 64 47 66
rect 49 64 53 66
rect 43 51 53 64
rect 55 65 62 77
rect 55 63 58 65
rect 60 63 62 65
rect 55 58 62 63
rect 55 56 58 58
rect 60 56 62 58
rect 55 51 62 56
rect 66 74 73 77
rect 66 72 68 74
rect 70 72 73 74
rect 66 67 73 72
rect 66 65 68 67
rect 70 65 73 67
rect 66 51 73 65
rect 75 65 85 77
rect 75 63 79 65
rect 81 63 85 65
rect 75 57 85 63
rect 75 55 79 57
rect 81 55 85 57
rect 75 51 85 55
rect 87 73 94 77
rect 87 71 90 73
rect 92 71 94 73
rect 87 66 94 71
rect 87 64 90 66
rect 92 64 94 66
rect 87 51 94 64
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 81 34 83
rect 62 85 66 90
rect 94 85 98 90
rect 62 83 63 85
rect 65 83 66 85
rect 62 81 66 83
rect 94 83 95 85
rect 97 83 98 85
rect 94 81 98 83
rect 3 74 7 81
rect 3 72 4 74
rect 6 72 7 74
rect 3 67 7 72
rect 25 74 29 81
rect 25 72 26 74
rect 28 72 29 74
rect 25 67 29 72
rect 3 65 4 67
rect 6 65 7 67
rect 3 63 7 65
rect 25 65 26 67
rect 28 65 29 67
rect 25 63 29 65
rect 78 65 82 67
rect 78 63 79 65
rect 81 63 82 65
rect 6 50 10 51
rect 6 46 27 50
rect 46 47 50 51
rect 6 44 7 46
rect 9 44 10 46
rect 6 37 10 44
rect 21 44 23 46
rect 25 44 27 46
rect 21 34 27 44
rect 37 46 59 47
rect 37 44 39 46
rect 41 44 49 46
rect 51 44 59 46
rect 37 43 59 44
rect 35 36 39 38
rect 35 34 36 36
rect 38 34 39 36
rect 21 30 39 34
rect 53 36 59 43
rect 53 34 55 36
rect 57 34 59 36
rect 53 30 59 34
rect 70 46 74 59
rect 70 44 71 46
rect 73 44 74 46
rect 70 36 74 44
rect 70 34 71 36
rect 73 34 74 36
rect 70 32 74 34
rect 78 57 82 63
rect 78 55 79 57
rect 81 55 82 57
rect 78 26 82 55
rect 35 25 82 26
rect 35 24 58 25
rect 35 22 36 24
rect 38 23 58 24
rect 60 23 68 25
rect 70 23 82 25
rect 38 22 82 23
rect 35 17 42 22
rect 57 18 61 22
rect 35 15 36 17
rect 38 15 42 17
rect 35 13 42 15
rect 46 16 50 18
rect 46 14 47 16
rect 49 14 50 16
rect 57 16 58 18
rect 60 16 61 18
rect 57 14 61 16
rect 67 18 71 22
rect 67 16 68 18
rect 70 16 71 18
rect 46 7 50 14
rect 67 13 71 16
rect 78 16 82 18
rect 78 14 79 16
rect 81 14 82 16
rect 78 7 82 14
rect -2 6 98 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 4 23 6
rect 25 5 84 6
rect 25 4 31 5
rect 1 3 31 4
rect 33 3 63 5
rect 65 4 84 5
rect 86 5 98 6
rect 86 4 95 5
rect 65 3 95 4
rect 97 3 98 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 -2 66 3
rect 94 -2 98 3
<< alu2 >>
rect -2 85 98 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 95 85
rect 97 83 98 85
rect -2 80 98 83
rect -2 5 98 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 95 5
rect 97 3 98 5
rect -2 -2 98 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
rect 93 5 99 7
rect 93 3 95 5
rect 97 3 99 5
rect 93 0 99 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
rect 93 85 99 88
rect 93 83 95 85
rect 97 83 99 85
rect 93 81 99 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polyct0 >>
rect 74 82 76 84
rect 84 82 86 84
<< polyct1 >>
rect 7 44 9 46
rect 23 44 25 46
rect 39 44 41 46
rect 49 44 51 46
rect 71 44 73 46
rect 36 34 38 36
rect 55 34 57 36
rect 71 34 73 36
rect 7 4 9 6
rect 23 4 25 6
rect 84 4 86 6
<< ndifct1 >>
rect 36 22 38 24
rect 36 15 38 17
rect 47 14 49 16
rect 58 23 60 25
rect 58 16 60 18
rect 68 23 70 25
rect 68 16 70 18
rect 79 14 81 16
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< pdifct0 >>
rect 15 63 17 65
rect 15 56 17 58
rect 36 63 38 65
rect 36 56 38 58
rect 47 71 49 73
rect 47 64 49 66
rect 58 63 60 65
rect 58 56 60 58
rect 68 72 70 74
rect 68 65 70 67
rect 90 71 92 73
rect 90 64 92 66
<< pdifct1 >>
rect 4 72 6 74
rect 4 65 6 67
rect 26 72 28 74
rect 26 65 28 67
rect 79 63 81 65
rect 79 55 81 57
<< alu0 >>
rect 72 84 88 85
rect 72 82 74 84
rect 76 82 84 84
rect 86 82 88 84
rect 72 81 88 82
rect 46 74 93 75
rect 46 73 68 74
rect 46 71 47 73
rect 49 72 68 73
rect 70 73 93 74
rect 70 72 90 73
rect 49 71 90 72
rect 92 71 93 73
rect 14 65 18 67
rect 14 63 15 65
rect 17 63 18 65
rect 35 65 39 67
rect 35 63 36 65
rect 38 63 39 65
rect 14 58 18 63
rect 35 58 39 63
rect 46 66 50 71
rect 67 67 71 71
rect 46 64 47 66
rect 49 64 50 66
rect 46 62 50 64
rect 57 65 61 67
rect 57 63 58 65
rect 60 63 61 65
rect 67 65 68 67
rect 70 65 71 67
rect 67 63 71 65
rect 57 58 61 63
rect 14 56 15 58
rect 17 56 36 58
rect 38 56 58 58
rect 60 56 61 58
rect 14 54 61 56
rect 89 66 93 71
rect 89 64 90 66
rect 92 64 93 66
rect 89 62 93 64
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< labels >>
rlabel alu1 8 44 8 44 6 a
rlabel alu1 16 48 16 48 6 a
rlabel alu1 40 20 40 20 6 z
rlabel alu1 24 40 24 40 6 a
rlabel alu1 32 32 32 32 6 a
rlabel alu1 56 24 56 24 6 z
rlabel alu1 64 24 64 24 6 z
rlabel alu1 48 24 48 24 6 z
rlabel alu1 56 36 56 36 6 b
rlabel alu1 48 48 48 48 6 b
rlabel alu1 72 24 72 24 6 z
rlabel alu1 80 48 80 48 6 z
rlabel alu1 72 48 72 48 6 c
rlabel alu2 48 4 48 4 6 vss
rlabel alu2 48 84 48 84 6 vdd
<< end >>
