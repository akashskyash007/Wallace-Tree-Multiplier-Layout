magic
tech scmos
timestamp 1199199122
<< checkpaint >>
rect -1813 -1800 2117 1880
<< ab >>
rect -13 0 317 80
<< alu1 >>
rect -10 69 -6 74
rect -10 67 -9 69
rect -7 67 -6 69
rect -10 53 -6 67
rect -10 51 -9 53
rect -7 51 -6 53
rect -10 37 -6 51
rect -10 35 -9 37
rect -7 35 -6 37
rect -10 21 -6 35
rect -10 19 -9 21
rect -7 19 -6 21
rect -10 12 -6 19
rect -12 8 316 12
rect -10 6 -6 8
<< alu2 >>
rect -13 69 317 70
rect -13 67 -9 69
rect -7 67 317 69
rect -13 66 317 67
rect -13 53 317 54
rect -13 51 -9 53
rect -7 51 317 53
rect -13 50 317 51
rect -13 37 317 38
rect -13 35 -9 37
rect -7 35 317 37
rect -13 34 317 35
rect -13 21 317 22
rect -13 19 -9 21
rect -7 19 3 21
rect 5 19 19 21
rect 21 19 35 21
rect 37 19 51 21
rect 53 19 67 21
rect 69 19 83 21
rect 85 19 99 21
rect 101 19 115 21
rect 117 19 131 21
rect 133 19 147 21
rect 149 19 163 21
rect 165 19 179 21
rect 181 19 195 21
rect 197 19 211 21
rect 213 19 227 21
rect 229 19 243 21
rect 245 19 259 21
rect 261 19 275 21
rect 277 19 291 21
rect 293 19 307 21
rect 309 19 317 21
rect -13 18 317 19
<< alu3 >>
rect 2 61 6 74
rect 2 59 3 61
rect 5 59 6 61
rect 2 45 6 59
rect 2 43 3 45
rect 5 43 6 45
rect 2 29 6 43
rect 2 27 3 29
rect 5 27 6 29
rect 2 21 6 27
rect 2 19 3 21
rect 5 19 6 21
rect 2 13 6 19
rect 2 11 3 13
rect 5 11 6 13
rect 2 6 6 11
rect 18 21 22 74
rect 18 19 19 21
rect 21 19 22 21
rect 18 6 22 19
rect 34 21 38 74
rect 34 19 35 21
rect 37 19 38 21
rect 34 6 38 19
rect 50 21 54 74
rect 50 19 51 21
rect 53 19 54 21
rect 50 6 54 19
rect 66 21 70 74
rect 66 19 67 21
rect 69 19 70 21
rect 66 6 70 19
rect 82 21 86 74
rect 82 19 83 21
rect 85 19 86 21
rect 82 6 86 19
rect 98 21 102 74
rect 98 19 99 21
rect 101 19 102 21
rect 98 6 102 19
rect 114 21 118 74
rect 114 19 115 21
rect 117 19 118 21
rect 114 6 118 19
rect 130 21 134 74
rect 130 19 131 21
rect 133 19 134 21
rect 130 6 134 19
rect 146 21 150 74
rect 146 19 147 21
rect 149 19 150 21
rect 146 6 150 19
rect 162 21 166 74
rect 162 19 163 21
rect 165 19 166 21
rect 162 6 166 19
rect 178 21 182 74
rect 178 19 179 21
rect 181 19 182 21
rect 178 6 182 19
rect 194 21 198 74
rect 194 19 195 21
rect 197 19 198 21
rect 194 6 198 19
rect 210 21 214 74
rect 210 19 211 21
rect 213 19 214 21
rect 210 6 214 19
rect 226 21 230 74
rect 226 19 227 21
rect 229 19 230 21
rect 226 6 230 19
rect 242 21 246 74
rect 242 19 243 21
rect 245 19 246 21
rect 242 6 246 19
rect 258 21 262 74
rect 258 19 259 21
rect 261 19 262 21
rect 258 6 262 19
rect 274 21 278 74
rect 274 19 275 21
rect 277 19 278 21
rect 274 6 278 19
rect 290 21 294 74
rect 290 19 291 21
rect 293 19 294 21
rect 290 6 294 19
rect 306 21 310 74
rect 306 19 307 21
rect 309 19 310 21
rect 306 6 310 19
<< alu4 >>
rect -13 61 317 62
rect -13 59 3 61
rect 5 59 317 61
rect -13 58 317 59
rect -13 45 317 46
rect -13 43 3 45
rect 5 43 317 45
rect -13 42 317 43
rect -13 29 317 30
rect -13 27 3 29
rect 5 27 317 29
rect -13 26 317 27
rect -13 13 317 14
rect -13 11 -5 13
rect -3 11 3 13
rect 5 11 11 13
rect 13 11 27 13
rect 29 11 43 13
rect 45 11 59 13
rect 61 11 75 13
rect 77 11 91 13
rect 93 11 107 13
rect 109 11 123 13
rect 125 11 139 13
rect 141 11 155 13
rect 157 11 171 13
rect 173 11 187 13
rect 189 11 203 13
rect 205 11 219 13
rect 221 11 235 13
rect 237 11 251 13
rect 253 11 267 13
rect 269 11 283 13
rect 285 11 299 13
rect 301 11 317 13
rect -13 10 317 11
<< alu5 >>
rect -6 13 -2 74
rect -6 11 -5 13
rect -3 11 -2 13
rect -6 6 -2 11
rect 10 13 14 74
rect 10 11 11 13
rect 13 11 14 13
rect 10 6 14 11
rect 26 13 30 74
rect 26 11 27 13
rect 29 11 30 13
rect 26 6 30 11
rect 42 13 46 74
rect 42 11 43 13
rect 45 11 46 13
rect 42 6 46 11
rect 58 13 62 74
rect 58 11 59 13
rect 61 11 62 13
rect 58 6 62 11
rect 74 13 78 74
rect 74 11 75 13
rect 77 11 78 13
rect 74 6 78 11
rect 90 13 94 74
rect 90 11 91 13
rect 93 11 94 13
rect 90 6 94 11
rect 106 13 110 74
rect 106 11 107 13
rect 109 11 110 13
rect 106 6 110 11
rect 122 13 126 74
rect 122 11 123 13
rect 125 11 126 13
rect 122 6 126 11
rect 138 13 142 74
rect 138 11 139 13
rect 141 11 142 13
rect 138 6 142 11
rect 154 13 158 74
rect 154 11 155 13
rect 157 11 158 13
rect 154 6 158 11
rect 170 13 174 74
rect 170 11 171 13
rect 173 11 174 13
rect 170 6 174 11
rect 186 13 190 74
rect 186 11 187 13
rect 189 11 190 13
rect 186 6 190 11
rect 202 13 206 74
rect 202 11 203 13
rect 205 11 206 13
rect 202 6 206 11
rect 218 13 222 74
rect 218 11 219 13
rect 221 11 222 13
rect 218 6 222 11
rect 234 13 238 74
rect 234 11 235 13
rect 237 11 238 13
rect 234 6 238 11
rect 250 13 254 74
rect 250 11 251 13
rect 253 11 254 13
rect 250 6 254 11
rect 266 13 270 74
rect 266 11 267 13
rect 269 11 270 13
rect 266 6 270 11
rect 282 13 286 74
rect 282 11 283 13
rect 285 11 286 13
rect 282 6 286 11
rect 298 13 302 74
rect 298 11 299 13
rect 301 11 302 13
rect 298 6 302 11
<< via1 >>
rect -9 67 -7 69
rect -9 51 -7 53
rect -9 35 -7 37
rect -9 19 -7 21
<< via2 >>
rect 3 19 5 21
rect 19 19 21 21
rect 35 19 37 21
rect 51 19 53 21
rect 67 19 69 21
rect 83 19 85 21
rect 99 19 101 21
rect 115 19 117 21
rect 131 19 133 21
rect 147 19 149 21
rect 163 19 165 21
rect 179 19 181 21
rect 195 19 197 21
rect 211 19 213 21
rect 227 19 229 21
rect 243 19 245 21
rect 259 19 261 21
rect 275 19 277 21
rect 291 19 293 21
rect 307 19 309 21
<< via3 >>
rect 3 59 5 61
rect 3 43 5 45
rect 3 27 5 29
rect 3 11 5 13
<< via4 >>
rect -5 11 -3 13
rect 11 11 13 13
rect 27 11 29 13
rect 43 11 45 13
rect 59 11 61 13
rect 75 11 77 13
rect 91 11 93 13
rect 107 11 109 13
rect 123 11 125 13
rect 139 11 141 13
rect 155 11 157 13
rect 171 11 173 13
rect 187 11 189 13
rect 203 11 205 13
rect 219 11 221 13
rect 235 11 237 13
rect 251 11 253 13
rect 267 11 269 13
rect 283 11 285 13
rect 299 11 301 13
<< end >>
