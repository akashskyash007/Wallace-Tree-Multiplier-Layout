magic
tech scmos
timestamp 1199203485
<< ab >>
rect 0 0 136 80
<< nwell >>
rect -5 36 141 88
<< pwell >>
rect -5 -8 141 36
<< poly >>
rect 18 70 20 74
rect 25 70 27 74
rect 35 70 37 74
rect 42 70 44 74
rect 52 70 54 74
rect 59 70 61 74
rect 73 70 75 74
rect 83 70 85 74
rect 93 70 95 74
rect 103 70 105 74
rect 115 70 117 74
rect 125 70 127 74
rect 18 22 20 42
rect 25 39 27 42
rect 35 39 37 42
rect 42 39 44 42
rect 52 39 54 42
rect 25 37 38 39
rect 32 35 34 37
rect 36 35 38 37
rect 32 33 38 35
rect 42 37 54 39
rect 59 39 61 42
rect 73 39 75 42
rect 83 39 85 42
rect 93 39 95 42
rect 59 37 68 39
rect 32 30 34 33
rect 42 30 44 37
rect 52 30 54 37
rect 62 35 64 37
rect 66 35 68 37
rect 62 33 68 35
rect 72 37 79 39
rect 83 37 99 39
rect 72 35 75 37
rect 77 35 79 37
rect 72 33 79 35
rect 93 35 95 37
rect 97 35 99 37
rect 93 33 99 35
rect 62 30 64 33
rect 72 30 74 33
rect 103 30 105 42
rect 115 39 117 42
rect 125 39 127 42
rect 109 37 127 39
rect 109 35 111 37
rect 113 35 127 37
rect 109 33 127 35
rect 115 30 117 33
rect 125 30 127 33
rect 17 20 23 22
rect 17 18 19 20
rect 21 18 23 20
rect 17 16 23 18
rect 21 8 23 16
rect 32 12 34 16
rect 42 8 44 16
rect 52 11 54 16
rect 62 11 64 16
rect 21 6 44 8
rect 72 8 74 16
rect 103 8 105 16
rect 115 11 117 16
rect 125 11 127 16
rect 72 6 105 8
<< ndif >>
rect 27 22 32 30
rect 25 20 32 22
rect 25 18 27 20
rect 29 18 32 20
rect 25 16 32 18
rect 34 28 42 30
rect 34 26 37 28
rect 39 26 42 28
rect 34 16 42 26
rect 44 28 52 30
rect 44 26 47 28
rect 49 26 52 28
rect 44 16 52 26
rect 54 28 62 30
rect 54 26 57 28
rect 59 26 62 28
rect 54 16 62 26
rect 64 21 72 30
rect 64 19 67 21
rect 69 19 72 21
rect 64 16 72 19
rect 74 16 82 30
rect 96 28 103 30
rect 96 26 98 28
rect 100 26 103 28
rect 96 21 103 26
rect 96 19 98 21
rect 100 19 103 21
rect 96 16 103 19
rect 105 27 115 30
rect 105 25 109 27
rect 111 25 115 27
rect 105 20 115 25
rect 105 18 109 20
rect 111 18 115 20
rect 105 16 115 18
rect 117 28 125 30
rect 117 26 120 28
rect 122 26 125 28
rect 117 21 125 26
rect 117 19 120 21
rect 122 19 125 21
rect 117 16 125 19
rect 127 27 134 30
rect 127 25 130 27
rect 132 25 134 27
rect 127 20 134 25
rect 127 18 130 20
rect 132 18 134 20
rect 127 16 134 18
rect 76 14 82 16
rect 76 12 78 14
rect 80 12 82 14
rect 76 10 82 12
<< pdif >>
rect 13 55 18 70
rect 11 53 18 55
rect 11 51 13 53
rect 15 51 18 53
rect 11 46 18 51
rect 11 44 13 46
rect 15 44 18 46
rect 11 42 18 44
rect 20 42 25 70
rect 27 68 35 70
rect 27 66 30 68
rect 32 66 35 68
rect 27 42 35 66
rect 37 42 42 70
rect 44 61 52 70
rect 44 59 47 61
rect 49 59 52 61
rect 44 46 52 59
rect 44 44 47 46
rect 49 44 52 46
rect 44 42 52 44
rect 54 42 59 70
rect 61 68 73 70
rect 61 66 66 68
rect 68 66 73 68
rect 61 42 73 66
rect 75 46 83 70
rect 75 44 78 46
rect 80 44 83 46
rect 75 42 83 44
rect 85 61 93 70
rect 85 59 88 61
rect 90 59 93 61
rect 85 42 93 59
rect 95 46 103 70
rect 95 44 98 46
rect 100 44 103 46
rect 95 42 103 44
rect 105 68 115 70
rect 105 66 109 68
rect 111 66 115 68
rect 105 61 115 66
rect 105 59 109 61
rect 111 59 115 61
rect 105 42 115 59
rect 117 54 125 70
rect 117 52 120 54
rect 122 52 125 54
rect 117 46 125 52
rect 117 44 120 46
rect 122 44 125 46
rect 117 42 125 44
rect 127 68 134 70
rect 127 66 130 68
rect 132 66 134 68
rect 127 61 134 66
rect 127 59 130 61
rect 132 59 134 61
rect 127 42 134 59
<< alu1 >>
rect -2 81 138 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 138 81
rect -2 68 138 79
rect 26 61 92 62
rect 26 59 47 61
rect 49 59 88 61
rect 90 59 92 61
rect 26 58 92 59
rect 10 53 16 55
rect 10 51 13 53
rect 15 51 16 53
rect 10 46 16 51
rect 26 46 30 58
rect 10 44 13 46
rect 15 44 30 46
rect 10 42 30 44
rect 26 29 30 42
rect 26 28 41 29
rect 26 26 37 28
rect 39 26 41 28
rect 26 25 41 26
rect 73 37 79 38
rect 73 35 75 37
rect 77 35 79 37
rect 73 30 79 35
rect 65 26 79 30
rect 106 38 110 47
rect 93 37 115 38
rect 93 35 95 37
rect 97 35 111 37
rect 113 35 115 37
rect 93 34 115 35
rect -2 1 138 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 138 1
rect -2 -2 138 -1
<< ptie >>
rect 0 1 136 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 136 1
rect 0 -3 136 -1
<< ntie >>
rect 0 81 136 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 136 81
rect 0 77 136 79
<< nmos >>
rect 32 16 34 30
rect 42 16 44 30
rect 52 16 54 30
rect 62 16 64 30
rect 72 16 74 30
rect 103 16 105 30
rect 115 16 117 30
rect 125 16 127 30
<< pmos >>
rect 18 42 20 70
rect 25 42 27 70
rect 35 42 37 70
rect 42 42 44 70
rect 52 42 54 70
rect 59 42 61 70
rect 73 42 75 70
rect 83 42 85 70
rect 93 42 95 70
rect 103 42 105 70
rect 115 42 117 70
rect 125 42 127 70
<< polyct0 >>
rect 34 35 36 37
rect 64 35 66 37
rect 19 18 21 20
<< polyct1 >>
rect 75 35 77 37
rect 95 35 97 37
rect 111 35 113 37
<< ndifct0 >>
rect 27 18 29 20
rect 47 26 49 28
rect 57 26 59 28
rect 67 19 69 21
rect 98 26 100 28
rect 98 19 100 21
rect 109 25 111 27
rect 109 18 111 20
rect 120 26 122 28
rect 120 19 122 21
rect 130 25 132 27
rect 130 18 132 20
rect 78 12 80 14
<< ndifct1 >>
rect 37 26 39 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
<< pdifct0 >>
rect 30 66 32 68
rect 47 44 49 46
rect 66 66 68 68
rect 78 44 80 46
rect 98 44 100 46
rect 109 66 111 68
rect 109 59 111 61
rect 120 52 122 54
rect 120 44 122 46
rect 130 66 132 68
rect 130 59 132 61
<< pdifct1 >>
rect 13 51 15 53
rect 13 44 15 46
rect 47 59 49 61
rect 88 59 90 61
<< alu0 >>
rect 28 66 30 68
rect 32 66 34 68
rect 28 65 34 66
rect 64 66 66 68
rect 68 66 70 68
rect 64 65 70 66
rect 107 66 109 68
rect 111 66 113 68
rect 107 61 113 66
rect 107 59 109 61
rect 111 59 113 61
rect 107 58 113 59
rect 128 66 130 68
rect 132 66 134 68
rect 128 61 134 66
rect 128 59 130 61
rect 132 59 134 61
rect 128 58 134 59
rect 119 54 123 56
rect 37 52 120 54
rect 122 52 123 54
rect 37 50 123 52
rect 37 39 41 50
rect 45 46 51 47
rect 45 44 47 46
rect 49 44 58 46
rect 45 42 58 44
rect 33 37 41 39
rect 33 35 34 37
rect 36 35 50 37
rect 33 33 50 35
rect 46 28 50 33
rect 46 26 47 28
rect 49 26 50 28
rect 46 24 50 26
rect 54 29 58 42
rect 63 37 67 50
rect 76 46 82 47
rect 96 46 102 47
rect 76 44 78 46
rect 80 44 98 46
rect 100 44 102 46
rect 76 42 102 44
rect 63 35 64 37
rect 66 35 67 37
rect 63 33 67 35
rect 54 28 61 29
rect 54 26 57 28
rect 59 26 61 28
rect 83 26 87 42
rect 119 46 123 50
rect 119 44 120 46
rect 122 44 123 46
rect 97 28 101 30
rect 97 26 98 28
rect 100 26 101 28
rect 54 25 61 26
rect 83 22 101 26
rect 65 21 87 22
rect 17 20 67 21
rect 17 18 19 20
rect 21 18 27 20
rect 29 19 67 20
rect 69 19 87 21
rect 29 18 87 19
rect 97 21 101 22
rect 97 19 98 21
rect 100 19 101 21
rect 17 17 70 18
rect 97 17 101 19
rect 108 27 112 29
rect 108 25 109 27
rect 111 25 112 27
rect 108 20 112 25
rect 108 18 109 20
rect 111 18 112 20
rect 76 14 82 15
rect 76 12 78 14
rect 80 12 82 14
rect 86 12 92 15
rect 108 12 112 18
rect 119 28 123 44
rect 119 26 120 28
rect 122 26 123 28
rect 119 21 123 26
rect 119 19 120 21
rect 122 19 123 21
rect 119 17 123 19
rect 129 27 133 29
rect 129 25 130 27
rect 132 25 133 27
rect 129 20 133 25
rect 129 18 130 20
rect 132 18 133 20
rect 129 12 133 18
<< labels >>
rlabel alu0 48 30 48 30 6 bn
rlabel alu0 39 43 39 43 6 bn
rlabel alu0 43 19 43 19 6 an
rlabel alu0 65 43 65 43 6 bn
rlabel alu0 76 20 76 20 6 an
rlabel alu0 99 23 99 23 6 an
rlabel alu0 89 44 89 44 6 an
rlabel alu0 99 44 99 44 6 an
rlabel alu0 121 36 121 36 6 bn
rlabel alu1 28 40 28 40 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 52 60 52 60 6 z
rlabel alu1 60 60 60 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 68 6 68 6 6 vss
rlabel alu1 68 28 68 28 6 a
rlabel alu1 100 36 100 36 6 b
rlabel alu1 76 32 76 32 6 a
rlabel alu1 76 60 76 60 6 z
rlabel alu1 84 60 84 60 6 z
rlabel alu1 68 60 68 60 6 z
rlabel alu1 68 74 68 74 6 vdd
rlabel alu1 108 40 108 40 6 b
<< end >>
