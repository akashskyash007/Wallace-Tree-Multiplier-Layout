magic
tech scmos
timestamp 1199202912
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 9 34 11 43
rect 16 40 18 43
rect 26 40 28 43
rect 16 38 28 40
rect 21 37 28 38
rect 21 35 24 37
rect 26 35 28 37
rect 9 32 17 34
rect 9 31 13 32
rect 11 30 13 31
rect 15 30 17 32
rect 11 28 17 30
rect 21 33 28 35
rect 11 25 13 28
rect 21 25 23 33
rect 33 31 35 43
rect 33 29 39 31
rect 33 27 35 29
rect 37 27 39 29
rect 33 25 39 27
rect 11 6 13 10
rect 21 6 23 10
<< ndif >>
rect 3 14 11 25
rect 3 12 6 14
rect 8 12 11 14
rect 3 10 11 12
rect 13 21 21 25
rect 13 19 16 21
rect 18 19 21 21
rect 13 10 21 19
rect 23 21 31 25
rect 23 19 26 21
rect 28 19 31 21
rect 23 14 31 19
rect 23 12 26 14
rect 28 12 31 14
rect 23 10 31 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 43 9 59
rect 11 43 16 70
rect 18 54 26 70
rect 18 52 21 54
rect 23 52 26 54
rect 18 47 26 52
rect 18 45 21 47
rect 23 45 26 47
rect 18 43 26 45
rect 28 43 33 70
rect 35 68 42 70
rect 35 66 38 68
rect 40 66 42 68
rect 35 61 42 66
rect 35 59 38 61
rect 40 59 42 61
rect 35 43 42 59
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 18 54 24 56
rect 18 52 21 54
rect 23 52 24 54
rect 18 47 24 52
rect 18 46 21 47
rect 2 45 21 46
rect 23 45 24 47
rect 2 42 24 45
rect 2 22 6 42
rect 34 38 39 47
rect 22 37 39 38
rect 22 35 24 37
rect 26 35 39 37
rect 22 34 39 35
rect 12 32 16 34
rect 12 30 13 32
rect 15 30 16 32
rect 12 29 39 30
rect 12 27 35 29
rect 37 27 39 29
rect 12 26 39 27
rect 2 21 20 22
rect 2 19 16 21
rect 18 19 20 21
rect 2 18 20 19
rect 34 17 39 26
rect -2 1 50 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 11 10 13 25
rect 21 10 23 25
<< pmos >>
rect 9 43 11 70
rect 16 43 18 70
rect 26 43 28 70
rect 33 43 35 70
<< polyct1 >>
rect 24 35 26 37
rect 13 30 15 32
rect 35 27 37 29
<< ndifct0 >>
rect 6 12 8 14
rect 26 19 28 21
rect 26 12 28 14
<< ndifct1 >>
rect 16 19 18 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 38 66 40 68
rect 38 59 40 61
<< pdifct1 >>
rect 21 52 23 54
rect 21 45 23 47
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 36 66 38 68
rect 40 66 42 68
rect 36 61 42 66
rect 36 59 38 61
rect 40 59 42 61
rect 36 58 42 59
rect 24 21 30 22
rect 24 19 26 21
rect 28 19 30 21
rect 4 14 10 15
rect 4 12 6 14
rect 8 12 10 14
rect 24 14 30 19
rect 24 12 26 14
rect 28 12 30 14
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 28 28 28 6 a
rlabel alu1 28 36 28 36 6 b
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 36 24 36 24 6 a
rlabel alu1 36 40 36 40 6 b
<< end >>
