magic
tech scmos
timestamp 1199470660
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 13 85 15 89
rect 21 85 23 89
rect 33 85 35 90
rect 45 85 47 90
rect 57 85 59 90
rect 13 53 15 65
rect 21 62 23 65
rect 33 62 35 65
rect 21 60 27 62
rect 13 51 21 53
rect 13 50 17 51
rect 11 49 17 50
rect 19 49 21 51
rect 11 47 21 49
rect 25 51 27 60
rect 33 60 41 62
rect 33 58 37 60
rect 39 58 41 60
rect 33 56 41 58
rect 25 49 41 51
rect 11 33 13 47
rect 25 39 27 49
rect 35 47 37 49
rect 39 47 41 49
rect 35 45 41 47
rect 23 36 27 39
rect 45 42 47 65
rect 57 62 59 65
rect 51 60 59 62
rect 51 58 53 60
rect 55 58 59 60
rect 51 56 59 58
rect 45 40 53 42
rect 45 38 49 40
rect 51 38 53 40
rect 35 36 53 38
rect 23 33 25 36
rect 35 33 37 36
rect 57 33 59 56
rect 11 19 13 24
rect 23 19 25 24
rect 35 19 37 24
rect 57 19 59 24
<< ndif >>
rect 6 30 11 33
rect 3 28 11 30
rect 3 26 5 28
rect 7 26 11 28
rect 3 24 11 26
rect 13 31 23 33
rect 13 29 17 31
rect 19 29 23 31
rect 13 24 23 29
rect 25 31 35 33
rect 25 29 29 31
rect 31 29 35 31
rect 25 24 35 29
rect 37 24 57 33
rect 59 31 67 33
rect 59 29 63 31
rect 65 29 67 31
rect 59 27 67 29
rect 59 24 64 27
rect 39 11 55 24
rect 39 9 41 11
rect 43 9 51 11
rect 53 9 55 11
rect 39 7 55 9
<< pdif >>
rect 49 91 55 93
rect 49 89 51 91
rect 53 89 55 91
rect 49 85 55 89
rect 4 81 13 85
rect 4 79 7 81
rect 9 79 13 81
rect 4 65 13 79
rect 15 65 21 85
rect 23 81 33 85
rect 23 79 27 81
rect 29 79 33 81
rect 23 65 33 79
rect 35 81 45 85
rect 35 79 39 81
rect 41 79 45 81
rect 35 73 45 79
rect 35 71 39 73
rect 41 71 45 73
rect 35 65 45 71
rect 47 65 57 85
rect 59 79 64 85
rect 59 77 67 79
rect 59 75 63 77
rect 65 75 67 77
rect 59 69 67 75
rect 59 67 63 69
rect 65 67 67 69
rect 59 65 67 67
<< alu1 >>
rect -2 95 72 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 72 95
rect -2 91 72 93
rect -2 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 6 81 10 88
rect 6 79 7 81
rect 9 79 10 81
rect 6 77 10 79
rect 18 81 33 83
rect 18 79 27 81
rect 29 79 33 81
rect 18 78 33 79
rect 38 81 42 83
rect 38 79 39 81
rect 41 79 42 81
rect 18 73 22 78
rect 8 67 22 73
rect 38 73 42 79
rect 38 72 39 73
rect 28 71 39 72
rect 41 71 42 73
rect 28 68 42 71
rect 8 43 12 67
rect 28 53 32 68
rect 48 62 52 83
rect 62 77 66 79
rect 62 75 63 77
rect 65 75 66 77
rect 62 69 66 75
rect 62 67 63 69
rect 65 67 66 69
rect 36 60 57 62
rect 36 58 37 60
rect 39 58 53 60
rect 55 58 57 60
rect 36 56 57 58
rect 16 51 32 53
rect 62 51 66 67
rect 16 49 17 51
rect 19 49 32 51
rect 16 47 32 49
rect 8 37 22 43
rect 16 31 22 37
rect 4 28 8 30
rect 4 26 5 28
rect 7 26 8 28
rect 16 29 17 31
rect 19 29 22 31
rect 16 27 22 29
rect 28 31 32 47
rect 28 29 29 31
rect 31 29 32 31
rect 28 27 32 29
rect 36 49 66 51
rect 36 47 37 49
rect 39 47 66 49
rect 4 22 8 26
rect 36 22 40 47
rect 4 18 40 22
rect 47 40 53 42
rect 47 38 49 40
rect 51 38 53 40
rect 47 22 53 38
rect 62 31 66 47
rect 62 29 63 31
rect 65 29 66 31
rect 62 27 66 29
rect 47 18 63 22
rect -2 11 72 12
rect -2 9 41 11
rect 43 9 51 11
rect 53 9 72 11
rect -2 7 72 9
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 72 7
rect -2 0 72 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 11 24 13 33
rect 23 24 25 33
rect 35 24 37 33
rect 57 24 59 33
<< pmos >>
rect 13 65 15 85
rect 21 65 23 85
rect 33 65 35 85
rect 45 65 47 85
rect 57 65 59 85
<< polyct1 >>
rect 17 49 19 51
rect 37 58 39 60
rect 37 47 39 49
rect 53 58 55 60
rect 49 38 51 40
<< ndifct1 >>
rect 5 26 7 28
rect 17 29 19 31
rect 29 29 31 31
rect 63 29 65 31
rect 41 9 43 11
rect 51 9 53 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 51 89 53 91
rect 7 79 9 81
rect 27 79 29 81
rect 39 79 41 81
rect 39 71 41 73
rect 63 75 65 77
rect 63 67 65 69
<< labels >>
rlabel alu1 6 24 6 24 6 bn
rlabel alu1 20 35 20 35 6 z
rlabel alu1 10 55 10 55 6 z
rlabel alu1 20 75 20 75 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 24 50 24 50 6 an
rlabel alu1 30 49 30 49 6 an
rlabel alu1 30 80 30 80 6 z
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 50 30 50 30 6 a
rlabel alu1 40 60 40 60 6 b
rlabel alu1 50 70 50 70 6 b
rlabel alu1 40 75 40 75 6 an
rlabel alu1 60 20 60 20 6 a
rlabel alu1 51 49 51 49 6 bn
rlabel alu1 64 53 64 53 6 bn
<< end >>
