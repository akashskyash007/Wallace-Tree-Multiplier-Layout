magic
tech scmos
timestamp 1199203653
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 18 70 20 74
rect 25 70 27 74
rect 36 70 38 74
rect 43 70 45 74
rect 2 61 8 63
rect 2 59 4 61
rect 6 59 8 61
rect 2 57 11 59
rect 9 54 11 57
rect 54 61 56 66
rect 54 46 56 50
rect 54 44 64 46
rect 9 30 11 43
rect 18 40 20 43
rect 15 38 21 40
rect 15 36 17 38
rect 19 36 21 38
rect 15 34 21 36
rect 25 30 27 43
rect 36 39 38 43
rect 43 40 45 43
rect 54 42 60 44
rect 62 42 64 44
rect 54 40 64 42
rect 9 28 27 30
rect 31 37 38 39
rect 31 35 33 37
rect 35 35 38 37
rect 31 33 38 35
rect 42 38 64 40
rect 9 25 11 28
rect 21 25 23 28
rect 31 25 33 33
rect 42 30 44 38
rect 51 32 57 34
rect 51 30 53 32
rect 55 30 57 32
rect 9 15 11 19
rect 51 28 57 30
rect 52 24 54 28
rect 61 26 63 38
rect 21 8 23 13
rect 31 9 33 14
rect 42 13 44 18
rect 61 16 63 20
rect 52 6 54 10
<< ndif >>
rect 35 28 42 30
rect 35 26 37 28
rect 39 26 42 28
rect 35 25 42 26
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 19 21 25
rect 13 17 21 19
rect 13 15 15 17
rect 17 15 21 17
rect 13 13 21 15
rect 23 21 31 25
rect 23 19 26 21
rect 28 19 31 21
rect 23 14 31 19
rect 33 18 42 25
rect 44 24 49 30
rect 56 24 61 26
rect 44 22 52 24
rect 44 20 47 22
rect 49 20 52 22
rect 44 18 52 20
rect 33 14 38 18
rect 23 13 28 14
rect 47 10 52 18
rect 54 20 61 24
rect 63 24 70 26
rect 63 22 66 24
rect 68 22 70 24
rect 63 20 70 22
rect 54 14 59 20
rect 54 12 62 14
rect 54 10 58 12
rect 60 10 62 12
rect 56 8 62 10
<< pdif >>
rect 11 65 18 70
rect 11 63 13 65
rect 15 63 18 65
rect 11 61 18 63
rect 13 54 18 61
rect 4 49 9 54
rect 2 47 9 49
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 43 18 54
rect 20 43 25 70
rect 27 47 36 70
rect 27 45 31 47
rect 33 45 36 47
rect 27 43 36 45
rect 38 43 43 70
rect 45 63 52 70
rect 45 61 48 63
rect 50 61 52 63
rect 45 50 54 61
rect 56 56 61 61
rect 56 54 63 56
rect 56 52 59 54
rect 61 52 63 54
rect 56 50 63 52
rect 45 43 52 50
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 61 7 63
rect 2 59 4 61
rect 6 59 7 61
rect 2 58 7 59
rect 2 54 14 58
rect 10 49 14 54
rect 29 47 35 48
rect 29 45 31 47
rect 33 45 46 47
rect 29 42 46 45
rect 42 30 46 42
rect 35 28 46 30
rect 66 47 70 55
rect 58 44 70 47
rect 58 42 60 44
rect 62 42 70 44
rect 58 41 70 42
rect 35 26 37 28
rect 39 26 46 28
rect 35 25 41 26
rect -2 10 58 12
rect 60 10 74 12
rect -2 1 74 10
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 9 19 11 25
rect 21 13 23 25
rect 31 14 33 25
rect 42 18 44 30
rect 52 10 54 24
rect 61 20 63 26
<< pmos >>
rect 9 43 11 54
rect 18 43 20 70
rect 25 43 27 70
rect 36 43 38 70
rect 43 43 45 70
rect 54 50 56 61
<< polyct0 >>
rect 17 36 19 38
rect 33 35 35 37
rect 53 30 55 32
<< polyct1 >>
rect 4 59 6 61
rect 60 42 62 44
<< ndifct0 >>
rect 4 21 6 23
rect 15 15 17 17
rect 26 19 28 21
rect 47 20 49 22
rect 66 22 68 24
<< ndifct1 >>
rect 37 26 39 28
rect 58 10 60 12
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 13 63 15 65
rect 4 45 6 47
rect 48 61 50 63
rect 59 52 61 54
<< pdifct1 >>
rect 31 45 33 47
<< alu0 >>
rect 11 65 17 68
rect 11 63 13 65
rect 15 63 17 65
rect 11 62 17 63
rect 47 63 51 68
rect 47 61 48 63
rect 50 61 51 63
rect 47 59 51 61
rect 18 54 63 55
rect 18 52 59 54
rect 61 52 63 54
rect 18 51 63 52
rect 3 47 7 49
rect 3 45 4 47
rect 6 45 7 47
rect 3 30 7 45
rect 18 39 22 51
rect 15 38 22 39
rect 15 36 17 38
rect 19 36 22 38
rect 15 35 22 36
rect 27 37 37 38
rect 27 35 33 37
rect 35 35 37 37
rect 27 34 37 35
rect 27 30 31 34
rect 3 26 31 30
rect 50 33 54 51
rect 50 32 69 33
rect 50 30 53 32
rect 55 30 69 32
rect 50 29 69 30
rect 3 23 7 26
rect 65 24 69 29
rect 3 21 4 23
rect 6 21 7 23
rect 45 22 51 23
rect 3 19 7 21
rect 24 21 47 22
rect 24 19 26 21
rect 28 20 47 21
rect 49 20 51 22
rect 65 22 66 24
rect 68 22 69 24
rect 65 20 69 22
rect 28 19 51 20
rect 14 17 18 19
rect 24 18 51 19
rect 14 15 15 17
rect 17 15 18 17
rect 14 12 18 15
rect 56 12 62 13
<< labels >>
rlabel alu0 5 34 5 34 6 bn
rlabel alu0 20 45 20 45 6 an
rlabel alu0 37 20 37 20 6 n3
rlabel alu0 32 36 32 36 6 bn
rlabel alu0 67 26 67 26 6 an
rlabel alu0 59 31 59 31 6 an
rlabel alu0 40 53 40 53 6 an
rlabel alu1 12 52 12 52 6 b
rlabel alu1 4 60 4 60 6 b
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 44 40 44 40 6 z
rlabel alu1 36 44 36 44 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 44 60 44 6 a
rlabel alu1 68 48 68 48 6 a
<< end >>
