magic
tech scmos
timestamp 1199543817
<< ab >>
rect 0 0 10 100
<< nwell >>
rect -2 48 12 104
<< pwell >>
rect -2 -4 12 48
<< alu1 >>
rect -2 88 12 100
rect -2 0 12 12
<< labels >>
rlabel alu1 5 6 5 6 6 vss
rlabel alu1 5 94 5 94 6 vdd
<< end >>
