magic
tech scmos
timestamp 1199541824
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -5 48 55 105
<< pwell >>
rect -5 -5 55 48
<< poly >>
rect 23 94 25 98
rect 35 94 37 98
rect 11 75 13 79
rect 11 53 13 56
rect 11 51 19 53
rect 11 49 15 51
rect 17 49 19 51
rect 11 47 19 49
rect 23 43 25 55
rect 35 43 37 55
rect 3 41 37 43
rect 3 39 5 41
rect 7 39 37 41
rect 3 37 37 39
rect 11 31 19 33
rect 11 29 15 31
rect 17 29 19 31
rect 11 27 19 29
rect 11 24 13 27
rect 23 25 25 37
rect 35 25 37 37
rect 11 10 13 14
rect 23 2 25 6
rect 35 2 37 6
<< ndif >>
rect 18 24 23 25
rect 3 21 11 24
rect 3 19 5 21
rect 7 19 11 21
rect 3 14 11 19
rect 13 14 23 24
rect 15 11 23 14
rect 15 9 17 11
rect 19 9 23 11
rect 15 6 23 9
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 6 35 19
rect 37 21 45 25
rect 37 19 41 21
rect 43 19 45 21
rect 37 11 45 19
rect 37 9 41 11
rect 43 9 45 11
rect 37 6 45 9
<< pdif >>
rect 15 91 23 94
rect 15 89 17 91
rect 19 89 23 91
rect 15 75 23 89
rect 3 71 11 75
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 56 11 59
rect 13 56 23 75
rect 18 55 23 56
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 91 45 94
rect 37 89 41 91
rect 43 89 45 91
rect 37 81 45 89
rect 37 79 41 81
rect 43 79 45 81
rect 37 71 45 79
rect 37 69 41 71
rect 43 69 45 71
rect 37 61 45 69
rect 37 59 41 61
rect 43 59 45 61
rect 37 55 45 59
<< alu1 >>
rect -2 95 52 100
rect -2 93 5 95
rect 7 93 52 95
rect -2 91 52 93
rect -2 89 17 91
rect 19 89 41 91
rect 43 89 52 91
rect -2 88 52 89
rect 4 85 8 88
rect 4 83 5 85
rect 7 83 8 85
rect 4 81 8 83
rect 4 71 8 73
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 4 59 5 61
rect 7 59 8 61
rect 4 41 8 59
rect 18 52 22 83
rect 13 51 22 52
rect 13 49 15 51
rect 17 49 22 51
rect 13 48 22 49
rect 4 39 5 41
rect 7 39 8 41
rect 4 21 8 39
rect 18 32 22 48
rect 13 31 22 32
rect 13 29 15 31
rect 17 29 22 31
rect 13 28 22 29
rect 4 19 5 21
rect 7 19 8 21
rect 4 17 8 19
rect 18 17 22 28
rect 28 81 32 83
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 28 21 32 59
rect 40 81 44 88
rect 40 79 41 81
rect 43 79 44 81
rect 40 71 44 79
rect 40 69 41 71
rect 43 69 44 71
rect 40 61 44 69
rect 40 59 41 61
rect 43 59 44 61
rect 40 57 44 59
rect 28 19 29 21
rect 31 19 32 21
rect 28 17 32 19
rect 40 21 44 23
rect 40 19 41 21
rect 43 19 44 21
rect 40 12 44 19
rect -2 11 52 12
rect -2 9 17 11
rect 19 9 41 11
rect 43 9 52 11
rect -2 0 52 9
<< ntie >>
rect 3 95 9 97
rect 3 93 5 95
rect 7 93 9 95
rect 3 85 9 93
rect 3 83 5 85
rect 7 83 9 85
rect 3 81 9 83
<< nmos >>
rect 11 14 13 24
rect 23 6 25 25
rect 35 6 37 25
<< pmos >>
rect 11 56 13 75
rect 23 55 25 94
rect 35 55 37 94
<< polyct1 >>
rect 15 49 17 51
rect 5 39 7 41
rect 15 29 17 31
<< ndifct1 >>
rect 5 19 7 21
rect 17 9 19 11
rect 29 19 31 21
rect 41 19 43 21
rect 41 9 43 11
<< ntiect1 >>
rect 5 93 7 95
rect 5 83 7 85
<< pdifct1 >>
rect 17 89 19 91
rect 5 69 7 71
rect 5 59 7 61
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
rect 41 89 43 91
rect 41 79 43 81
rect 41 69 43 71
rect 41 59 43 61
<< labels >>
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 50 30 50 6 q
rlabel alu1 20 50 20 50 6 i
rlabel alu1 25 94 25 94 6 vdd
<< end >>
