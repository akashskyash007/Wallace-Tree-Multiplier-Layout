magic
tech scmos
timestamp 1199202038
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 38 11 42
rect 19 38 21 42
rect 29 39 31 42
rect 9 36 22 38
rect 9 34 18 36
rect 20 34 22 36
rect 9 32 22 34
rect 26 37 32 39
rect 26 35 28 37
rect 30 35 32 37
rect 26 33 32 35
rect 9 29 11 32
rect 19 29 21 32
rect 29 29 31 33
rect 9 10 11 15
rect 19 10 21 15
rect 29 10 31 15
<< ndif >>
rect 2 27 9 29
rect 2 25 4 27
rect 6 25 9 27
rect 2 19 9 25
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 21 19 29
rect 11 19 14 21
rect 16 19 19 21
rect 11 15 19 19
rect 21 19 29 29
rect 21 17 24 19
rect 26 17 29 19
rect 21 15 29 17
rect 31 27 38 29
rect 31 25 34 27
rect 36 25 38 27
rect 31 20 38 25
rect 31 18 34 20
rect 36 18 38 20
rect 31 15 38 18
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 55 36 70
rect 31 53 38 55
rect 31 51 34 53
rect 36 51 38 53
rect 31 46 38 51
rect 31 44 34 46
rect 36 44 38 46
rect 31 42 38 44
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 37 6 50
rect 17 42 30 46
rect 26 39 30 42
rect 2 33 14 37
rect 10 23 14 33
rect 26 37 31 39
rect 26 35 28 37
rect 30 35 31 37
rect 26 33 31 35
rect 10 21 17 23
rect 10 19 14 21
rect 16 19 17 21
rect 10 17 17 19
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 15 11 29
rect 19 15 21 29
rect 29 15 31 29
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
<< polyct0 >>
rect 18 34 20 36
<< polyct1 >>
rect 28 35 30 37
<< ndifct0 >>
rect 4 25 6 27
rect 4 17 6 19
rect 24 17 26 19
rect 34 25 36 27
rect 34 18 36 20
<< ndifct1 >>
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 66 26 68
rect 24 59 26 61
rect 34 51 36 53
rect 34 44 36 46
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 61 28 66
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 33 53 38 55
rect 33 51 34 53
rect 36 51 38 53
rect 33 46 38 51
rect 33 44 34 46
rect 36 44 38 46
rect 33 42 38 44
rect 3 27 7 29
rect 3 25 4 27
rect 6 25 7 27
rect 3 19 7 25
rect 3 17 4 19
rect 6 17 7 19
rect 17 36 21 38
rect 17 34 18 36
rect 20 34 21 36
rect 17 30 21 34
rect 34 30 38 42
rect 17 27 38 30
rect 17 26 34 27
rect 32 25 34 26
rect 36 25 38 27
rect 23 19 27 21
rect 23 17 24 19
rect 26 17 27 19
rect 32 20 38 25
rect 32 18 34 20
rect 36 18 38 20
rect 32 17 38 18
rect 3 12 7 17
rect 23 12 27 17
<< labels >>
rlabel alu0 19 32 19 32 6 an
rlabel alu0 36 36 36 36 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 36 28 36 6 a
rlabel alu1 20 44 20 44 6 a
rlabel alu1 20 74 20 74 6 vdd
<< end >>
