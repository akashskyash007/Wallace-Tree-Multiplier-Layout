magic
tech scmos
timestamp 1199543067
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 35 94 37 98
rect 47 94 49 98
rect 57 94 59 98
rect 11 84 13 88
rect 23 85 25 89
rect 11 43 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 21 51 25 53
rect 33 51 37 53
rect 21 43 23 51
rect 33 43 35 51
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 35 43
rect 27 39 29 41
rect 31 39 35 41
rect 47 43 49 55
rect 57 43 59 55
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 27 37 35 39
rect 11 34 13 37
rect 21 34 23 37
rect 33 34 35 37
rect 45 37 53 39
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 45 34 47 37
rect 57 34 59 37
rect 11 12 13 16
rect 21 13 23 17
rect 33 13 35 17
rect 45 13 47 17
rect 57 12 59 16
<< ndif >>
rect 3 16 11 34
rect 13 17 21 34
rect 23 21 33 34
rect 23 19 27 21
rect 29 19 33 21
rect 23 17 33 19
rect 35 21 45 34
rect 35 19 39 21
rect 41 19 45 21
rect 35 17 45 19
rect 47 17 57 34
rect 13 16 18 17
rect 3 11 9 16
rect 49 16 57 17
rect 59 21 67 34
rect 59 19 63 21
rect 65 19 67 21
rect 59 16 67 19
rect 49 11 55 16
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 30 85 35 94
rect 15 84 23 85
rect 3 81 11 84
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 56 23 84
rect 25 81 35 85
rect 25 79 29 81
rect 31 79 35 81
rect 25 56 35 79
rect 37 71 47 94
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 13 55 18 56
rect 42 55 47 56
rect 49 55 57 94
rect 59 81 67 94
rect 59 79 63 81
rect 65 79 67 81
rect 59 55 67 79
<< alu1 >>
rect -2 91 72 100
rect -2 89 17 91
rect 19 89 72 91
rect -2 88 72 89
rect 3 81 67 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 79 63 81
rect 65 79 67 81
rect 3 78 67 79
rect 8 41 12 73
rect 8 39 9 41
rect 11 39 12 41
rect 8 17 12 39
rect 18 41 22 73
rect 18 39 19 41
rect 21 39 22 41
rect 18 27 22 39
rect 28 41 32 73
rect 28 39 29 41
rect 31 39 32 41
rect 28 37 32 39
rect 38 72 42 73
rect 38 71 45 72
rect 38 69 41 71
rect 43 69 45 71
rect 38 68 45 69
rect 28 32 32 33
rect 38 32 42 68
rect 28 28 42 32
rect 28 22 32 28
rect 38 27 42 28
rect 48 41 52 63
rect 48 39 49 41
rect 51 39 52 41
rect 48 27 52 39
rect 58 41 62 73
rect 58 39 59 41
rect 61 39 62 41
rect 58 27 62 39
rect 25 21 32 22
rect 25 19 27 21
rect 29 19 32 21
rect 25 18 32 19
rect 37 21 67 22
rect 37 19 39 21
rect 41 19 63 21
rect 65 19 67 21
rect 37 18 67 19
rect 28 17 32 18
rect -2 11 72 12
rect -2 9 5 11
rect 7 9 51 11
rect 53 9 72 11
rect -2 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 72 9
rect -2 0 72 7
<< ptie >>
rect 21 9 43 11
rect 21 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 43 9
rect 21 5 43 7
<< nmos >>
rect 11 16 13 34
rect 21 17 23 34
rect 33 17 35 34
rect 45 17 47 34
rect 57 16 59 34
<< pmos >>
rect 11 55 13 84
rect 23 56 25 85
rect 35 56 37 94
rect 47 55 49 94
rect 57 55 59 94
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 49 39 51 41
rect 59 39 61 41
<< ndifct1 >>
rect 27 19 29 21
rect 39 19 41 21
rect 63 19 65 21
rect 5 9 7 11
rect 51 9 53 11
<< ptiect1 >>
rect 23 7 25 9
rect 31 7 33 9
rect 39 7 41 9
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 29 79 31 81
rect 41 69 43 71
rect 63 79 65 81
<< labels >>
rlabel alu1 10 45 10 45 6 i0
rlabel alu1 30 25 30 25 6 nq
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 30 55 30 55 6 i4
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 40 50 40 50 6 nq
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 50 60 50 6 i3
<< end >>
