magic
tech scmos
timestamp 1199202561
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 56 11 60
rect 19 58 21 63
rect 29 58 31 63
rect 39 60 41 64
rect 49 60 51 65
rect 9 34 11 40
rect 19 35 21 40
rect 29 35 31 40
rect 9 32 15 34
rect 9 30 11 32
rect 13 30 15 32
rect 9 28 15 30
rect 19 33 31 35
rect 19 31 27 33
rect 29 31 31 33
rect 19 29 31 31
rect 12 25 14 28
rect 19 25 21 29
rect 29 18 31 29
rect 39 27 41 40
rect 49 35 51 38
rect 45 33 51 35
rect 45 31 47 33
rect 49 31 51 33
rect 45 29 51 31
rect 35 25 41 27
rect 49 26 51 29
rect 35 23 37 25
rect 39 23 41 25
rect 35 21 41 23
rect 36 18 38 21
rect 49 11 51 15
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 7
rect 36 2 38 7
<< ndif >>
rect 4 10 12 25
rect 4 8 7 10
rect 9 8 12 10
rect 4 6 12 8
rect 14 6 19 25
rect 21 18 26 25
rect 43 18 49 26
rect 21 16 29 18
rect 21 14 24 16
rect 26 14 29 16
rect 21 7 29 14
rect 31 7 36 18
rect 38 15 49 18
rect 51 24 58 26
rect 51 22 54 24
rect 56 22 58 24
rect 51 20 58 22
rect 51 15 56 20
rect 38 13 43 15
rect 45 13 47 15
rect 38 7 47 13
rect 21 6 26 7
<< pdif >>
rect 34 58 39 60
rect 14 56 19 58
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 40 9 52
rect 11 49 19 56
rect 11 47 14 49
rect 16 47 19 49
rect 11 40 19 47
rect 21 56 29 58
rect 21 54 24 56
rect 26 54 29 56
rect 21 40 29 54
rect 31 56 39 58
rect 31 54 34 56
rect 36 54 39 56
rect 31 49 39 54
rect 31 47 34 49
rect 36 47 39 49
rect 31 40 39 47
rect 41 56 49 60
rect 41 54 44 56
rect 46 54 49 56
rect 41 49 49 54
rect 41 47 44 49
rect 46 47 49 49
rect 41 40 49 47
rect 43 38 49 40
rect 51 51 56 60
rect 51 49 58 51
rect 51 47 54 49
rect 56 47 58 49
rect 51 42 58 47
rect 51 40 54 42
rect 56 40 58 42
rect 51 38 58 40
<< alu1 >>
rect -2 67 66 72
rect -2 65 7 67
rect 9 65 66 67
rect -2 64 66 65
rect 33 56 38 59
rect 33 54 34 56
rect 36 54 38 56
rect 33 50 38 54
rect 12 49 38 50
rect 12 47 14 49
rect 16 47 34 49
rect 36 47 38 49
rect 12 46 38 47
rect 2 18 6 43
rect 17 38 30 42
rect 26 33 30 38
rect 41 35 47 42
rect 26 31 27 33
rect 29 31 30 33
rect 26 29 30 31
rect 34 33 50 35
rect 34 31 47 33
rect 49 31 50 33
rect 34 29 50 31
rect 2 16 28 18
rect 2 14 24 16
rect 26 14 28 16
rect 22 13 28 14
rect -2 7 66 8
rect -2 5 53 7
rect 55 5 66 7
rect -2 0 66 5
<< ptie >>
rect 51 7 57 9
rect 51 5 53 7
rect 55 5 57 7
rect 51 3 57 5
<< ntie >>
rect 3 67 13 69
rect 3 65 7 67
rect 9 65 13 67
rect 3 63 13 65
<< nmos >>
rect 12 6 14 25
rect 19 6 21 25
rect 29 7 31 18
rect 36 7 38 18
rect 49 15 51 26
<< pmos >>
rect 9 40 11 56
rect 19 40 21 58
rect 29 40 31 58
rect 39 40 41 60
rect 49 38 51 60
<< polyct0 >>
rect 11 30 13 32
rect 37 23 39 25
<< polyct1 >>
rect 27 31 29 33
rect 47 31 49 33
<< ndifct0 >>
rect 7 8 9 10
rect 54 22 56 24
rect 43 13 45 15
<< ndifct1 >>
rect 24 14 26 16
<< ntiect1 >>
rect 7 65 9 67
<< ptiect1 >>
rect 53 5 55 7
<< pdifct0 >>
rect 4 52 6 54
rect 24 54 26 56
rect 44 54 46 56
rect 44 47 46 49
rect 54 47 56 49
rect 54 40 56 42
<< pdifct1 >>
rect 14 47 16 49
rect 34 54 36 56
rect 34 47 36 49
<< alu0 >>
rect 3 54 7 64
rect 3 52 4 54
rect 6 52 7 54
rect 22 56 28 64
rect 22 54 24 56
rect 26 54 28 56
rect 22 53 28 54
rect 3 50 7 52
rect 10 46 12 50
rect 42 56 48 64
rect 42 54 44 56
rect 46 54 48 56
rect 42 49 48 54
rect 42 47 44 49
rect 46 47 48 49
rect 42 46 48 47
rect 53 49 57 51
rect 53 47 54 49
rect 56 47 57 49
rect 10 43 14 46
rect 6 39 14 43
rect 53 42 57 47
rect 10 32 14 34
rect 10 30 11 32
rect 13 30 14 32
rect 10 26 14 30
rect 53 40 54 42
rect 56 40 57 42
rect 53 26 57 40
rect 10 25 57 26
rect 10 23 37 25
rect 39 24 57 25
rect 39 23 54 24
rect 10 22 54 23
rect 56 22 57 24
rect 53 20 57 22
rect 42 15 46 17
rect 42 13 43 15
rect 45 13 46 15
rect 5 10 11 11
rect 5 8 7 10
rect 9 8 11 10
rect 42 8 46 13
<< labels >>
rlabel alu0 12 28 12 28 6 an
rlabel alu0 33 24 33 24 6 an
rlabel alu0 55 35 55 35 6 an
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 16 20 16 6 z
rlabel polyct1 28 32 28 32 6 b
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 32 36 32 6 a
rlabel alu1 44 36 44 36 6 a
rlabel alu1 36 56 36 56 6 z
rlabel alu1 32 68 32 68 6 vdd
<< end >>
