magic
tech scmos
timestamp 1199202062
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 54 11 59
rect 21 61 27 63
rect 21 59 23 61
rect 25 59 27 61
rect 21 57 27 59
rect 21 54 23 57
rect 9 39 11 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 30 11 33
rect 21 30 23 42
rect 9 19 11 24
rect 21 19 23 24
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 11 28 21 30
rect 11 26 15 28
rect 17 26 21 28
rect 11 24 21 26
rect 23 28 30 30
rect 23 26 26 28
rect 28 26 30 28
rect 23 24 30 26
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 54 19 69
rect 4 48 9 54
rect 2 46 9 48
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 42 21 54
rect 23 48 28 54
rect 23 46 30 48
rect 23 44 26 46
rect 28 44 30 46
rect 23 42 30 44
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 71 34 79
rect -2 69 15 71
rect 17 69 34 71
rect -2 68 34 69
rect 18 61 30 63
rect 18 59 23 61
rect 25 59 30 61
rect 18 57 30 59
rect 2 49 14 55
rect 18 49 22 57
rect 2 46 6 49
rect 2 44 4 46
rect 2 29 6 44
rect 2 28 8 29
rect 2 26 4 28
rect 6 26 8 28
rect 2 25 8 26
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 24 11 30
rect 21 24 23 30
<< pmos >>
rect 9 42 11 54
rect 21 42 23 54
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 23 59 25 61
<< ndifct0 >>
rect 15 26 17 28
rect 26 26 28 28
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 26 44 28 46
<< pdifct1 >>
rect 15 69 17 71
rect 4 44 6 46
<< alu0 >>
rect 6 42 7 49
rect 25 46 29 48
rect 25 44 26 46
rect 28 44 29 46
rect 25 38 29 44
rect 9 37 29 38
rect 9 35 11 37
rect 13 35 29 37
rect 9 34 29 35
rect 14 28 18 30
rect 14 26 15 28
rect 17 26 18 28
rect 14 12 18 26
rect 25 28 29 34
rect 25 26 26 28
rect 28 26 29 28
rect 25 24 29 26
<< labels >>
rlabel alu0 27 36 27 36 6 an
rlabel alu0 19 36 19 36 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 20 56 20 56 6 a
rlabel alu1 28 60 28 60 6 a
<< end >>
