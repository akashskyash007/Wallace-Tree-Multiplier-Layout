magic
tech scmos
timestamp 1199201834
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 29 68 31 73
rect 9 58 11 63
rect 19 58 21 63
rect 45 54 47 58
rect 29 47 31 52
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 9 39 11 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 12 22 14 33
rect 19 31 21 42
rect 29 41 35 43
rect 19 29 25 31
rect 19 27 21 29
rect 23 27 25 29
rect 19 25 25 27
rect 22 22 24 25
rect 29 22 31 41
rect 45 39 47 42
rect 45 37 54 39
rect 45 35 50 37
rect 52 35 54 37
rect 41 33 54 35
rect 41 25 43 33
rect 12 11 14 16
rect 22 10 24 15
rect 29 10 31 15
rect 41 14 43 19
<< ndif >>
rect 33 22 41 25
rect 2 20 12 22
rect 2 18 4 20
rect 6 18 12 20
rect 2 16 12 18
rect 14 20 22 22
rect 14 18 17 20
rect 19 18 22 20
rect 14 16 22 18
rect 17 15 22 16
rect 24 15 29 22
rect 31 20 41 22
rect 31 18 35 20
rect 37 19 41 20
rect 43 23 50 25
rect 43 21 46 23
rect 48 21 50 23
rect 43 19 50 21
rect 37 18 39 19
rect 31 15 39 18
<< pdif >>
rect 21 71 27 73
rect 21 69 23 71
rect 25 69 27 71
rect 21 68 27 69
rect 21 65 29 68
rect 23 58 29 65
rect 4 55 9 58
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 56 19 58
rect 11 54 14 56
rect 16 54 19 56
rect 11 42 19 54
rect 21 52 29 58
rect 31 64 36 68
rect 48 64 54 66
rect 31 62 38 64
rect 31 60 34 62
rect 36 60 38 62
rect 48 62 50 64
rect 52 62 54 64
rect 48 60 54 62
rect 31 58 38 60
rect 31 52 36 58
rect 49 54 54 60
rect 21 42 27 52
rect 40 48 45 54
rect 38 46 45 48
rect 38 44 40 46
rect 42 44 45 46
rect 38 42 45 44
rect 47 42 54 54
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 23 71
rect 25 69 58 71
rect -2 68 58 69
rect 49 64 53 68
rect 49 62 50 64
rect 52 62 53 64
rect 49 60 53 62
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 26 46 30 55
rect 41 50 54 55
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 17 45 35 46
rect 17 43 31 45
rect 33 43 35 45
rect 17 42 35 43
rect 2 31 6 42
rect 50 39 54 50
rect 2 25 14 31
rect 18 29 38 31
rect 18 27 21 29
rect 23 27 38 29
rect 18 25 38 27
rect 10 21 14 25
rect 10 20 21 21
rect 10 18 17 20
rect 19 18 21 20
rect 10 17 21 18
rect 26 17 30 25
rect 49 37 54 39
rect 49 35 50 37
rect 52 35 54 37
rect 49 33 54 35
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 12 16 14 22
rect 22 15 24 22
rect 29 15 31 22
rect 41 19 43 25
<< pmos >>
rect 9 42 11 58
rect 19 42 21 58
rect 29 52 31 68
rect 45 42 47 54
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 21 27 23 29
rect 50 35 52 37
<< ndifct0 >>
rect 4 18 6 20
rect 35 18 37 20
rect 46 21 48 23
<< ndifct1 >>
rect 17 18 19 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 14 54 16 56
rect 34 60 36 62
rect 40 44 42 46
<< pdifct1 >>
rect 23 69 25 71
rect 4 51 6 53
rect 4 44 6 46
rect 50 62 52 64
<< alu0 >>
rect 13 62 38 63
rect 13 60 34 62
rect 36 60 38 62
rect 13 59 38 60
rect 13 56 17 59
rect 13 54 14 56
rect 16 54 17 56
rect 13 52 17 54
rect 38 46 44 47
rect 38 44 40 46
rect 42 44 44 46
rect 38 38 44 44
rect 9 37 46 38
rect 9 35 11 37
rect 13 35 46 37
rect 9 34 46 35
rect 3 20 7 22
rect 3 18 4 20
rect 6 18 7 20
rect 3 12 7 18
rect 42 24 46 34
rect 42 23 50 24
rect 34 20 38 22
rect 42 21 46 23
rect 48 21 50 23
rect 42 20 50 21
rect 34 18 35 20
rect 37 18 38 20
rect 34 12 38 18
<< labels >>
rlabel alu0 15 57 15 57 6 n1
rlabel alu0 25 61 25 61 6 n1
rlabel alu0 44 29 44 29 6 bn
rlabel alu0 27 36 27 36 6 bn
rlabel alu0 41 40 41 40 6 bn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 20 28 20 28 6 a2
rlabel alu1 20 44 20 44 6 a1
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 24 28 24 6 a2
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 28 48 28 48 6 a1
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 52 44 52 44 6 b
rlabel alu1 44 52 44 52 6 b
<< end >>
