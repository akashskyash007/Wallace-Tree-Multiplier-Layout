magic
tech scmos
timestamp 1199203142
<< ab >>
rect 0 0 192 80
<< nwell >>
rect -5 36 197 88
<< pwell >>
rect -5 -8 197 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 56 70 58 74
rect 66 70 68 74
rect 73 70 75 74
rect 83 70 85 74
rect 90 70 92 74
rect 100 70 102 74
rect 107 70 109 74
rect 117 70 119 74
rect 124 70 126 74
rect 134 70 136 74
rect 141 70 143 74
rect 151 70 153 74
rect 158 70 160 74
rect 168 63 170 68
rect 175 63 177 68
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 9 37 41 39
rect 9 35 27 37
rect 29 35 31 37
rect 9 33 31 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 37
rect 45 37 51 39
rect 56 39 58 42
rect 66 39 68 42
rect 56 37 68 39
rect 73 39 75 42
rect 83 39 85 42
rect 73 37 85 39
rect 90 39 92 42
rect 100 39 102 42
rect 90 37 102 39
rect 107 39 109 42
rect 117 39 119 42
rect 124 39 126 42
rect 134 39 136 42
rect 107 37 119 39
rect 123 37 136 39
rect 141 39 143 42
rect 151 39 153 42
rect 141 37 153 39
rect 158 39 160 42
rect 168 39 170 42
rect 158 37 170 39
rect 175 39 177 42
rect 175 37 183 39
rect 45 35 47 37
rect 49 35 51 37
rect 45 33 51 35
rect 59 29 61 37
rect 76 35 78 37
rect 80 35 82 37
rect 76 33 82 35
rect 70 29 72 33
rect 80 29 82 33
rect 90 35 92 37
rect 94 35 96 37
rect 90 33 96 35
rect 107 35 112 37
rect 114 35 116 37
rect 107 33 116 35
rect 123 35 129 37
rect 123 33 125 35
rect 127 33 129 35
rect 141 35 143 37
rect 145 35 147 37
rect 141 33 147 35
rect 158 35 162 37
rect 164 35 168 37
rect 158 33 168 35
rect 175 35 179 37
rect 181 35 183 37
rect 175 33 183 35
rect 49 25 51 29
rect 90 28 92 33
rect 100 31 116 33
rect 122 31 129 33
rect 134 31 147 33
rect 156 31 168 33
rect 100 28 102 31
rect 112 28 114 31
rect 122 28 124 31
rect 134 28 136 31
rect 144 28 146 31
rect 156 28 158 31
rect 166 28 168 31
rect 177 30 179 33
rect 80 12 82 16
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
rect 39 8 41 11
rect 49 8 51 11
rect 39 6 51 8
rect 59 8 61 11
rect 70 8 72 11
rect 90 8 92 16
rect 59 6 92 8
rect 100 6 102 10
rect 112 6 114 10
rect 122 6 124 10
rect 177 15 179 19
rect 134 6 136 10
rect 144 6 146 10
rect 156 8 158 13
rect 166 8 168 13
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 10 19 26
rect 21 20 29 30
rect 21 18 24 20
rect 26 18 29 20
rect 21 10 29 18
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 11 39 26
rect 41 25 46 30
rect 54 25 59 29
rect 41 20 49 25
rect 41 18 44 20
rect 46 18 49 20
rect 41 11 49 18
rect 51 23 59 25
rect 51 21 54 23
rect 56 21 59 23
rect 51 11 59 21
rect 61 15 70 29
rect 61 13 65 15
rect 67 13 70 15
rect 61 11 70 13
rect 72 25 80 29
rect 72 23 75 25
rect 77 23 80 25
rect 72 16 80 23
rect 82 28 87 29
rect 170 28 177 30
rect 82 20 90 28
rect 82 18 85 20
rect 87 18 90 20
rect 82 16 90 18
rect 92 25 100 28
rect 92 23 95 25
rect 97 23 100 25
rect 92 16 100 23
rect 72 11 77 16
rect 31 10 36 11
rect 95 10 100 16
rect 102 11 112 28
rect 102 10 106 11
rect 104 9 106 10
rect 108 10 112 11
rect 114 20 122 28
rect 114 18 117 20
rect 119 18 122 20
rect 114 10 122 18
rect 124 11 134 28
rect 124 10 128 11
rect 108 9 110 10
rect 104 7 110 9
rect 126 9 128 10
rect 130 10 134 11
rect 136 20 144 28
rect 136 18 139 20
rect 141 18 144 20
rect 136 10 144 18
rect 146 13 156 28
rect 158 20 166 28
rect 158 18 161 20
rect 163 18 166 20
rect 158 13 166 18
rect 168 19 177 28
rect 179 28 186 30
rect 179 26 182 28
rect 184 26 186 28
rect 179 24 186 26
rect 179 19 184 24
rect 168 17 175 19
rect 168 15 171 17
rect 173 15 175 17
rect 168 13 175 15
rect 146 11 154 13
rect 146 10 150 11
rect 130 9 132 10
rect 126 7 132 9
rect 148 9 150 10
rect 152 9 154 11
rect 148 7 154 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 61 49 66
rect 41 59 44 61
rect 46 59 49 61
rect 41 42 49 59
rect 51 42 56 70
rect 58 61 66 70
rect 58 59 61 61
rect 63 59 66 61
rect 58 53 66 59
rect 58 51 61 53
rect 63 51 66 53
rect 58 42 66 51
rect 68 42 73 70
rect 75 68 83 70
rect 75 66 78 68
rect 80 66 83 68
rect 75 61 83 66
rect 75 59 78 61
rect 80 59 83 61
rect 75 42 83 59
rect 85 42 90 70
rect 92 60 100 70
rect 92 58 95 60
rect 97 58 100 60
rect 92 53 100 58
rect 92 51 95 53
rect 97 51 100 53
rect 92 42 100 51
rect 102 42 107 70
rect 109 68 117 70
rect 109 66 112 68
rect 114 66 117 68
rect 109 61 117 66
rect 109 59 112 61
rect 114 59 117 61
rect 109 42 117 59
rect 119 42 124 70
rect 126 61 134 70
rect 126 59 129 61
rect 131 59 134 61
rect 126 53 134 59
rect 126 51 129 53
rect 131 51 134 53
rect 126 42 134 51
rect 136 42 141 70
rect 143 68 151 70
rect 143 66 146 68
rect 148 66 151 68
rect 143 61 151 66
rect 143 59 146 61
rect 148 59 151 61
rect 143 42 151 59
rect 153 42 158 70
rect 160 63 165 70
rect 160 61 168 63
rect 160 59 163 61
rect 165 59 168 61
rect 160 54 168 59
rect 160 52 163 54
rect 165 52 168 54
rect 160 42 168 52
rect 170 42 175 63
rect 177 61 185 63
rect 177 59 180 61
rect 182 59 185 61
rect 177 54 185 59
rect 177 52 180 54
rect 182 52 185 54
rect 177 42 185 52
<< alu1 >>
rect -2 81 194 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 194 81
rect -2 68 194 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 58 61 64 63
rect 58 59 61 61
rect 63 59 64 61
rect 58 54 64 59
rect 128 61 134 63
rect 128 59 129 61
rect 131 59 134 61
rect 128 54 134 59
rect 162 61 166 63
rect 162 59 163 61
rect 165 59 166 61
rect 162 54 166 59
rect 12 53 163 54
rect 12 51 14 53
rect 16 51 34 53
rect 36 51 61 53
rect 63 51 95 53
rect 97 51 129 53
rect 131 52 163 53
rect 165 52 166 54
rect 131 51 166 52
rect 12 50 166 51
rect 12 47 17 50
rect 2 46 17 47
rect 170 46 174 55
rect 2 44 14 46
rect 16 44 17 46
rect 2 42 17 44
rect 25 42 39 46
rect 78 42 183 46
rect 2 28 6 42
rect 2 26 4 28
rect 2 21 6 26
rect 25 38 31 42
rect 78 38 82 42
rect 17 37 31 38
rect 17 35 27 37
rect 29 35 31 37
rect 17 34 31 35
rect 41 37 82 38
rect 41 35 47 37
rect 49 35 78 37
rect 80 35 82 37
rect 41 34 82 35
rect 89 37 106 38
rect 89 35 92 37
rect 94 35 106 37
rect 89 34 106 35
rect 102 30 106 34
rect 153 37 167 38
rect 153 35 162 37
rect 164 35 167 37
rect 153 34 167 35
rect 177 37 183 42
rect 177 35 179 37
rect 181 35 183 37
rect 177 34 183 35
rect 153 30 159 34
rect 102 26 159 30
rect 2 19 4 21
rect 6 20 48 21
rect 6 19 24 20
rect 2 18 24 19
rect 26 18 44 20
rect 46 18 48 20
rect 2 17 48 18
rect -2 11 194 12
rect -2 9 106 11
rect 108 9 128 11
rect 130 9 150 11
rect 152 9 194 11
rect -2 1 194 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 194 1
rect -2 -2 194 -1
<< ptie >>
rect 0 1 192 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 192 1
rect 0 -3 192 -1
<< ntie >>
rect 0 81 192 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 192 81
rect 0 77 192 79
<< nmos >>
rect 9 10 11 30
rect 19 10 21 30
rect 29 10 31 30
rect 39 11 41 30
rect 49 11 51 25
rect 59 11 61 29
rect 70 11 72 29
rect 80 16 82 29
rect 90 16 92 28
rect 100 10 102 28
rect 112 10 114 28
rect 122 10 124 28
rect 134 10 136 28
rect 144 10 146 28
rect 156 13 158 28
rect 166 13 168 28
rect 177 19 179 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 56 42 58 70
rect 66 42 68 70
rect 73 42 75 70
rect 83 42 85 70
rect 90 42 92 70
rect 100 42 102 70
rect 107 42 109 70
rect 117 42 119 70
rect 124 42 126 70
rect 134 42 136 70
rect 141 42 143 70
rect 151 42 153 70
rect 158 42 160 70
rect 168 42 170 63
rect 175 42 177 63
<< polyct0 >>
rect 112 35 114 37
rect 125 33 127 35
rect 143 35 145 37
<< polyct1 >>
rect 27 35 29 37
rect 47 35 49 37
rect 78 35 80 37
rect 92 35 94 37
rect 162 35 164 37
rect 179 35 181 37
<< ndifct0 >>
rect 14 26 16 28
rect 34 26 36 28
rect 54 21 56 23
rect 65 13 67 15
rect 75 23 77 25
rect 85 18 87 20
rect 95 23 97 25
rect 117 18 119 20
rect 139 18 141 20
rect 161 18 163 20
rect 182 26 184 28
rect 171 15 173 17
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
rect 24 18 26 20
rect 44 18 46 20
rect 106 9 108 11
rect 128 9 130 11
rect 150 9 152 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
rect 171 79 173 81
rect 179 79 181 81
rect 187 79 189 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
rect 171 -1 173 1
rect 179 -1 181 1
rect 187 -1 189 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 66 26 68
rect 24 59 26 61
rect 44 66 46 68
rect 44 59 46 61
rect 78 66 80 68
rect 78 59 80 61
rect 95 58 97 60
rect 112 66 114 68
rect 112 59 114 61
rect 146 66 148 68
rect 146 59 148 61
rect 180 59 182 61
rect 180 52 182 54
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
rect 34 59 36 61
rect 34 51 36 53
rect 61 59 63 61
rect 61 51 63 53
rect 95 51 97 53
rect 129 59 131 61
rect 129 51 131 53
rect 163 59 165 61
rect 163 52 165 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 42 66 44 68
rect 46 66 48 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 42 61 48 66
rect 76 66 78 68
rect 80 66 82 68
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 76 61 82 66
rect 110 66 112 68
rect 114 66 116 68
rect 76 59 78 61
rect 80 59 82 61
rect 76 58 82 59
rect 94 60 98 62
rect 94 58 95 60
rect 97 58 98 60
rect 110 61 116 66
rect 144 66 146 68
rect 148 66 150 68
rect 110 59 112 61
rect 114 59 116 61
rect 110 58 116 59
rect 94 54 98 58
rect 144 61 150 66
rect 144 59 146 61
rect 148 59 150 61
rect 144 58 150 59
rect 179 61 183 68
rect 179 59 180 61
rect 182 59 183 61
rect 179 54 183 59
rect 179 52 180 54
rect 182 52 183 54
rect 179 50 183 52
rect 6 21 7 42
rect 110 37 116 42
rect 141 37 147 42
rect 110 35 112 37
rect 114 35 116 37
rect 110 34 116 35
rect 124 35 128 37
rect 124 33 125 35
rect 127 33 128 35
rect 141 35 143 37
rect 145 35 147 37
rect 141 34 147 35
rect 124 30 128 33
rect 12 28 98 29
rect 12 26 14 28
rect 16 26 34 28
rect 36 26 98 28
rect 162 28 186 29
rect 162 26 182 28
rect 184 26 186 28
rect 12 25 98 26
rect 53 23 57 25
rect 53 21 54 23
rect 56 21 57 23
rect 74 23 75 25
rect 77 23 78 25
rect 74 21 78 23
rect 94 23 95 25
rect 97 23 98 25
rect 94 21 98 23
rect 162 25 186 26
rect 162 21 166 25
rect 53 19 57 21
rect 83 20 89 21
rect 83 18 85 20
rect 87 18 89 20
rect 64 15 68 17
rect 64 13 65 15
rect 67 13 68 15
rect 64 12 68 13
rect 83 12 89 18
rect 94 20 166 21
rect 94 18 117 20
rect 119 18 139 20
rect 141 18 161 20
rect 163 18 166 20
rect 94 17 166 18
rect 170 17 174 19
rect 170 15 171 17
rect 173 15 174 17
rect 170 12 174 15
<< labels >>
rlabel alu0 55 24 55 24 6 n1
rlabel alu0 55 27 55 27 6 n1
rlabel alu0 96 23 96 23 6 n1
rlabel alu0 130 19 130 19 6 n1
rlabel alu0 174 27 174 27 6 n1
rlabel alu1 4 32 4 32 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 36 20 36 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 44 36 44 6 b
rlabel alu1 68 36 68 36 6 a1
rlabel alu1 60 36 60 36 6 a1
rlabel alu1 52 36 52 36 6 a1
rlabel alu1 44 36 44 36 6 a1
rlabel alu1 44 52 44 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 60 56 60 56 6 z
rlabel alu1 96 6 96 6 6 vss
rlabel alu1 108 28 108 28 6 a2
rlabel alu1 76 36 76 36 6 a1
rlabel alu1 100 44 100 44 6 a1
rlabel alu1 108 44 108 44 6 a1
rlabel alu1 100 36 100 36 6 a2
rlabel alu1 84 44 84 44 6 a1
rlabel alu1 92 44 92 44 6 a1
rlabel alu1 92 36 92 36 6 a2
rlabel alu1 84 52 84 52 6 z
rlabel alu1 92 52 92 52 6 z
rlabel alu1 100 52 100 52 6 z
rlabel alu1 108 52 108 52 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 96 74 96 74 6 vdd
rlabel alu1 116 28 116 28 6 a2
rlabel alu1 132 28 132 28 6 a2
rlabel alu1 140 28 140 28 6 a2
rlabel alu1 148 28 148 28 6 a2
rlabel alu1 124 28 124 28 6 a2
rlabel alu1 116 44 116 44 6 a1
rlabel alu1 132 44 132 44 6 a1
rlabel alu1 140 44 140 44 6 a1
rlabel alu1 148 44 148 44 6 a1
rlabel alu1 124 44 124 44 6 a1
rlabel alu1 124 52 124 52 6 z
rlabel alu1 140 52 140 52 6 z
rlabel alu1 148 52 148 52 6 z
rlabel alu1 116 52 116 52 6 z
rlabel alu1 132 56 132 56 6 z
rlabel alu1 156 32 156 32 6 a2
rlabel alu1 156 44 156 44 6 a1
rlabel alu1 164 44 164 44 6 a1
rlabel alu1 180 40 180 40 6 a1
rlabel alu1 164 36 164 36 6 a2
rlabel alu1 172 48 172 48 6 a1
rlabel alu1 156 52 156 52 6 z
rlabel pdifct1 164 60 164 60 6 z
<< end >>
