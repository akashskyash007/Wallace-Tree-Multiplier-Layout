magic
tech scmos
timestamp 1199470679
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 13 94 15 98
rect 21 94 23 98
rect 33 94 35 98
rect 45 94 47 98
rect 57 94 59 98
rect 13 48 15 57
rect 21 54 23 57
rect 33 54 35 57
rect 21 52 27 54
rect 33 52 41 54
rect 25 48 27 52
rect 35 50 41 52
rect 35 48 37 50
rect 39 48 41 50
rect 13 46 21 48
rect 13 45 17 46
rect 11 44 17 45
rect 19 44 21 46
rect 11 42 21 44
rect 25 46 31 48
rect 35 46 41 48
rect 25 44 27 46
rect 29 44 31 46
rect 25 42 31 44
rect 45 42 47 57
rect 57 53 59 57
rect 51 51 59 53
rect 51 49 53 51
rect 55 49 59 51
rect 51 47 59 49
rect 11 33 13 42
rect 25 38 27 42
rect 45 40 53 42
rect 45 38 49 40
rect 51 38 53 40
rect 23 36 27 38
rect 35 36 53 38
rect 23 33 25 36
rect 35 33 37 36
rect 57 33 59 47
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 57 12 59 17
<< ndif >>
rect 6 23 11 33
rect 3 21 11 23
rect 3 19 5 21
rect 7 19 11 21
rect 3 17 11 19
rect 13 29 23 33
rect 13 27 17 29
rect 19 27 23 29
rect 13 17 23 27
rect 25 31 35 33
rect 25 29 29 31
rect 31 29 35 31
rect 25 17 35 29
rect 37 17 57 33
rect 59 31 67 33
rect 59 29 63 31
rect 65 29 67 31
rect 59 23 67 29
rect 59 21 63 23
rect 65 21 67 23
rect 59 19 67 21
rect 59 17 64 19
rect 39 11 55 17
rect 39 9 41 11
rect 43 9 51 11
rect 53 9 55 11
rect 39 7 55 9
<< pdif >>
rect 4 91 13 94
rect 4 89 7 91
rect 9 89 13 91
rect 4 57 13 89
rect 15 57 21 94
rect 23 81 33 94
rect 23 79 27 81
rect 29 79 33 81
rect 23 57 33 79
rect 35 81 45 94
rect 35 79 39 81
rect 41 79 45 81
rect 35 73 45 79
rect 35 71 39 73
rect 41 71 45 73
rect 35 57 45 71
rect 47 91 57 94
rect 47 89 51 91
rect 53 89 57 91
rect 47 81 57 89
rect 47 79 51 81
rect 53 79 57 81
rect 47 71 57 79
rect 47 69 51 71
rect 53 69 57 71
rect 47 57 57 69
rect 59 71 64 94
rect 59 69 67 71
rect 59 67 63 69
rect 65 67 67 69
rect 59 61 67 67
rect 59 59 63 61
rect 65 59 67 61
rect 59 57 67 59
<< alu1 >>
rect -2 91 72 100
rect -2 89 7 91
rect 9 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 8 81 33 83
rect 8 79 27 81
rect 29 79 33 81
rect 8 78 33 79
rect 38 81 42 83
rect 38 79 39 81
rect 41 79 42 81
rect 8 30 12 78
rect 38 73 42 79
rect 38 72 39 73
rect 18 71 39 72
rect 41 71 42 73
rect 18 68 42 71
rect 50 81 54 88
rect 50 79 51 81
rect 53 79 54 81
rect 50 71 54 79
rect 50 69 51 71
rect 53 69 54 71
rect 18 48 22 68
rect 50 67 54 69
rect 62 69 66 71
rect 62 67 63 69
rect 65 67 66 69
rect 62 62 66 67
rect 16 46 22 48
rect 16 44 17 46
rect 19 44 22 46
rect 16 42 22 44
rect 26 61 66 62
rect 26 59 63 61
rect 65 59 66 61
rect 26 58 66 59
rect 26 46 30 58
rect 26 44 27 46
rect 29 44 30 46
rect 26 42 30 44
rect 36 51 57 52
rect 36 50 53 51
rect 36 48 37 50
rect 39 49 53 50
rect 55 49 57 51
rect 39 48 57 49
rect 18 38 22 42
rect 18 34 32 38
rect 36 37 42 48
rect 47 40 53 42
rect 47 38 49 40
rect 51 38 53 40
rect 28 31 32 34
rect 47 32 53 38
rect 8 29 21 30
rect 8 27 17 29
rect 19 27 21 29
rect 28 29 29 31
rect 31 29 32 31
rect 28 27 32 29
rect 37 28 53 32
rect 62 31 66 58
rect 62 29 63 31
rect 65 29 66 31
rect 8 26 21 27
rect 62 23 66 29
rect 62 22 63 23
rect 3 21 63 22
rect 65 21 66 23
rect 3 19 5 21
rect 7 19 66 21
rect 3 18 66 19
rect -2 11 72 12
rect -2 9 41 11
rect 43 9 51 11
rect 53 9 72 11
rect -2 7 72 9
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 72 7
rect -2 0 72 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< nmos >>
rect 11 17 13 33
rect 23 17 25 33
rect 35 17 37 33
rect 57 17 59 33
<< pmos >>
rect 13 57 15 94
rect 21 57 23 94
rect 33 57 35 94
rect 45 57 47 94
rect 57 57 59 94
<< polyct1 >>
rect 37 48 39 50
rect 17 44 19 46
rect 27 44 29 46
rect 53 49 55 51
rect 49 38 51 40
<< ndifct1 >>
rect 5 19 7 21
rect 17 27 19 29
rect 29 29 31 31
rect 63 29 65 31
rect 63 21 65 23
rect 41 9 43 11
rect 51 9 53 11
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 7 89 9 91
rect 27 79 29 81
rect 39 79 41 81
rect 39 71 41 73
rect 51 89 53 91
rect 51 79 53 81
rect 51 69 53 71
rect 63 67 65 69
rect 63 59 65 61
<< labels >>
rlabel alu1 10 55 10 55 6 z
rlabel alu1 30 32 30 32 6 an
rlabel alu1 28 52 28 52 6 bn
rlabel alu1 20 53 20 53 6 an
rlabel alu1 20 80 20 80 6 z
rlabel alu1 30 80 30 80 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 45 40 45 6 b
rlabel alu1 40 30 40 30 6 a
rlabel alu1 50 35 50 35 6 a
rlabel alu1 50 50 50 50 6 b
rlabel alu1 40 75 40 75 6 an
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 34 20 34 20 6 bn
rlabel alu1 64 44 64 44 6 bn
rlabel alu1 46 60 46 60 6 bn
<< end >>
