magic
tech scmos
timestamp 1199469020
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -2 48 52 104
<< pwell >>
rect -2 -4 52 48
<< poly >>
rect 13 94 15 98
rect 25 94 27 98
rect 37 94 39 98
rect 13 52 15 55
rect 25 52 27 55
rect 13 50 21 52
rect 13 48 17 50
rect 19 48 21 50
rect 13 46 21 48
rect 25 50 33 52
rect 25 48 29 50
rect 31 48 33 50
rect 25 46 33 48
rect 13 27 15 46
rect 25 34 27 46
rect 37 43 39 55
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 33 37 43 39
rect 33 34 35 37
rect 13 12 15 17
rect 25 12 27 17
rect 33 12 35 17
<< ndif >>
rect 20 27 25 34
rect 4 21 13 27
rect 4 19 7 21
rect 9 19 13 21
rect 4 17 13 19
rect 15 21 25 27
rect 15 19 19 21
rect 21 19 25 21
rect 15 17 25 19
rect 27 17 33 34
rect 35 21 44 34
rect 35 19 39 21
rect 41 19 44 21
rect 35 17 44 19
<< pdif >>
rect 8 69 13 94
rect 5 67 13 69
rect 5 65 7 67
rect 9 65 13 67
rect 5 59 13 65
rect 5 57 7 59
rect 9 57 13 59
rect 5 55 13 57
rect 15 81 25 94
rect 15 79 19 81
rect 21 79 25 81
rect 15 73 25 79
rect 15 71 19 73
rect 21 71 25 73
rect 15 55 25 71
rect 27 91 37 94
rect 27 89 31 91
rect 33 89 37 91
rect 27 81 37 89
rect 27 79 31 81
rect 33 79 37 81
rect 27 55 37 79
rect 39 83 44 94
rect 39 81 47 83
rect 39 79 43 81
rect 45 79 47 81
rect 39 73 47 79
rect 39 71 43 73
rect 45 71 47 73
rect 39 69 47 71
rect 39 55 44 69
<< alu1 >>
rect -2 91 52 100
rect -2 89 31 91
rect 33 89 52 91
rect -2 88 52 89
rect 18 81 22 83
rect 18 79 19 81
rect 21 79 22 81
rect 18 73 22 79
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 77 34 79
rect 42 81 46 83
rect 42 79 43 81
rect 45 79 46 81
rect 6 67 12 73
rect 18 71 19 73
rect 21 72 22 73
rect 42 73 46 79
rect 42 72 43 73
rect 21 71 43 72
rect 45 71 46 73
rect 18 68 46 71
rect 6 65 7 67
rect 9 65 12 67
rect 6 59 12 65
rect 6 57 7 59
rect 9 57 12 59
rect 6 55 12 57
rect 8 32 12 55
rect 18 58 33 63
rect 18 52 22 58
rect 38 53 42 63
rect 16 50 22 52
rect 16 48 17 50
rect 19 48 22 50
rect 16 46 22 48
rect 18 37 22 46
rect 28 50 42 53
rect 28 48 29 50
rect 31 48 42 50
rect 28 47 42 48
rect 28 37 32 47
rect 38 41 42 43
rect 38 39 39 41
rect 41 39 42 41
rect 38 33 42 39
rect 8 27 23 32
rect 6 21 10 23
rect 6 19 7 21
rect 9 19 10 21
rect 6 12 10 19
rect 17 21 23 27
rect 17 19 19 21
rect 21 19 23 21
rect 17 18 23 19
rect 28 27 42 33
rect 28 17 32 27
rect 38 21 42 23
rect 38 19 39 21
rect 41 19 42 21
rect 38 12 42 19
rect -2 7 52 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 52 7
rect -2 0 52 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< nmos >>
rect 13 17 15 27
rect 25 17 27 34
rect 33 17 35 34
<< pmos >>
rect 13 55 15 94
rect 25 55 27 94
rect 37 55 39 94
<< polyct1 >>
rect 17 48 19 50
rect 29 48 31 50
rect 39 39 41 41
<< ndifct1 >>
rect 7 19 9 21
rect 19 19 21 21
rect 39 19 41 21
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 7 65 9 67
rect 7 57 9 59
rect 19 79 21 81
rect 19 71 21 73
rect 31 89 33 91
rect 31 79 33 81
rect 43 79 45 81
rect 43 71 45 73
<< labels >>
rlabel alu1 20 25 20 25 6 z
rlabel alu1 20 50 20 50 6 b
rlabel alu1 10 50 10 50 6 z
rlabel alu1 20 75 20 75 6 n2
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 25 30 25 6 a1
rlabel alu1 30 45 30 45 6 a2
rlabel alu1 30 60 30 60 6 b
rlabel alu1 25 94 25 94 6 vdd
rlabel alu1 40 35 40 35 6 a1
rlabel alu1 40 55 40 55 6 a2
rlabel alu1 32 70 32 70 6 n2
rlabel alu1 44 75 44 75 6 n2
<< end >>
