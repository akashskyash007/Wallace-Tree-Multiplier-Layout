magic
tech scmos
timestamp 1199203324
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 70 11 74
rect 28 70 30 74
rect 35 70 37 74
rect 42 70 44 74
rect 49 70 51 74
rect 9 39 11 42
rect 28 39 30 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 30 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 24 11 33
rect 20 22 22 33
rect 35 31 37 42
rect 30 29 37 31
rect 30 27 33 29
rect 35 27 37 29
rect 30 25 37 27
rect 42 31 44 42
rect 49 39 51 42
rect 49 37 59 39
rect 52 35 55 37
rect 57 35 59 37
rect 52 33 59 35
rect 42 29 48 31
rect 42 27 44 29
rect 46 27 48 29
rect 42 25 48 27
rect 30 22 32 25
rect 42 22 44 25
rect 52 22 54 33
rect 9 6 11 10
rect 20 9 22 14
rect 30 9 32 14
rect 42 9 44 14
rect 52 9 54 14
<< ndif >>
rect 2 22 9 24
rect 2 20 4 22
rect 6 20 9 22
rect 2 18 9 20
rect 4 10 9 18
rect 11 22 18 24
rect 11 21 20 22
rect 11 19 14 21
rect 16 19 20 21
rect 11 14 20 19
rect 22 20 30 22
rect 22 18 25 20
rect 27 18 30 20
rect 22 14 30 18
rect 32 14 42 22
rect 44 20 52 22
rect 44 18 47 20
rect 49 18 52 20
rect 44 14 52 18
rect 54 14 62 22
rect 11 12 14 14
rect 16 12 18 14
rect 11 10 18 12
rect 34 11 40 14
rect 34 9 36 11
rect 38 9 40 11
rect 56 11 62 14
rect 56 9 58 11
rect 60 9 62 11
rect 34 7 40 9
rect 56 7 62 9
<< pdif >>
rect 13 70 19 72
rect 4 56 9 70
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 69 19 70
rect 11 67 15 69
rect 17 67 19 69
rect 11 59 19 67
rect 11 42 17 59
rect 23 55 28 70
rect 21 53 28 55
rect 21 51 23 53
rect 25 51 28 53
rect 21 49 28 51
rect 23 42 28 49
rect 30 42 35 70
rect 37 42 42 70
rect 44 42 49 70
rect 51 68 59 70
rect 51 66 54 68
rect 56 66 59 68
rect 51 61 59 66
rect 51 59 54 61
rect 56 59 59 61
rect 51 42 59 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 69 66 79
rect -2 68 15 69
rect 17 68 66 69
rect 2 57 14 63
rect 2 54 6 57
rect 2 52 4 54
rect 2 24 6 52
rect 34 46 38 63
rect 19 42 38 46
rect 42 46 46 55
rect 42 42 59 46
rect 19 37 25 42
rect 19 35 21 37
rect 23 35 25 37
rect 19 34 25 35
rect 32 34 47 38
rect 53 37 59 42
rect 53 35 55 37
rect 57 35 59 37
rect 53 34 59 35
rect 2 22 7 24
rect 2 20 4 22
rect 6 20 7 22
rect 2 17 7 20
rect 32 29 38 34
rect 32 27 33 29
rect 35 27 38 29
rect 32 25 38 27
rect 42 29 62 30
rect 42 27 44 29
rect 46 27 62 29
rect 42 26 62 27
rect 58 17 62 26
rect -2 11 66 12
rect -2 9 36 11
rect 38 9 58 11
rect 60 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 10 11 24
rect 20 14 22 22
rect 30 14 32 22
rect 42 14 44 22
rect 52 14 54 22
<< pmos >>
rect 9 42 11 70
rect 28 42 30 70
rect 35 42 37 70
rect 42 42 44 70
rect 49 42 51 70
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 21 35 23 37
rect 33 27 35 29
rect 55 35 57 37
rect 44 27 46 29
<< ndifct0 >>
rect 14 19 16 21
rect 25 18 27 20
rect 47 18 49 20
rect 14 12 16 14
<< ndifct1 >>
rect 4 20 6 22
rect 36 9 38 11
rect 58 9 60 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 15 67 17 68
rect 23 51 25 53
rect 54 66 56 68
rect 54 59 56 61
<< pdifct1 >>
rect 4 52 6 54
rect 15 68 17 69
<< alu0 >>
rect 13 67 15 68
rect 17 67 19 68
rect 13 66 19 67
rect 52 66 54 68
rect 56 66 58 68
rect 6 50 7 57
rect 11 53 27 54
rect 11 51 23 53
rect 25 51 27 53
rect 11 50 27 51
rect 11 39 15 50
rect 52 61 58 66
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
rect 10 37 15 39
rect 10 35 11 37
rect 13 35 15 37
rect 10 33 15 35
rect 11 30 15 33
rect 11 26 27 30
rect 12 21 18 22
rect 12 19 14 21
rect 16 19 18 21
rect 12 14 18 19
rect 23 21 27 26
rect 23 20 51 21
rect 23 18 25 20
rect 27 18 47 20
rect 49 18 51 20
rect 23 17 51 18
rect 12 12 14 14
rect 16 12 18 14
<< labels >>
rlabel alu0 13 40 13 40 6 zn
rlabel alu0 19 52 19 52 6 zn
rlabel alu0 37 19 37 19 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 44 28 44 6 d
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 32 36 32 6 c
rlabel alu1 44 36 44 36 6 c
rlabel alu1 36 56 36 56 6 d
rlabel alu1 44 52 44 52 6 a
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 60 20 60 20 6 b
rlabel alu1 52 28 52 28 6 b
rlabel alu1 52 44 52 44 6 a
<< end >>
