magic
tech scmos
timestamp 1199202100
<< ab >>
rect 0 0 88 72
<< nwell >>
rect -5 32 93 77
<< pwell >>
rect -5 -5 93 32
<< poly >>
rect 9 58 11 63
rect 19 58 21 63
rect 39 59 41 64
rect 46 59 48 64
rect 56 59 58 64
rect 66 59 68 64
rect 76 63 78 68
rect 9 35 11 38
rect 19 35 21 42
rect 39 35 41 43
rect 46 35 48 43
rect 56 35 58 43
rect 66 35 68 43
rect 76 35 78 43
rect 5 33 11 35
rect 5 31 7 33
rect 9 31 11 33
rect 5 29 11 31
rect 17 33 23 35
rect 17 31 19 33
rect 21 31 23 33
rect 17 29 23 31
rect 32 33 42 35
rect 32 31 34 33
rect 36 31 42 33
rect 46 32 49 35
rect 32 29 42 31
rect 9 22 11 29
rect 19 19 21 29
rect 40 26 42 29
rect 47 26 49 32
rect 55 33 61 35
rect 55 31 57 33
rect 59 31 61 33
rect 55 29 61 31
rect 65 33 71 35
rect 65 31 67 33
rect 69 31 71 33
rect 65 29 71 31
rect 76 33 86 35
rect 76 31 82 33
rect 84 31 86 33
rect 76 29 86 31
rect 57 26 59 29
rect 67 26 69 29
rect 77 26 79 29
rect 9 7 11 12
rect 19 7 21 12
rect 40 14 42 19
rect 47 10 49 19
rect 57 14 59 19
rect 67 16 69 19
rect 63 14 69 16
rect 63 10 65 14
rect 47 8 65 10
rect 77 11 79 16
<< ndif >>
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 4 12 9 16
rect 11 19 16 22
rect 32 19 40 26
rect 42 19 47 26
rect 49 24 57 26
rect 49 22 52 24
rect 54 22 57 24
rect 49 19 57 22
rect 59 23 67 26
rect 59 21 62 23
rect 64 21 67 23
rect 59 19 67 21
rect 69 19 77 26
rect 11 16 19 19
rect 11 14 14 16
rect 16 14 19 16
rect 11 12 19 14
rect 21 16 28 19
rect 21 14 24 16
rect 26 14 28 16
rect 21 12 28 14
rect 32 7 38 19
rect 71 16 77 19
rect 79 24 86 26
rect 79 22 82 24
rect 84 22 86 24
rect 79 20 86 22
rect 79 16 84 20
rect 71 12 75 16
rect 69 10 75 12
rect 69 8 71 10
rect 73 8 75 10
rect 32 5 34 7
rect 36 5 38 7
rect 69 6 75 8
rect 32 3 38 5
<< pdif >>
rect 70 59 76 63
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 4 38 9 45
rect 11 56 19 58
rect 11 54 14 56
rect 16 54 19 56
rect 11 42 19 54
rect 21 56 28 58
rect 21 54 24 56
rect 26 54 28 56
rect 21 49 28 54
rect 21 47 24 49
rect 26 47 28 49
rect 21 45 28 47
rect 32 57 39 59
rect 32 55 34 57
rect 36 55 39 57
rect 21 42 26 45
rect 32 43 39 55
rect 41 43 46 59
rect 48 48 56 59
rect 48 46 51 48
rect 53 46 56 48
rect 48 43 56 46
rect 58 57 66 59
rect 58 55 61 57
rect 63 55 66 57
rect 58 43 66 55
rect 68 57 76 59
rect 68 55 71 57
rect 73 55 76 57
rect 68 43 76 55
rect 78 59 83 63
rect 78 57 85 59
rect 78 55 81 57
rect 83 55 85 57
rect 78 50 85 55
rect 78 48 81 50
rect 83 48 85 50
rect 78 46 85 48
rect 78 43 83 46
rect 11 38 17 42
<< alu1 >>
rect -2 67 90 72
rect -2 65 29 67
rect 31 65 90 67
rect -2 64 90 65
rect 50 48 54 51
rect 50 46 51 48
rect 53 46 54 48
rect 50 43 54 46
rect 2 35 6 43
rect 2 33 14 35
rect 2 31 7 33
rect 9 31 14 33
rect 2 29 14 31
rect 42 39 54 43
rect 42 25 46 39
rect 58 35 62 51
rect 50 33 62 35
rect 50 31 57 33
rect 59 31 62 33
rect 50 29 62 31
rect 74 37 86 43
rect 81 33 86 37
rect 81 31 82 33
rect 84 31 86 33
rect 81 29 86 31
rect 42 24 56 25
rect 42 22 52 24
rect 54 22 56 24
rect 42 21 56 22
rect -2 7 90 8
rect -2 5 34 7
rect 36 5 81 7
rect 83 5 90 7
rect -2 0 90 5
<< ptie >>
rect 79 7 85 9
rect 79 5 81 7
rect 83 5 85 7
rect 79 3 85 5
<< ntie >>
rect 27 67 33 69
rect 27 65 29 67
rect 31 65 33 67
rect 27 63 33 65
<< nmos >>
rect 9 12 11 22
rect 40 19 42 26
rect 47 19 49 26
rect 57 19 59 26
rect 67 19 69 26
rect 19 12 21 19
rect 77 16 79 26
<< pmos >>
rect 9 38 11 58
rect 19 42 21 58
rect 39 43 41 59
rect 46 43 48 59
rect 56 43 58 59
rect 66 43 68 59
rect 76 43 78 63
<< polyct0 >>
rect 19 31 21 33
rect 34 31 36 33
rect 67 31 69 33
<< polyct1 >>
rect 7 31 9 33
rect 57 31 59 33
rect 82 31 84 33
<< ndifct0 >>
rect 4 18 6 20
rect 62 21 64 23
rect 14 14 16 16
rect 24 14 26 16
rect 82 22 84 24
rect 71 8 73 10
<< ndifct1 >>
rect 52 22 54 24
rect 34 5 36 7
<< ntiect1 >>
rect 29 65 31 67
<< ptiect1 >>
rect 81 5 83 7
<< pdifct0 >>
rect 4 54 6 56
rect 4 47 6 49
rect 14 54 16 56
rect 24 54 26 56
rect 24 47 26 49
rect 34 55 36 57
rect 61 55 63 57
rect 71 55 73 57
rect 81 55 83 57
rect 81 48 83 50
<< pdifct1 >>
rect 51 46 53 48
<< alu0 >>
rect 2 56 8 57
rect 2 54 4 56
rect 6 54 8 56
rect 2 50 8 54
rect 12 56 18 64
rect 32 57 38 64
rect 12 54 14 56
rect 16 54 18 56
rect 12 53 18 54
rect 22 56 28 57
rect 22 54 24 56
rect 26 54 28 56
rect 32 55 34 57
rect 36 55 38 57
rect 32 54 38 55
rect 42 57 65 58
rect 42 55 61 57
rect 63 55 65 57
rect 42 54 65 55
rect 69 57 75 64
rect 69 55 71 57
rect 73 55 75 57
rect 69 54 75 55
rect 80 57 84 59
rect 80 55 81 57
rect 83 55 84 57
rect 22 50 28 54
rect 42 50 46 54
rect 2 49 17 50
rect 2 47 4 49
rect 6 47 17 49
rect 2 46 17 47
rect 22 49 46 50
rect 22 47 24 49
rect 26 47 46 49
rect 22 46 46 47
rect 13 43 17 46
rect 13 39 22 43
rect 18 34 22 39
rect 18 33 38 34
rect 18 31 19 33
rect 21 31 34 33
rect 36 31 38 33
rect 18 30 38 31
rect 18 25 22 30
rect 3 21 22 25
rect 80 50 84 55
rect 66 48 81 50
rect 83 48 84 50
rect 66 46 84 48
rect 66 33 70 46
rect 66 31 67 33
rect 69 31 76 33
rect 66 29 76 31
rect 72 25 76 29
rect 61 23 65 25
rect 61 21 62 23
rect 64 21 65 23
rect 72 24 86 25
rect 72 22 82 24
rect 84 22 86 24
rect 72 21 86 22
rect 3 20 7 21
rect 3 18 4 20
rect 6 18 7 20
rect 3 16 7 18
rect 61 17 65 21
rect 12 16 18 17
rect 12 14 14 16
rect 16 14 18 16
rect 12 8 18 14
rect 22 16 65 17
rect 22 14 24 16
rect 26 14 65 16
rect 22 13 65 14
rect 70 10 74 12
rect 70 8 71 10
rect 73 8 74 10
<< labels >>
rlabel alu0 5 20 5 20 6 an
rlabel alu0 9 48 9 48 6 an
rlabel alu0 5 51 5 51 6 an
rlabel alu0 28 32 28 32 6 an
rlabel alu0 25 51 25 51 6 n1
rlabel alu0 43 15 43 15 6 n3
rlabel alu0 63 19 63 19 6 n3
rlabel alu0 34 48 34 48 6 n1
rlabel alu0 53 56 53 56 6 n1
rlabel alu0 79 23 79 23 6 bn
rlabel alu0 68 39 68 39 6 bn
rlabel alu0 82 52 82 52 6 bn
rlabel alu1 12 32 12 32 6 a
rlabel alu1 4 36 4 36 6 a
rlabel alu1 44 4 44 4 6 vss
rlabel alu1 44 32 44 32 6 z
rlabel alu1 52 32 52 32 6 c
rlabel alu1 60 40 60 40 6 c
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 68 44 68 6 vdd
rlabel alu1 76 40 76 40 6 b
rlabel alu1 84 36 84 36 6 b
<< end >>
