magic
tech scmos
timestamp 1199543760
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -2 48 52 104
<< pwell >>
rect -2 -4 52 48
<< poly >>
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 11 63 13 65
rect 11 61 19 63
rect 11 59 15 61
rect 17 59 19 61
rect 11 57 19 59
rect 3 51 9 53
rect 23 51 25 65
rect 3 49 5 51
rect 7 49 25 51
rect 3 47 9 49
rect 11 41 19 43
rect 11 39 15 41
rect 17 39 19 41
rect 11 37 19 39
rect 11 35 13 37
rect 23 35 25 49
rect 35 43 37 65
rect 35 41 43 43
rect 35 39 39 41
rect 41 39 43 41
rect 31 37 43 39
rect 31 35 33 37
rect 11 22 13 25
rect 23 12 25 15
rect 31 12 33 15
<< ndif >>
rect 3 31 11 35
rect 3 29 5 31
rect 7 29 11 31
rect 3 25 11 29
rect 13 25 23 35
rect 15 15 23 25
rect 25 15 31 35
rect 33 21 41 35
rect 33 19 37 21
rect 39 19 41 21
rect 33 15 41 19
rect 15 11 21 15
rect 15 9 17 11
rect 19 9 21 11
rect 15 7 21 9
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 39 91 45 93
rect 39 89 41 91
rect 43 89 45 91
rect 39 85 45 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 65 23 85
rect 25 81 35 85
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 65 35 69
rect 37 65 45 85
<< alu1 >>
rect -2 91 52 100
rect -2 89 17 91
rect 19 89 41 91
rect 43 89 52 91
rect -2 88 52 89
rect 4 81 8 82
rect 4 79 5 81
rect 7 79 8 81
rect 4 78 8 79
rect 5 72 7 78
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 52 7 68
rect 18 62 22 82
rect 14 61 22 62
rect 14 59 15 61
rect 17 59 22 61
rect 14 58 22 59
rect 4 51 8 52
rect 4 49 5 51
rect 7 49 8 51
rect 4 48 8 49
rect 5 32 7 48
rect 18 42 22 58
rect 14 41 22 42
rect 14 39 15 41
rect 17 39 22 41
rect 14 38 22 39
rect 4 31 8 32
rect 4 29 5 31
rect 7 29 8 31
rect 4 28 8 29
rect 18 18 22 38
rect 28 81 32 82
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 22 32 69
rect 38 41 42 82
rect 38 39 39 41
rect 41 39 42 41
rect 38 28 42 39
rect 28 21 40 22
rect 28 19 37 21
rect 39 19 40 21
rect 28 18 40 19
rect -2 11 52 12
rect -2 9 17 11
rect 19 9 52 11
rect -2 7 52 9
rect -2 5 5 7
rect 7 5 29 7
rect 31 5 43 7
rect 45 5 52 7
rect -2 0 52 5
<< ptie >>
rect 3 7 9 15
rect 27 7 47 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 27 5 29 7
rect 31 5 43 7
rect 45 5 47 7
rect 27 3 47 5
<< nmos >>
rect 11 25 13 35
rect 23 15 25 35
rect 31 15 33 35
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
<< polyct1 >>
rect 15 59 17 61
rect 5 49 7 51
rect 15 39 17 41
rect 39 39 41 41
<< ndifct1 >>
rect 5 29 7 31
rect 37 19 39 21
rect 17 9 19 11
<< ptiect1 >>
rect 5 5 7 7
rect 29 5 31 7
rect 43 5 45 7
<< pdifct1 >>
rect 17 89 19 91
rect 41 89 43 91
rect 5 79 7 81
rect 5 69 7 71
rect 29 79 31 81
rect 29 69 31 71
<< labels >>
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 50 30 50 6 q
rlabel alu1 25 94 25 94 6 vdd
rlabel alu1 40 55 40 55 6 i0
<< end >>
