magic
tech scmos
timestamp 1199202680
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 9 62 11 67
rect 19 62 21 67
rect 29 62 31 67
rect 39 62 41 67
rect 50 52 52 57
rect 60 52 62 57
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 50 35 52 38
rect 60 35 62 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 31 35
rect 19 31 27 33
rect 29 31 31 33
rect 19 29 31 31
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 33 52 35
rect 56 33 62 35
rect 36 31 43 33
rect 45 31 47 33
rect 36 29 47 31
rect 56 31 58 33
rect 60 31 62 33
rect 56 29 62 31
rect 36 26 38 29
rect 12 8 14 13
rect 19 8 21 13
rect 29 8 31 13
rect 36 8 38 13
<< ndif >>
rect 3 13 12 26
rect 14 13 19 26
rect 21 17 29 26
rect 21 15 24 17
rect 26 15 29 17
rect 21 13 29 15
rect 31 13 36 26
rect 38 13 47 26
rect 3 7 10 13
rect 3 5 6 7
rect 8 5 10 7
rect 3 3 10 5
rect 40 7 47 13
rect 40 5 42 7
rect 44 5 47 7
rect 40 3 47 5
<< pdif >>
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 38 9 58
rect 11 57 19 62
rect 11 55 14 57
rect 16 55 19 57
rect 11 49 19 55
rect 11 47 14 49
rect 16 47 19 49
rect 11 38 19 47
rect 21 60 29 62
rect 21 58 24 60
rect 26 58 29 60
rect 21 38 29 58
rect 31 57 39 62
rect 31 55 34 57
rect 36 55 39 57
rect 31 49 39 55
rect 31 47 34 49
rect 36 47 39 49
rect 31 38 39 47
rect 41 60 48 62
rect 41 58 44 60
rect 46 58 48 60
rect 41 52 48 58
rect 41 38 50 52
rect 52 49 60 52
rect 52 47 55 49
rect 57 47 60 49
rect 52 38 60 47
rect 62 50 70 52
rect 62 48 65 50
rect 67 48 70 50
rect 62 42 70 48
rect 62 40 65 42
rect 67 40 70 42
rect 62 38 70 40
<< alu1 >>
rect -2 67 74 72
rect -2 65 54 67
rect 56 65 65 67
rect 67 65 74 67
rect -2 64 74 65
rect 33 57 38 59
rect 33 55 34 57
rect 36 55 38 57
rect 33 50 38 55
rect 2 49 59 50
rect 2 47 14 49
rect 16 47 34 49
rect 36 47 55 49
rect 57 47 59 49
rect 2 46 59 47
rect 2 18 6 46
rect 25 38 57 42
rect 10 33 21 35
rect 10 31 11 33
rect 13 31 21 33
rect 10 29 21 31
rect 25 33 31 38
rect 53 34 57 38
rect 25 31 27 33
rect 29 31 31 33
rect 25 30 31 31
rect 41 33 47 34
rect 41 31 43 33
rect 45 31 47 33
rect 17 26 21 29
rect 41 26 47 31
rect 53 33 63 34
rect 53 31 58 33
rect 60 31 63 33
rect 53 30 63 31
rect 17 22 47 26
rect 2 17 31 18
rect 2 15 24 17
rect 26 15 31 17
rect 2 14 31 15
rect -2 7 74 8
rect -2 5 6 7
rect 8 5 42 7
rect 44 5 54 7
rect 56 5 65 7
rect 67 5 74 7
rect -2 0 74 5
<< ptie >>
rect 52 7 69 9
rect 52 5 54 7
rect 56 5 65 7
rect 67 5 69 7
rect 52 3 69 5
<< ntie >>
rect 52 67 69 69
rect 52 65 54 67
rect 56 65 65 67
rect 67 65 69 67
rect 52 63 69 65
<< nmos >>
rect 12 13 14 26
rect 19 13 21 26
rect 29 13 31 26
rect 36 13 38 26
<< pmos >>
rect 9 38 11 62
rect 19 38 21 62
rect 29 38 31 62
rect 39 38 41 62
rect 50 38 52 52
rect 60 38 62 52
<< polyct1 >>
rect 11 31 13 33
rect 27 31 29 33
rect 43 31 45 33
rect 58 31 60 33
<< ndifct1 >>
rect 24 15 26 17
rect 6 5 8 7
rect 42 5 44 7
<< ntiect1 >>
rect 54 65 56 67
rect 65 65 67 67
<< ptiect1 >>
rect 54 5 56 7
rect 65 5 67 7
<< pdifct0 >>
rect 4 58 6 60
rect 14 55 16 57
rect 24 58 26 60
rect 44 58 46 60
rect 65 48 67 50
rect 65 40 67 42
<< pdifct1 >>
rect 14 47 16 49
rect 34 55 36 57
rect 34 47 36 49
rect 55 47 57 49
<< alu0 >>
rect 3 60 7 64
rect 3 58 4 60
rect 6 58 7 60
rect 23 60 27 64
rect 3 56 7 58
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 23 58 24 60
rect 26 58 27 60
rect 43 60 47 64
rect 23 56 27 58
rect 13 50 17 55
rect 43 58 44 60
rect 46 58 47 60
rect 43 56 47 58
rect 64 50 68 64
rect 64 48 65 50
rect 67 48 68 50
rect 64 42 68 48
rect 64 40 65 42
rect 67 40 68 42
rect 64 38 68 40
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 24 20 24 6 a
rlabel alu1 28 24 28 24 6 a
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 40 44 40 6 b
rlabel alu1 52 40 52 40 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 32 60 32 6 b
<< end >>
