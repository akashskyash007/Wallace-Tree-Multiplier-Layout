magic
tech scmos
timestamp 1199201978
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 9 66 11 70
rect 21 55 23 60
rect 9 35 11 38
rect 21 35 23 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 21 33 27 35
rect 21 31 23 33
rect 25 31 27 33
rect 21 29 27 31
rect 9 26 11 29
rect 21 26 23 29
rect 9 7 11 12
rect 21 11 23 16
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 12 9 15
rect 11 16 21 26
rect 23 24 30 26
rect 23 22 26 24
rect 28 22 30 24
rect 23 20 30 22
rect 23 16 28 20
rect 11 14 15 16
rect 17 14 19 16
rect 11 12 19 14
<< pdif >>
rect 13 67 19 69
rect 13 66 15 67
rect 4 59 9 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 4 38 9 46
rect 11 65 15 66
rect 17 65 19 67
rect 11 55 19 65
rect 11 38 21 55
rect 23 51 28 55
rect 23 49 30 51
rect 23 47 26 49
rect 28 47 30 49
rect 23 45 30 47
rect 23 38 28 45
<< alu1 >>
rect -2 67 34 72
rect -2 65 15 67
rect 17 65 25 67
rect 27 65 34 67
rect -2 64 34 65
rect 2 57 15 59
rect 2 55 4 57
rect 6 55 15 57
rect 2 54 15 55
rect 2 50 6 54
rect 2 48 4 50
rect 2 26 6 48
rect 26 35 30 43
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 17 7 22
rect 18 33 30 35
rect 18 31 23 33
rect 25 31 30 33
rect 18 29 30 31
rect 2 15 4 17
rect 6 15 7 17
rect 2 13 7 15
rect -2 7 34 8
rect -2 5 25 7
rect 27 5 34 7
rect -2 0 34 5
<< ptie >>
rect 23 7 29 9
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< ntie >>
rect 23 67 29 69
rect 23 65 25 67
rect 27 65 29 67
rect 23 63 29 65
<< nmos >>
rect 9 12 11 26
rect 21 16 23 26
<< pmos >>
rect 9 38 11 66
rect 21 38 23 55
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 23 31 25 33
<< ndifct0 >>
rect 26 22 28 24
rect 15 14 17 16
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
<< ntiect1 >>
rect 25 65 27 67
<< ptiect1 >>
rect 25 5 27 7
<< pdifct0 >>
rect 26 47 28 49
<< pdifct1 >>
rect 4 55 6 57
rect 4 48 6 50
rect 15 65 17 67
<< alu0 >>
rect 6 46 7 54
rect 10 49 30 50
rect 10 47 26 49
rect 28 47 30 49
rect 10 46 30 47
rect 10 33 14 46
rect 10 31 11 33
rect 13 31 14 33
rect 10 25 14 31
rect 10 24 30 25
rect 10 22 26 24
rect 28 22 30 24
rect 10 21 30 22
rect 13 16 19 17
rect 13 14 15 16
rect 17 14 19 16
rect 13 8 19 14
<< labels >>
rlabel alu0 12 35 12 35 6 an
rlabel alu0 20 23 20 23 6 an
rlabel alu0 20 48 20 48 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 12 56 12 56 6 z
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 20 32 20 32 6 a
rlabel alu1 28 36 28 36 6 a
<< end >>
