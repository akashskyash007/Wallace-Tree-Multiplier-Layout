magic
tech scmos
timestamp 1199542387
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 45 94 47 98
rect 57 94 59 98
rect 11 83 13 87
rect 23 83 25 87
rect 35 83 37 87
rect 11 43 13 63
rect 23 53 25 63
rect 17 51 25 53
rect 17 49 19 51
rect 21 49 25 51
rect 17 47 25 49
rect 7 41 15 43
rect 7 39 9 41
rect 11 39 15 41
rect 7 37 15 39
rect 13 34 15 37
rect 21 34 23 47
rect 35 43 37 63
rect 67 82 73 84
rect 67 80 69 82
rect 71 80 73 82
rect 67 78 73 80
rect 67 75 69 78
rect 45 43 47 55
rect 57 43 59 55
rect 27 41 37 43
rect 43 41 63 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 43 39 59 41
rect 61 39 63 41
rect 43 37 63 39
rect 29 34 31 37
rect 43 25 45 37
rect 55 25 57 37
rect 67 25 69 55
rect 13 11 15 15
rect 21 11 23 15
rect 29 11 31 15
rect 67 11 69 15
rect 43 2 45 6
rect 55 2 57 6
<< ndif >>
rect 5 21 13 34
rect 5 19 7 21
rect 9 19 13 21
rect 5 15 13 19
rect 15 15 21 34
rect 23 15 29 34
rect 31 25 41 34
rect 31 15 43 25
rect 33 11 43 15
rect 33 9 37 11
rect 39 9 43 11
rect 33 6 43 9
rect 45 21 55 25
rect 45 19 49 21
rect 51 19 55 21
rect 45 6 55 19
rect 57 15 67 25
rect 69 21 77 25
rect 69 19 73 21
rect 75 19 77 21
rect 69 15 77 19
rect 57 11 65 15
rect 57 9 61 11
rect 63 9 65 11
rect 57 6 65 9
<< pdif >>
rect 37 94 43 95
rect 61 94 67 95
rect 37 93 45 94
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 37 91 39 93
rect 41 91 45 93
rect 37 89 45 91
rect 15 83 21 89
rect 39 83 45 89
rect 3 81 11 83
rect 3 79 5 81
rect 7 79 11 81
rect 3 63 11 79
rect 13 63 23 83
rect 25 81 35 83
rect 25 79 29 81
rect 31 79 35 81
rect 25 63 35 79
rect 37 63 45 83
rect 39 55 45 63
rect 47 71 57 94
rect 47 69 51 71
rect 53 69 57 71
rect 47 61 57 69
rect 47 59 51 61
rect 53 59 57 61
rect 47 55 57 59
rect 59 93 67 94
rect 59 91 63 93
rect 65 91 67 93
rect 59 89 67 91
rect 59 75 65 89
rect 59 55 67 75
rect 69 71 77 75
rect 69 69 73 71
rect 75 69 77 71
rect 69 61 77 69
rect 69 59 73 61
rect 75 59 77 61
rect 69 55 77 59
<< alu1 >>
rect -2 93 82 100
rect -2 91 39 93
rect 41 91 63 93
rect 65 91 82 93
rect -2 89 17 91
rect 19 89 82 91
rect -2 88 82 89
rect 67 82 73 83
rect 3 81 69 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 80 69 81
rect 71 80 73 82
rect 31 79 73 80
rect 3 78 72 79
rect 8 41 12 73
rect 8 39 9 41
rect 11 39 12 41
rect 8 27 12 39
rect 18 51 22 73
rect 18 49 19 51
rect 21 49 22 51
rect 18 27 22 49
rect 28 41 32 73
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 22 42 78
rect 5 21 42 22
rect 5 19 7 21
rect 9 19 42 21
rect 5 18 42 19
rect 48 72 52 73
rect 48 71 55 72
rect 48 69 51 71
rect 53 69 55 71
rect 48 68 55 69
rect 72 71 76 73
rect 72 69 73 71
rect 75 69 76 71
rect 48 62 52 68
rect 48 61 55 62
rect 48 59 51 61
rect 53 59 55 61
rect 48 58 55 59
rect 72 61 76 69
rect 72 59 73 61
rect 75 59 76 61
rect 48 21 52 58
rect 72 42 76 59
rect 57 41 76 42
rect 57 39 59 41
rect 61 39 76 41
rect 57 38 76 39
rect 48 19 49 21
rect 51 19 52 21
rect 48 17 52 19
rect 72 21 76 38
rect 72 19 73 21
rect 75 19 76 21
rect 72 17 76 19
rect -2 11 82 12
rect -2 9 37 11
rect 39 9 61 11
rect 63 9 82 11
rect -2 7 82 9
rect -2 5 5 7
rect 7 5 13 7
rect 15 5 21 7
rect 23 5 82 7
rect -2 0 82 5
<< ptie >>
rect 3 7 25 9
rect 3 5 5 7
rect 7 5 13 7
rect 15 5 21 7
rect 23 5 25 7
rect 3 3 25 5
<< nmos >>
rect 13 15 15 34
rect 21 15 23 34
rect 29 15 31 34
rect 43 6 45 25
rect 55 6 57 25
rect 67 15 69 25
<< pmos >>
rect 11 63 13 83
rect 23 63 25 83
rect 35 63 37 83
rect 45 55 47 94
rect 57 55 59 94
rect 67 55 69 75
<< polyct1 >>
rect 19 49 21 51
rect 9 39 11 41
rect 69 80 71 82
rect 29 39 31 41
rect 59 39 61 41
<< ndifct1 >>
rect 7 19 9 21
rect 37 9 39 11
rect 49 19 51 21
rect 73 19 75 21
rect 61 9 63 11
<< ptiect1 >>
rect 5 5 7 7
rect 13 5 15 7
rect 21 5 23 7
<< pdifct1 >>
rect 17 89 19 91
rect 39 91 41 93
rect 5 79 7 81
rect 29 79 31 81
rect 51 69 53 71
rect 51 59 53 61
rect 63 91 65 93
rect 73 69 75 71
rect 73 59 75 61
<< labels >>
rlabel alu1 10 50 10 50 6 i0
rlabel alu1 30 50 30 50 6 i1
rlabel polyct1 20 50 20 50 6 i2
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 50 45 50 45 6 nq
rlabel alu1 40 94 40 94 6 vdd
<< end >>
