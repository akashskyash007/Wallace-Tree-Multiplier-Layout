magic
tech scmos
timestamp 1199203318
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 33 70 35 74
rect 40 70 42 74
rect 47 70 49 74
rect 54 70 56 74
rect 64 70 66 74
rect 71 70 73 74
rect 78 70 80 74
rect 85 70 87 74
rect 9 61 11 65
rect 19 63 21 68
rect 9 39 11 42
rect 19 39 21 42
rect 33 39 35 42
rect 9 37 21 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 28 37 35 39
rect 28 35 30 37
rect 32 36 35 37
rect 32 35 34 36
rect 28 33 34 35
rect 9 30 11 33
rect 28 22 30 33
rect 40 32 42 42
rect 47 39 49 42
rect 54 39 56 42
rect 64 39 66 42
rect 47 36 50 39
rect 54 37 66 39
rect 38 30 44 32
rect 38 28 40 30
rect 42 28 44 30
rect 38 26 44 28
rect 48 31 50 36
rect 58 35 60 37
rect 62 35 64 37
rect 58 33 64 35
rect 48 29 54 31
rect 48 27 50 29
rect 52 27 54 29
rect 38 22 40 26
rect 48 25 54 27
rect 50 22 52 25
rect 60 22 62 33
rect 71 31 73 42
rect 78 33 80 42
rect 85 39 87 42
rect 85 37 94 39
rect 88 35 90 37
rect 92 35 94 37
rect 88 33 94 35
rect 78 31 84 33
rect 68 29 74 31
rect 68 27 70 29
rect 72 27 74 29
rect 78 29 80 31
rect 82 29 84 31
rect 78 27 84 29
rect 68 25 74 27
rect 9 6 11 10
rect 28 9 30 14
rect 38 9 40 14
rect 50 9 52 14
rect 60 9 62 14
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 22 26 30
rect 11 20 28 22
rect 11 18 14 20
rect 16 18 28 20
rect 11 14 28 18
rect 30 20 38 22
rect 30 18 33 20
rect 35 18 38 20
rect 30 14 38 18
rect 40 14 50 22
rect 52 20 60 22
rect 52 18 55 20
rect 57 18 60 20
rect 52 14 60 18
rect 62 14 71 22
rect 11 11 26 14
rect 11 10 15 11
rect 13 9 15 10
rect 17 9 22 11
rect 24 9 26 11
rect 42 11 48 14
rect 42 9 44 11
rect 46 9 48 11
rect 64 11 71 14
rect 64 9 66 11
rect 68 9 71 11
rect 13 7 26 9
rect 42 7 48 9
rect 64 7 71 9
<< pdif >>
rect 23 68 33 70
rect 23 66 26 68
rect 28 66 33 68
rect 23 63 33 66
rect 14 61 19 63
rect 2 59 9 61
rect 2 57 4 59
rect 6 57 9 59
rect 2 52 9 57
rect 2 50 4 52
rect 6 50 9 52
rect 2 42 9 50
rect 11 53 19 61
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 42 33 63
rect 35 42 40 70
rect 42 42 47 70
rect 49 42 54 70
rect 56 61 64 70
rect 56 59 59 61
rect 61 59 64 61
rect 56 42 64 59
rect 66 42 71 70
rect 73 42 78 70
rect 80 42 85 70
rect 87 68 94 70
rect 87 66 90 68
rect 92 66 94 68
rect 87 61 94 66
rect 87 59 90 61
rect 92 59 94 61
rect 87 42 94 59
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 13 46 17 51
rect 2 44 14 46
rect 16 44 17 46
rect 2 42 17 44
rect 2 30 6 42
rect 74 54 78 63
rect 2 28 15 30
rect 2 26 4 28
rect 6 26 15 28
rect 2 21 7 26
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect 29 50 94 54
rect 29 37 33 50
rect 29 35 30 37
rect 32 35 33 37
rect 29 33 33 35
rect 39 42 79 46
rect 39 30 43 42
rect 73 38 79 42
rect 49 37 64 38
rect 49 35 60 37
rect 62 35 64 37
rect 49 34 64 35
rect 73 34 83 38
rect 79 31 83 34
rect 89 37 94 50
rect 89 35 90 37
rect 92 35 94 37
rect 89 33 94 35
rect 39 28 40 30
rect 42 28 43 30
rect 39 26 43 28
rect 48 29 74 30
rect 48 27 50 29
rect 52 27 70 29
rect 72 27 74 29
rect 79 29 80 31
rect 82 29 83 31
rect 79 27 83 29
rect 48 26 74 27
rect 66 17 70 26
rect -2 11 98 12
rect -2 9 15 11
rect 17 9 22 11
rect 24 9 44 11
rect 46 9 66 11
rect 68 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 9 10 11 30
rect 28 14 30 22
rect 38 14 40 22
rect 50 14 52 22
rect 60 14 62 22
<< pmos >>
rect 9 42 11 61
rect 19 42 21 63
rect 33 42 35 70
rect 40 42 42 70
rect 47 42 49 70
rect 54 42 56 70
rect 64 42 66 70
rect 71 42 73 70
rect 78 42 80 70
rect 85 42 87 70
<< polyct0 >>
rect 17 35 19 37
<< polyct1 >>
rect 30 35 32 37
rect 40 28 42 30
rect 60 35 62 37
rect 50 27 52 29
rect 90 35 92 37
rect 70 27 72 29
rect 80 29 82 31
<< ndifct0 >>
rect 14 18 16 20
rect 33 18 35 20
rect 55 18 57 20
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
rect 15 9 17 11
rect 22 9 24 11
rect 44 9 46 11
rect 66 9 68 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 26 66 28 68
rect 4 57 6 59
rect 4 50 6 52
rect 59 59 61 61
rect 90 66 92 68
rect 90 59 92 61
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
<< alu0 >>
rect 2 59 8 68
rect 24 66 26 68
rect 28 66 30 68
rect 24 65 30 66
rect 88 66 90 68
rect 92 66 94 68
rect 2 57 4 59
rect 6 57 8 59
rect 2 52 8 57
rect 21 61 63 62
rect 21 59 59 61
rect 61 59 63 61
rect 21 58 63 59
rect 2 50 4 52
rect 6 50 8 52
rect 2 49 8 50
rect 21 38 25 58
rect 88 61 94 66
rect 88 59 90 61
rect 92 59 94 61
rect 88 58 94 59
rect 15 37 25 38
rect 15 35 17 37
rect 19 35 25 37
rect 15 34 25 35
rect 13 20 17 22
rect 13 18 14 20
rect 16 18 17 20
rect 13 12 17 18
rect 21 21 25 34
rect 21 20 59 21
rect 21 18 33 20
rect 35 18 55 20
rect 57 18 59 20
rect 21 17 59 18
<< labels >>
rlabel alu0 20 36 20 36 6 zn
rlabel alu0 40 19 40 19 6 zn
rlabel alu0 42 60 42 60 6 zn
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 52 28 52 28 6 c
rlabel alu1 44 44 44 44 6 b
rlabel alu1 52 36 52 36 6 d
rlabel alu1 52 44 52 44 6 b
rlabel alu1 44 52 44 52 6 a
rlabel alu1 52 52 52 52 6 a
rlabel alu1 36 52 36 52 6 a
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 60 28 60 28 6 c
rlabel alu1 68 20 68 20 6 c
rlabel alu1 68 24 68 24 6 c
rlabel alu1 60 36 60 36 6 d
rlabel alu1 60 44 60 44 6 b
rlabel alu1 68 44 68 44 6 b
rlabel alu1 76 40 76 40 6 b
rlabel alu1 68 52 68 52 6 a
rlabel alu1 60 52 60 52 6 a
rlabel alu1 76 56 76 56 6 a
rlabel alu1 92 40 92 40 6 a
rlabel alu1 84 52 84 52 6 a
<< end >>
