magic
tech scmos
timestamp 1199542525
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 23 95 25 98
rect 33 95 35 98
rect 45 95 47 98
rect 57 95 59 98
rect 11 85 13 88
rect 11 41 13 65
rect 23 53 25 55
rect 17 51 25 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 33 43 35 55
rect 45 53 47 55
rect 57 53 59 55
rect 45 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 57 51 63 53
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 27 41 35 43
rect 11 39 29 41
rect 31 39 47 41
rect 11 25 13 39
rect 27 37 33 39
rect 17 31 23 33
rect 17 29 19 31
rect 21 29 23 31
rect 29 31 35 33
rect 29 29 31 31
rect 33 29 35 31
rect 17 27 25 29
rect 29 27 35 29
rect 23 25 25 27
rect 33 25 35 27
rect 45 25 47 39
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 57 27 63 29
rect 57 25 59 27
rect 11 12 13 15
rect 23 2 25 5
rect 33 2 35 5
rect 45 2 47 5
rect 57 2 59 5
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 15 11 23 15
rect 15 9 17 11
rect 19 9 23 11
rect 15 5 23 9
rect 25 5 33 25
rect 35 21 45 25
rect 35 19 39 21
rect 41 19 45 21
rect 35 5 45 19
rect 47 5 57 25
rect 59 11 67 25
rect 59 9 63 11
rect 65 9 67 11
rect 59 5 67 9
<< pdif >>
rect 15 91 23 95
rect 15 89 17 91
rect 19 89 23 91
rect 15 85 23 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 65 23 85
rect 15 55 23 65
rect 25 55 33 95
rect 35 71 45 95
rect 35 69 39 71
rect 41 69 45 71
rect 35 61 45 69
rect 35 59 39 61
rect 41 59 45 61
rect 35 55 45 59
rect 47 55 57 95
rect 59 91 67 95
rect 59 89 63 91
rect 65 89 67 91
rect 59 55 67 89
<< alu1 >>
rect -2 91 72 100
rect -2 89 17 91
rect 19 89 63 91
rect 65 89 72 91
rect -2 88 72 89
rect 4 81 8 82
rect 4 79 5 81
rect 7 79 51 81
rect 4 78 8 79
rect 5 72 7 78
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 22 7 68
rect 18 51 22 72
rect 18 49 19 51
rect 21 49 22 51
rect 18 31 22 49
rect 28 41 32 72
rect 28 39 29 41
rect 31 39 32 41
rect 28 38 32 39
rect 38 71 42 72
rect 38 69 39 71
rect 41 69 42 71
rect 38 61 42 69
rect 38 59 39 61
rect 41 59 42 61
rect 38 42 42 59
rect 49 52 51 79
rect 48 51 52 52
rect 48 49 49 51
rect 51 49 52 51
rect 48 48 52 49
rect 58 51 62 82
rect 58 49 59 51
rect 61 49 62 51
rect 38 38 44 42
rect 40 32 44 38
rect 18 29 19 31
rect 21 29 22 31
rect 18 28 22 29
rect 30 31 34 32
rect 30 29 31 31
rect 33 29 34 31
rect 30 28 34 29
rect 40 28 52 32
rect 58 31 62 49
rect 58 29 59 31
rect 61 29 62 31
rect 4 21 8 22
rect 30 21 32 28
rect 40 22 44 28
rect 4 19 5 21
rect 7 19 32 21
rect 38 21 44 22
rect 38 19 39 21
rect 41 19 44 21
rect 4 18 8 19
rect 38 18 44 19
rect 58 18 62 29
rect -2 11 72 12
rect -2 9 17 11
rect 19 9 63 11
rect 65 9 72 11
rect -2 0 72 9
<< nmos >>
rect 11 15 13 25
rect 23 5 25 25
rect 33 5 35 25
rect 45 5 47 25
rect 57 5 59 25
<< pmos >>
rect 11 65 13 85
rect 23 55 25 95
rect 33 55 35 95
rect 45 55 47 95
rect 57 55 59 95
<< polyct1 >>
rect 19 49 21 51
rect 49 49 51 51
rect 59 49 61 51
rect 29 39 31 41
rect 19 29 21 31
rect 31 29 33 31
rect 59 29 61 31
<< ndifct1 >>
rect 5 19 7 21
rect 17 9 19 11
rect 39 19 41 21
rect 63 9 65 11
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 5 69 7 71
rect 39 69 41 71
rect 39 59 41 61
rect 63 89 65 91
<< labels >>
rlabel alu1 30 55 30 55 6 cmd
rlabel polyct1 20 50 20 50 6 i0
rlabel ndifct1 40 20 40 20 6 nq
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 50 30 50 30 6 nq
rlabel alu1 40 55 40 55 6 nq
rlabel alu1 35 94 35 94 6 vdd
rlabel polyct1 60 50 60 50 6 i1
<< end >>
