magic
tech scmos
timestamp 1199201993
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 69 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 22 39
rect 9 35 18 37
rect 20 35 22 37
rect 9 33 22 35
rect 26 37 32 39
rect 26 35 28 37
rect 30 35 32 37
rect 26 33 32 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 9 11 11 16
rect 19 11 21 16
rect 29 10 31 15
<< ndif >>
rect 2 27 9 30
rect 2 25 4 27
rect 6 25 9 27
rect 2 20 9 25
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 21 19 30
rect 11 19 14 21
rect 16 19 19 21
rect 11 16 19 19
rect 21 20 29 30
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 23 15 29 16
rect 31 28 38 30
rect 31 26 34 28
rect 36 26 38 28
rect 31 21 38 26
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
rect 31 15 36 17
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 69 27 70
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 62 36 69
rect 31 60 38 62
rect 31 58 34 60
rect 36 58 38 60
rect 31 53 38 58
rect 31 51 34 53
rect 36 51 38 53
rect 31 49 38 51
rect 31 42 36 49
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 37 6 50
rect 17 42 31 46
rect 2 33 14 37
rect 10 23 14 33
rect 26 37 31 42
rect 26 35 28 37
rect 30 35 31 37
rect 26 33 31 35
rect 10 21 17 23
rect 10 19 14 21
rect 16 19 17 21
rect 10 17 17 19
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 15 31 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 69
<< polyct0 >>
rect 18 35 20 37
<< polyct1 >>
rect 28 35 30 37
<< ndifct0 >>
rect 4 25 6 27
rect 4 18 6 20
rect 24 18 26 20
rect 34 26 36 28
rect 34 19 36 21
<< ndifct1 >>
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 65 26 67
rect 24 58 26 60
rect 34 58 36 60
rect 34 51 36 53
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 23 67 27 68
rect 23 65 24 67
rect 26 65 27 67
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 23 60 27 65
rect 23 58 24 60
rect 26 58 27 60
rect 23 56 27 58
rect 33 60 38 62
rect 33 58 34 60
rect 36 58 38 60
rect 33 53 38 58
rect 33 51 34 53
rect 36 51 38 53
rect 33 49 38 51
rect 17 37 21 39
rect 3 27 7 29
rect 3 25 4 27
rect 6 25 7 27
rect 3 20 7 25
rect 3 18 4 20
rect 6 18 7 20
rect 3 12 7 18
rect 17 35 18 37
rect 20 35 21 37
rect 17 30 21 35
rect 34 30 38 49
rect 17 28 38 30
rect 17 26 34 28
rect 36 26 38 28
rect 23 20 27 22
rect 23 18 24 20
rect 26 18 27 20
rect 23 12 27 18
rect 33 21 37 26
rect 33 19 34 21
rect 36 19 37 21
rect 33 17 37 19
<< labels >>
rlabel alu0 19 32 19 32 6 an
rlabel alu0 35 23 35 23 6 an
rlabel alu0 36 44 36 44 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 40 28 40 6 a
rlabel alu1 20 44 20 44 6 a
rlabel alu1 20 74 20 74 6 vdd
<< end >>
