magic
tech scmos
timestamp 1199201853
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 51 70 53 74
rect 61 70 63 74
rect 9 40 11 43
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 19 39 21 43
rect 29 39 31 43
rect 19 37 31 39
rect 39 40 41 43
rect 51 40 53 43
rect 61 40 63 43
rect 39 38 54 40
rect 19 35 27 37
rect 29 35 31 37
rect 19 33 31 35
rect 41 37 54 38
rect 41 35 43 37
rect 45 35 54 37
rect 20 29 22 33
rect 35 29 37 34
rect 41 33 54 35
rect 58 38 64 40
rect 58 36 60 38
rect 62 36 64 38
rect 58 34 64 36
rect 42 29 44 33
rect 52 29 54 33
rect 59 29 61 34
rect 20 9 22 14
rect 35 8 37 16
rect 42 12 44 16
rect 52 12 54 16
rect 59 8 61 16
rect 35 6 61 8
<< ndif >>
rect 15 23 20 29
rect 13 21 20 23
rect 13 19 15 21
rect 17 19 20 21
rect 13 17 20 19
rect 15 14 20 17
rect 22 16 35 29
rect 37 16 42 29
rect 44 21 52 29
rect 44 19 47 21
rect 49 19 52 21
rect 44 16 52 19
rect 54 16 59 29
rect 61 16 69 29
rect 22 14 33 16
rect 24 12 27 14
rect 29 12 33 14
rect 24 10 33 12
rect 63 11 69 16
rect 63 9 65 11
rect 67 9 69 11
rect 63 7 69 9
<< pdif >>
rect 43 71 49 73
rect 43 70 45 71
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 43 9 59
rect 11 62 19 70
rect 11 60 14 62
rect 16 60 19 62
rect 11 43 19 60
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 43 29 51
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 43 39 52
rect 41 69 45 70
rect 47 70 49 71
rect 47 69 51 70
rect 41 43 51 69
rect 53 61 61 70
rect 53 59 56 61
rect 58 59 61 61
rect 53 54 61 59
rect 53 52 56 54
rect 58 52 61 54
rect 53 43 61 52
rect 63 68 70 70
rect 63 66 66 68
rect 68 66 70 68
rect 63 60 70 66
rect 63 58 66 60
rect 68 58 70 60
rect 63 43 70 58
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 71 74 79
rect -2 69 45 71
rect 47 69 74 71
rect -2 68 74 69
rect 2 53 28 55
rect 2 51 24 53
rect 26 51 28 53
rect 2 50 28 51
rect 2 22 6 50
rect 42 46 46 55
rect 10 42 63 46
rect 10 38 14 42
rect 57 38 63 42
rect 10 36 11 38
rect 13 36 14 38
rect 10 34 14 36
rect 25 37 31 38
rect 25 35 27 37
rect 29 35 31 37
rect 25 30 31 35
rect 17 26 31 30
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 30 47 35
rect 57 36 60 38
rect 62 36 63 38
rect 57 34 63 36
rect 41 26 55 30
rect 2 21 55 22
rect 2 19 15 21
rect 17 19 47 21
rect 49 19 55 21
rect 2 18 55 19
rect -2 11 74 12
rect -2 9 65 11
rect 67 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 20 14 22 29
rect 35 16 37 29
rect 42 16 44 29
rect 52 16 54 29
rect 59 16 61 29
<< pmos >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
rect 51 43 53 70
rect 61 43 63 70
<< polyct1 >>
rect 11 36 13 38
rect 27 35 29 37
rect 43 35 45 37
rect 60 36 62 38
<< ndifct0 >>
rect 27 12 29 14
<< ndifct1 >>
rect 15 19 17 21
rect 47 19 49 21
rect 65 9 67 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 60 16 62
rect 34 59 36 61
rect 34 52 36 54
rect 56 59 58 61
rect 56 52 58 54
rect 66 66 68 68
rect 66 58 68 60
<< pdifct1 >>
rect 24 51 26 53
rect 45 69 47 71
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 65 66 66 68
rect 68 66 69 68
rect 2 59 4 61
rect 6 59 8 61
rect 12 62 59 63
rect 12 60 14 62
rect 16 61 59 62
rect 16 60 34 61
rect 12 59 34 60
rect 36 59 56 61
rect 58 59 59 61
rect 2 58 8 59
rect 33 54 37 59
rect 33 52 34 54
rect 36 52 37 54
rect 33 50 37 52
rect 55 54 59 59
rect 65 60 69 66
rect 65 58 66 60
rect 68 58 69 60
rect 65 56 69 58
rect 55 52 56 54
rect 58 52 59 54
rect 55 50 59 52
rect 25 14 31 15
rect 25 12 27 14
rect 29 12 31 14
<< labels >>
rlabel alu0 35 56 35 56 6 n1
rlabel alu0 57 56 57 56 6 n1
rlabel alu0 35 61 35 61 6 n1
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 32 28 32 6 b
rlabel alu1 28 44 28 44 6 a1
rlabel alu1 20 44 20 44 6 a1
rlabel alu1 20 52 20 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 44 32 44 32 6 a2
rlabel alu1 52 28 52 28 6 a2
rlabel alu1 52 44 52 44 6 a1
rlabel alu1 36 44 36 44 6 a1
rlabel alu1 44 48 44 48 6 a1
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 40 60 40 6 a1
<< end >>
