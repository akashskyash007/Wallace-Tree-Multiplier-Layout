magic
tech scmos
timestamp 1199542816
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -5 48 105 105
<< pwell >>
rect -5 -5 105 48
<< poly >>
rect 19 94 21 98
rect 27 94 29 98
rect 35 94 37 98
rect 43 94 45 98
rect 63 94 65 98
rect 75 94 77 98
rect 19 53 21 56
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 11 47 23 49
rect 11 25 13 47
rect 27 43 29 56
rect 35 53 37 56
rect 43 53 45 56
rect 87 76 89 80
rect 35 51 39 53
rect 43 51 49 53
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 23 37 33 39
rect 23 25 25 37
rect 37 33 39 51
rect 47 43 49 51
rect 63 43 65 55
rect 75 43 77 55
rect 87 53 89 56
rect 81 51 89 53
rect 81 49 83 51
rect 85 49 89 51
rect 81 47 89 49
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 63 41 97 43
rect 63 39 93 41
rect 95 39 97 41
rect 63 37 97 39
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 35 27 43 29
rect 35 24 37 27
rect 47 25 49 37
rect 63 25 65 37
rect 75 25 77 37
rect 81 31 89 33
rect 81 29 83 31
rect 85 29 89 31
rect 81 27 89 29
rect 11 11 13 15
rect 23 11 25 15
rect 35 10 37 14
rect 47 11 49 15
rect 87 24 89 27
rect 87 10 89 14
rect 63 2 65 6
rect 75 2 77 6
<< ndif >>
rect 3 15 11 25
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 15 23 19
rect 25 24 30 25
rect 67 31 73 33
rect 67 29 69 31
rect 71 29 73 31
rect 67 25 73 29
rect 42 24 47 25
rect 25 15 35 24
rect 3 11 9 15
rect 27 14 35 15
rect 37 21 47 24
rect 37 19 41 21
rect 43 19 47 21
rect 37 15 47 19
rect 49 15 63 25
rect 37 14 45 15
rect 27 11 33 14
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 27 9 29 11
rect 31 9 33 11
rect 51 11 63 15
rect 27 7 33 9
rect 51 9 55 11
rect 57 9 63 11
rect 51 6 63 9
rect 65 6 75 25
rect 77 24 82 25
rect 77 14 87 24
rect 89 21 97 24
rect 89 19 93 21
rect 95 19 97 21
rect 89 14 97 19
rect 77 11 85 14
rect 77 9 81 11
rect 83 9 85 11
rect 77 6 85 9
<< pdif >>
rect 14 85 19 94
rect 7 81 19 85
rect 7 79 9 81
rect 11 79 19 81
rect 7 71 19 79
rect 7 69 9 71
rect 11 69 19 71
rect 7 61 19 69
rect 7 59 9 61
rect 11 59 19 61
rect 7 56 19 59
rect 21 56 27 94
rect 29 56 35 94
rect 37 56 43 94
rect 45 91 63 94
rect 45 89 49 91
rect 51 89 57 91
rect 59 89 63 91
rect 45 56 63 89
rect 7 55 13 56
rect 52 55 63 56
rect 65 81 75 94
rect 65 79 69 81
rect 71 79 75 81
rect 65 71 75 79
rect 65 69 69 71
rect 71 69 75 71
rect 65 61 75 69
rect 65 59 69 61
rect 71 59 75 61
rect 65 55 75 59
rect 77 91 85 94
rect 77 89 81 91
rect 83 89 85 91
rect 77 81 85 89
rect 77 79 81 81
rect 83 79 85 81
rect 77 76 85 79
rect 77 71 87 76
rect 77 69 81 71
rect 83 69 87 71
rect 77 61 87 69
rect 77 59 81 61
rect 83 59 87 61
rect 77 56 87 59
rect 89 71 97 76
rect 89 69 93 71
rect 95 69 97 71
rect 89 61 97 69
rect 89 59 93 61
rect 95 59 97 61
rect 89 56 97 59
rect 77 55 82 56
<< alu1 >>
rect -2 95 102 100
rect -2 93 93 95
rect 95 93 102 95
rect -2 91 102 93
rect -2 89 49 91
rect 51 89 57 91
rect 59 89 81 91
rect 83 89 102 91
rect -2 88 102 89
rect 8 81 12 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 71 12 79
rect 8 69 9 71
rect 11 69 12 71
rect 8 61 12 69
rect 8 59 9 61
rect 11 59 12 61
rect 8 22 12 59
rect 18 51 22 83
rect 18 49 19 51
rect 21 49 22 51
rect 18 27 22 49
rect 28 41 32 83
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 31 42 83
rect 38 29 39 31
rect 41 29 42 31
rect 38 27 42 29
rect 48 41 52 83
rect 48 39 49 41
rect 51 39 52 41
rect 48 27 52 39
rect 68 81 72 83
rect 68 79 69 81
rect 71 79 72 81
rect 68 71 72 79
rect 68 69 69 71
rect 71 69 72 71
rect 68 61 72 69
rect 68 59 69 61
rect 71 59 72 61
rect 68 31 72 59
rect 80 81 84 88
rect 80 79 81 81
rect 83 79 84 81
rect 80 71 84 79
rect 80 69 81 71
rect 83 69 84 71
rect 80 61 84 69
rect 80 59 81 61
rect 83 59 84 61
rect 80 57 84 59
rect 92 71 96 73
rect 92 69 93 71
rect 95 69 96 71
rect 92 61 96 69
rect 92 59 93 61
rect 95 59 96 61
rect 68 29 69 31
rect 71 29 72 31
rect 68 27 72 29
rect 78 51 87 52
rect 78 49 83 51
rect 85 49 87 51
rect 78 48 87 49
rect 78 32 82 48
rect 92 41 96 59
rect 92 39 93 41
rect 95 39 96 41
rect 78 31 87 32
rect 78 29 83 31
rect 85 29 87 31
rect 78 28 87 29
rect 78 22 82 28
rect 8 21 82 22
rect 8 19 17 21
rect 19 19 41 21
rect 43 19 82 21
rect 8 18 82 19
rect 92 21 96 39
rect 92 19 93 21
rect 95 19 96 21
rect 92 17 96 19
rect -2 11 102 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 55 11
rect 57 9 81 11
rect 83 9 102 11
rect -2 0 102 9
<< ntie >>
rect 91 95 97 97
rect 91 93 93 95
rect 95 93 97 95
rect 91 86 97 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 14 37 24
rect 47 15 49 25
rect 63 6 65 25
rect 75 6 77 25
rect 87 14 89 24
<< pmos >>
rect 19 56 21 94
rect 27 56 29 94
rect 35 56 37 94
rect 43 56 45 94
rect 63 55 65 94
rect 75 55 77 94
rect 87 56 89 76
<< polyct1 >>
rect 19 49 21 51
rect 29 39 31 41
rect 83 49 85 51
rect 49 39 51 41
rect 93 39 95 41
rect 39 29 41 31
rect 83 29 85 31
<< ndifct1 >>
rect 17 19 19 21
rect 69 29 71 31
rect 41 19 43 21
rect 5 9 7 11
rect 29 9 31 11
rect 55 9 57 11
rect 93 19 95 21
rect 81 9 83 11
<< ntiect1 >>
rect 93 93 95 95
<< pdifct1 >>
rect 9 79 11 81
rect 9 69 11 71
rect 9 59 11 61
rect 49 89 51 91
rect 57 89 59 91
rect 69 79 71 81
rect 69 69 71 71
rect 69 59 71 61
rect 81 89 83 91
rect 81 79 83 81
rect 81 69 83 71
rect 81 59 83 61
rect 93 69 95 71
rect 93 59 95 61
<< labels >>
rlabel alu1 20 55 20 55 6 i1
rlabel alu1 30 55 30 55 6 i0
rlabel alu1 40 55 40 55 6 i2
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 50 55 50 55 6 i3
rlabel alu1 70 55 70 55 6 nq
rlabel alu1 50 94 50 94 6 vdd
<< end >>
