magic
tech scmos
timestamp 1199203562
<< ab >>
rect 0 0 136 80
<< nwell >>
rect -5 36 141 88
<< pwell >>
rect -5 -8 141 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 66 70 68 74
rect 78 72 104 74
rect 78 63 80 72
rect 85 66 97 68
rect 85 63 87 66
rect 95 63 97 66
rect 102 63 104 72
rect 115 70 117 74
rect 125 61 127 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 37 21 39
rect 25 37 51 39
rect 55 37 61 39
rect 66 39 68 42
rect 78 39 80 42
rect 66 37 80 39
rect 85 39 87 42
rect 85 37 91 39
rect 95 38 97 42
rect 102 39 104 42
rect 115 39 117 42
rect 125 39 127 42
rect 9 35 15 37
rect 9 33 11 35
rect 13 33 15 35
rect 25 35 27 37
rect 29 35 31 37
rect 25 33 31 35
rect 55 35 57 37
rect 59 35 61 37
rect 55 33 61 35
rect 85 35 87 37
rect 89 35 91 37
rect 85 33 91 35
rect 101 37 107 39
rect 101 35 103 37
rect 105 35 107 37
rect 9 31 15 33
rect 19 31 31 33
rect 12 28 14 31
rect 19 28 21 31
rect 29 28 31 31
rect 36 28 38 33
rect 55 30 57 33
rect 12 8 14 16
rect 19 12 21 16
rect 29 12 31 16
rect 36 8 38 16
rect 12 6 38 8
rect 75 29 77 33
rect 85 29 87 33
rect 95 30 97 34
rect 101 33 107 35
rect 105 30 107 33
rect 115 37 127 39
rect 115 35 123 37
rect 125 35 127 37
rect 115 33 127 35
rect 115 30 117 33
rect 125 30 127 33
rect 55 10 57 15
rect 85 12 87 16
rect 95 14 97 17
rect 105 14 107 17
rect 95 12 107 14
rect 75 8 77 11
rect 115 8 117 17
rect 125 15 127 19
rect 75 6 117 8
<< ndif >>
rect 40 28 55 30
rect 3 16 12 28
rect 14 16 19 28
rect 21 21 29 28
rect 21 19 24 21
rect 26 19 29 21
rect 21 16 29 19
rect 31 16 36 28
rect 38 16 55 28
rect 3 11 10 16
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
rect 40 15 55 16
rect 57 28 64 30
rect 89 29 95 30
rect 57 26 60 28
rect 62 26 64 28
rect 57 24 64 26
rect 57 15 62 24
rect 70 23 75 29
rect 68 21 75 23
rect 68 19 70 21
rect 72 19 75 21
rect 68 17 75 19
rect 40 11 53 15
rect 40 9 42 11
rect 44 9 49 11
rect 51 9 53 11
rect 70 11 75 17
rect 77 27 85 29
rect 77 25 80 27
rect 82 25 85 27
rect 77 20 85 25
rect 77 18 80 20
rect 82 18 85 20
rect 77 16 85 18
rect 87 21 95 29
rect 87 19 90 21
rect 92 19 95 21
rect 87 17 95 19
rect 97 28 105 30
rect 97 26 100 28
rect 102 26 105 28
rect 97 21 105 26
rect 97 19 100 21
rect 102 19 105 21
rect 97 17 105 19
rect 107 21 115 30
rect 107 19 110 21
rect 112 19 115 21
rect 107 17 115 19
rect 117 28 125 30
rect 117 26 120 28
rect 122 26 125 28
rect 117 19 125 26
rect 127 24 134 30
rect 127 22 130 24
rect 132 22 134 24
rect 127 20 134 22
rect 127 19 132 20
rect 117 17 122 19
rect 87 16 93 17
rect 77 11 82 16
rect 40 7 53 9
<< pdif >>
rect 70 71 76 73
rect 70 70 72 71
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 61 29 70
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 46 39 70
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 61 49 70
rect 41 59 44 61
rect 46 59 49 61
rect 41 42 49 59
rect 51 46 59 70
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 42 66 70
rect 68 69 72 70
rect 74 69 76 71
rect 68 63 76 69
rect 106 71 113 73
rect 106 69 109 71
rect 111 70 113 71
rect 111 69 115 70
rect 106 63 115 69
rect 68 42 78 63
rect 80 42 85 63
rect 87 53 95 63
rect 87 51 90 53
rect 92 51 95 53
rect 87 46 95 51
rect 87 44 90 46
rect 92 44 95 46
rect 87 42 95 44
rect 97 42 102 63
rect 104 42 115 63
rect 117 61 122 70
rect 117 55 125 61
rect 117 53 120 55
rect 122 53 125 55
rect 117 47 125 53
rect 117 45 120 47
rect 122 45 125 47
rect 117 42 125 45
rect 127 59 134 61
rect 127 57 130 59
rect 132 57 134 59
rect 127 42 134 57
<< alu1 >>
rect -2 81 138 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 138 81
rect -2 71 138 79
rect -2 69 72 71
rect 74 69 109 71
rect 111 69 138 71
rect -2 68 138 69
rect 2 61 48 62
rect 2 59 4 61
rect 6 59 24 61
rect 26 59 44 61
rect 46 59 48 61
rect 2 58 48 59
rect 2 54 6 58
rect 2 52 4 54
rect 2 22 6 52
rect 74 38 78 47
rect 106 39 110 47
rect 49 37 91 38
rect 49 35 57 37
rect 59 35 87 37
rect 89 35 91 37
rect 49 34 91 35
rect 98 37 110 39
rect 98 35 103 37
rect 105 35 110 37
rect 98 33 110 35
rect 2 21 74 22
rect 2 19 24 21
rect 26 19 70 21
rect 72 19 74 21
rect 2 18 74 19
rect 106 25 110 33
rect 130 39 134 47
rect 122 37 134 39
rect 122 35 123 37
rect 125 35 134 37
rect 122 33 134 35
rect -2 11 138 12
rect -2 9 6 11
rect 8 9 42 11
rect 44 9 49 11
rect 51 9 138 11
rect -2 1 138 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 138 1
rect -2 -2 138 -1
<< ptie >>
rect 0 1 136 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 136 1
rect 0 -3 136 -1
<< ntie >>
rect 0 81 136 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 136 81
rect 0 77 136 79
<< nmos >>
rect 12 16 14 28
rect 19 16 21 28
rect 29 16 31 28
rect 36 16 38 28
rect 55 15 57 30
rect 75 11 77 29
rect 85 16 87 29
rect 95 17 97 30
rect 105 17 107 30
rect 115 17 117 30
rect 125 19 127 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 66 42 68 70
rect 78 42 80 63
rect 85 42 87 63
rect 95 42 97 63
rect 102 42 104 63
rect 115 42 117 70
rect 125 42 127 61
<< polyct0 >>
rect 11 33 13 35
rect 27 35 29 37
<< polyct1 >>
rect 57 35 59 37
rect 87 35 89 37
rect 103 35 105 37
rect 123 35 125 37
<< ndifct0 >>
rect 60 26 62 28
rect 80 25 82 27
rect 80 18 82 20
rect 90 19 92 21
rect 100 26 102 28
rect 100 19 102 21
rect 110 19 112 21
rect 120 26 122 28
rect 130 22 132 24
<< ndifct1 >>
rect 24 19 26 21
rect 6 9 8 11
rect 70 19 72 21
rect 42 9 44 11
rect 49 9 51 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
<< pdifct0 >>
rect 14 51 16 53
rect 14 44 16 46
rect 34 44 36 46
rect 54 44 56 46
rect 90 51 92 53
rect 90 44 92 46
rect 120 53 122 55
rect 120 45 122 47
rect 130 57 132 59
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
rect 24 59 26 61
rect 44 59 46 61
rect 72 69 74 71
rect 109 69 111 71
<< alu0 >>
rect 54 58 123 62
rect 6 50 7 58
rect 54 54 58 58
rect 119 55 123 58
rect 129 59 133 68
rect 129 57 130 59
rect 132 57 133 59
rect 129 55 133 57
rect 12 53 58 54
rect 12 51 14 53
rect 16 51 58 53
rect 12 50 58 51
rect 64 53 94 54
rect 64 51 90 53
rect 92 51 94 53
rect 64 50 94 51
rect 12 46 18 50
rect 12 44 14 46
rect 16 44 18 46
rect 12 43 18 44
rect 24 38 28 50
rect 32 46 38 47
rect 52 46 58 47
rect 64 46 68 50
rect 32 44 34 46
rect 36 44 54 46
rect 56 44 68 46
rect 32 42 68 44
rect 24 37 31 38
rect 10 35 14 37
rect 10 33 11 35
rect 13 33 14 35
rect 24 35 27 37
rect 29 35 31 37
rect 24 34 31 35
rect 10 30 14 33
rect 34 30 38 42
rect 89 46 94 50
rect 119 53 120 55
rect 122 53 123 55
rect 119 47 123 53
rect 89 44 90 46
rect 92 44 94 46
rect 89 42 94 44
rect 10 28 103 30
rect 10 26 60 28
rect 62 27 100 28
rect 62 26 80 27
rect 58 25 64 26
rect 78 25 80 26
rect 82 26 100 27
rect 102 26 103 28
rect 82 25 84 26
rect 78 20 84 25
rect 78 18 80 20
rect 82 18 84 20
rect 78 17 84 18
rect 88 21 94 22
rect 88 19 90 21
rect 92 19 94 21
rect 88 12 94 19
rect 99 21 103 26
rect 114 45 120 47
rect 122 45 123 47
rect 114 43 123 45
rect 114 29 118 43
rect 114 28 124 29
rect 114 26 120 28
rect 122 26 124 28
rect 114 25 124 26
rect 129 24 133 26
rect 129 22 130 24
rect 132 22 133 24
rect 99 19 100 21
rect 102 19 103 21
rect 99 17 103 19
rect 108 21 114 22
rect 108 19 110 21
rect 112 19 114 21
rect 108 12 114 19
rect 129 12 133 22
<< labels >>
rlabel alu0 12 31 12 31 6 an
rlabel alu0 15 48 15 48 6 bn
rlabel alu0 26 44 26 44 6 bn
rlabel alu0 55 44 55 44 6 an
rlabel alu0 50 44 50 44 6 an
rlabel alu0 81 23 81 23 6 an
rlabel alu0 56 28 56 28 6 an
rlabel alu0 101 23 101 23 6 an
rlabel alu0 91 48 91 48 6 an
rlabel alu0 79 52 79 52 6 an
rlabel alu0 119 27 119 27 6 bn
rlabel alu0 121 52 121 52 6 bn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 60 36 60 36 6 a2
rlabel alu1 52 36 52 36 6 a2
rlabel alu1 44 60 44 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 68 6 68 6 6 vss
rlabel alu1 68 20 68 20 6 z
rlabel alu1 68 36 68 36 6 a2
rlabel alu1 100 36 100 36 6 a1
rlabel alu1 84 36 84 36 6 a2
rlabel alu1 76 40 76 40 6 a2
rlabel alu1 68 74 68 74 6 vdd
rlabel polyct1 124 36 124 36 6 b
rlabel alu1 108 36 108 36 6 a1
rlabel alu1 132 40 132 40 6 b
<< end >>
