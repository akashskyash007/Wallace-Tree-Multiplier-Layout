magic
tech scmos
timestamp 1199202242
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 60 11 65
rect 9 39 11 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 30 11 33
rect 9 16 11 21
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 21 9 24
rect 11 25 22 30
rect 11 23 18 25
rect 20 23 22 25
rect 11 21 22 23
<< pdif >>
rect 13 61 20 63
rect 13 60 15 61
rect 4 55 9 60
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 59 15 60
rect 17 59 20 61
rect 11 42 20 59
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 68 26 79
rect 2 53 14 55
rect 2 51 4 53
rect 6 51 14 53
rect 2 49 14 51
rect 2 46 6 49
rect 2 44 4 46
rect 2 28 6 44
rect 10 37 22 39
rect 10 35 11 37
rect 13 35 22 37
rect 10 33 22 35
rect 2 26 4 28
rect 2 17 6 26
rect 10 25 14 33
rect -2 1 26 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 21 11 30
<< pmos >>
rect 9 42 11 60
<< polyct1 >>
rect 11 35 13 37
<< ndifct0 >>
rect 18 23 20 25
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct0 >>
rect 15 59 17 61
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 13 61 19 68
rect 13 59 15 61
rect 17 59 19 61
rect 13 58 19 59
rect 6 42 7 49
rect 6 24 7 30
rect 17 25 21 27
rect 17 23 18 25
rect 20 23 21 25
rect 17 12 21 23
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 32 12 32 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 36 20 36 6 a
<< end >>
