magic
tech scmos
timestamp 1199203072
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 38 70 40 74
rect 45 70 47 74
rect 10 61 12 65
rect 20 61 22 65
rect 10 38 12 46
rect 20 39 22 46
rect 38 40 40 43
rect 9 36 15 38
rect 9 34 11 36
rect 13 34 15 36
rect 9 32 15 34
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 34 38 40 40
rect 34 36 36 38
rect 38 36 40 38
rect 19 33 25 35
rect 29 34 40 36
rect 45 38 47 43
rect 45 36 54 38
rect 45 34 50 36
rect 52 34 54 36
rect 12 29 14 32
rect 19 29 21 33
rect 29 29 31 34
rect 45 32 54 34
rect 45 29 47 32
rect 12 7 14 12
rect 19 7 21 12
rect 29 7 31 12
rect 45 7 47 12
<< ndif >>
rect 7 22 12 29
rect 5 20 12 22
rect 5 18 7 20
rect 9 18 12 20
rect 5 16 12 18
rect 7 12 12 16
rect 14 12 19 29
rect 21 20 29 29
rect 21 18 24 20
rect 26 18 29 20
rect 21 12 29 18
rect 31 12 45 29
rect 47 22 52 29
rect 47 20 54 22
rect 47 18 50 20
rect 52 18 54 20
rect 47 16 54 18
rect 47 12 52 16
rect 33 11 43 12
rect 33 9 37 11
rect 39 9 43 11
rect 33 7 43 9
<< pdif >>
rect 24 68 38 70
rect 24 66 29 68
rect 31 66 38 68
rect 2 63 8 65
rect 2 61 4 63
rect 6 61 8 63
rect 24 61 38 66
rect 2 46 10 61
rect 12 59 20 61
rect 12 57 15 59
rect 17 57 20 59
rect 12 46 20 57
rect 22 46 38 61
rect 24 43 38 46
rect 40 43 45 70
rect 47 62 52 70
rect 47 60 54 62
rect 47 58 50 60
rect 52 58 54 60
rect 47 53 54 58
rect 47 51 50 53
rect 52 51 54 53
rect 47 49 54 51
rect 47 43 52 49
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 14 60 54 62
rect 14 59 50 60
rect 14 57 15 59
rect 17 58 50 59
rect 52 58 54 60
rect 17 57 18 58
rect 14 55 18 57
rect 2 50 18 55
rect 25 50 39 54
rect 2 21 6 50
rect 10 42 23 46
rect 33 42 39 50
rect 49 53 54 58
rect 49 51 50 53
rect 52 51 54 53
rect 49 49 54 51
rect 10 36 14 42
rect 35 38 39 42
rect 10 34 11 36
rect 13 34 14 36
rect 10 25 14 34
rect 18 37 31 38
rect 18 35 21 37
rect 23 35 31 37
rect 18 34 31 35
rect 35 36 36 38
rect 38 36 39 38
rect 35 34 39 36
rect 49 36 54 39
rect 49 34 50 36
rect 52 34 54 36
rect 18 25 22 34
rect 49 30 54 34
rect 41 25 54 30
rect 2 20 11 21
rect 2 18 7 20
rect 9 18 11 20
rect 2 17 11 18
rect -2 11 58 12
rect -2 9 37 11
rect 39 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 12 12 14 29
rect 19 12 21 29
rect 29 12 31 29
rect 45 12 47 29
<< pmos >>
rect 10 46 12 61
rect 20 46 22 61
rect 38 43 40 70
rect 45 43 47 70
<< polyct1 >>
rect 11 34 13 36
rect 21 35 23 37
rect 36 36 38 38
rect 50 34 52 36
<< ndifct0 >>
rect 24 18 26 20
rect 50 18 52 20
<< ndifct1 >>
rect 7 18 9 20
rect 37 9 39 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 29 66 31 68
rect 4 61 6 63
<< pdifct1 >>
rect 15 57 17 59
rect 50 58 52 60
rect 50 51 52 53
<< alu0 >>
rect 3 63 7 68
rect 27 66 29 68
rect 31 66 33 68
rect 27 65 33 66
rect 3 61 4 63
rect 6 61 7 63
rect 3 59 7 61
rect 22 20 54 21
rect 22 18 24 20
rect 26 18 50 20
rect 52 18 54 20
rect 22 17 54 18
<< labels >>
rlabel alu0 38 19 38 19 6 n1
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 32 12 32 6 c
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 44 20 44 6 c
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 36 28 36 6 b
rlabel alu1 28 52 28 52 6 a1
rlabel alu1 36 48 36 48 6 a1
rlabel alu1 36 60 36 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 52 32 52 32 6 a2
rlabel alu1 52 52 52 52 6 z
rlabel alu1 44 60 44 60 6 z
<< end >>
