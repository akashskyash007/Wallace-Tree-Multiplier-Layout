magic
tech scmos
timestamp 1199203128
<< ab >>
rect 0 0 104 80
<< nwell >>
rect -5 36 109 88
<< pwell >>
rect -5 -8 109 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 46 70 48 74
rect 53 70 55 74
rect 63 70 65 74
rect 70 70 72 74
rect 80 62 82 67
rect 87 62 89 67
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 21 39
rect 9 35 11 37
rect 13 35 21 37
rect 9 33 21 35
rect 25 37 31 39
rect 25 35 27 37
rect 29 35 31 37
rect 25 33 31 35
rect 36 33 38 42
rect 46 33 48 42
rect 53 39 55 42
rect 63 39 65 42
rect 70 39 72 42
rect 80 39 82 42
rect 53 37 65 39
rect 69 37 82 39
rect 87 39 89 42
rect 87 37 95 39
rect 55 35 57 37
rect 59 35 61 37
rect 55 33 61 35
rect 9 30 11 33
rect 19 30 21 33
rect 36 31 51 33
rect 39 28 41 31
rect 49 28 51 31
rect 59 28 61 33
rect 69 35 71 37
rect 73 35 75 37
rect 69 33 75 35
rect 87 35 91 37
rect 93 35 95 37
rect 87 33 95 35
rect 69 28 71 33
rect 79 31 95 33
rect 79 28 81 31
rect 91 28 93 31
rect 29 22 31 27
rect 59 12 61 16
rect 9 6 11 11
rect 19 8 21 11
rect 29 8 31 11
rect 19 6 31 8
rect 39 6 41 11
rect 49 8 51 11
rect 69 8 71 16
rect 49 6 71 8
rect 79 6 81 11
rect 91 6 93 11
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 11 9 17
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 11 19 26
rect 21 22 26 30
rect 34 22 39 28
rect 21 20 29 22
rect 21 18 24 20
rect 26 18 29 20
rect 21 11 29 18
rect 31 20 39 22
rect 31 18 34 20
rect 36 18 39 20
rect 31 11 39 18
rect 41 15 49 28
rect 41 13 44 15
rect 46 13 49 15
rect 41 11 49 13
rect 51 25 59 28
rect 51 23 54 25
rect 56 23 59 25
rect 51 16 59 23
rect 61 20 69 28
rect 61 18 64 20
rect 66 18 69 20
rect 61 16 69 18
rect 71 25 79 28
rect 71 23 74 25
rect 76 23 79 25
rect 71 16 79 23
rect 51 11 56 16
rect 74 11 79 16
rect 81 11 91 28
rect 93 22 98 28
rect 93 20 100 22
rect 93 18 96 20
rect 98 18 100 20
rect 93 16 100 18
rect 93 11 98 16
rect 83 9 85 11
rect 87 9 89 11
rect 83 7 89 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 60 19 70
rect 11 58 14 60
rect 16 58 19 60
rect 11 53 19 58
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 42 36 70
rect 38 60 46 70
rect 38 58 41 60
rect 43 58 46 60
rect 38 53 46 58
rect 38 51 41 53
rect 43 51 46 53
rect 38 42 46 51
rect 48 42 53 70
rect 55 68 63 70
rect 55 66 58 68
rect 60 66 63 68
rect 55 61 63 66
rect 55 59 58 61
rect 60 59 63 61
rect 55 42 63 59
rect 65 42 70 70
rect 72 62 77 70
rect 72 60 80 62
rect 72 58 75 60
rect 77 58 80 60
rect 72 53 80 58
rect 72 51 75 53
rect 77 51 80 53
rect 72 42 80 51
rect 82 42 87 62
rect 89 60 97 62
rect 89 58 92 60
rect 94 58 97 60
rect 89 53 97 58
rect 89 51 92 53
rect 94 51 97 53
rect 89 42 97 51
<< alu1 >>
rect -2 81 106 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 106 81
rect -2 68 106 79
rect 40 60 46 63
rect 40 58 41 60
rect 43 58 46 60
rect 73 60 79 63
rect 73 58 75 60
rect 77 58 79 60
rect 40 54 46 58
rect 73 54 79 58
rect 2 53 79 54
rect 2 51 14 53
rect 16 51 41 53
rect 43 51 75 53
rect 77 51 79 53
rect 2 50 79 51
rect 2 28 6 50
rect 10 42 23 46
rect 57 42 95 46
rect 10 37 14 42
rect 57 38 61 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 25 37 61 38
rect 25 35 27 37
rect 29 35 57 37
rect 59 35 61 37
rect 25 34 61 35
rect 65 37 85 38
rect 65 35 71 37
rect 73 35 85 37
rect 65 34 85 35
rect 89 37 95 42
rect 89 35 91 37
rect 93 35 95 37
rect 89 34 95 35
rect 81 30 85 34
rect 2 26 4 28
rect 2 21 6 26
rect 81 26 95 30
rect 2 19 4 21
rect 6 20 28 21
rect 6 19 24 20
rect 2 18 24 19
rect 26 18 28 20
rect 2 17 28 18
rect -2 11 106 12
rect -2 9 85 11
rect 87 9 106 11
rect -2 1 106 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 106 1
rect -2 -2 106 -1
<< ptie >>
rect 0 1 104 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 104 1
rect 0 -3 104 -1
<< ntie >>
rect 0 81 104 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 104 81
rect 0 77 104 79
<< nmos >>
rect 9 11 11 30
rect 19 11 21 30
rect 29 11 31 22
rect 39 11 41 28
rect 49 11 51 28
rect 59 16 61 28
rect 69 16 71 28
rect 79 11 81 28
rect 91 11 93 28
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 36 42 38 70
rect 46 42 48 70
rect 53 42 55 70
rect 63 42 65 70
rect 70 42 72 70
rect 80 42 82 62
rect 87 42 89 62
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 57 35 59 37
rect 71 35 73 37
rect 91 35 93 37
<< ndifct0 >>
rect 14 26 16 28
rect 34 18 36 20
rect 44 13 46 15
rect 54 23 56 25
rect 64 18 66 20
rect 74 23 76 25
rect 96 18 98 20
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
rect 24 18 26 20
rect 85 9 87 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 58 16 60
rect 24 66 26 68
rect 24 59 26 61
rect 58 66 60 68
rect 58 59 60 61
rect 92 58 94 60
rect 92 51 94 53
<< pdifct1 >>
rect 14 51 16 53
rect 41 58 43 60
rect 41 51 43 53
rect 75 58 77 60
rect 75 51 77 53
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 60 17 62
rect 13 58 14 60
rect 16 58 17 60
rect 22 61 28 66
rect 56 66 58 68
rect 60 66 62 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 56 61 62 66
rect 56 59 58 61
rect 60 59 62 61
rect 56 58 62 59
rect 13 54 17 58
rect 90 60 96 68
rect 90 58 92 60
rect 94 58 96 60
rect 90 53 96 58
rect 90 51 92 53
rect 94 51 96 53
rect 90 50 96 51
rect 6 21 8 29
rect 12 28 77 29
rect 12 26 14 28
rect 16 26 77 28
rect 12 25 77 26
rect 32 20 38 25
rect 53 23 54 25
rect 56 23 57 25
rect 53 21 57 23
rect 73 23 74 25
rect 76 23 77 25
rect 73 21 77 23
rect 32 18 34 20
rect 36 18 38 20
rect 32 17 38 18
rect 62 20 68 21
rect 62 18 64 20
rect 66 18 68 20
rect 43 15 47 17
rect 43 13 44 15
rect 46 13 47 15
rect 43 12 47 13
rect 62 12 68 18
rect 73 20 100 21
rect 73 18 96 20
rect 98 18 100 20
rect 73 17 100 18
<< labels >>
rlabel alu0 35 23 35 23 6 n1
rlabel alu0 44 27 44 27 6 n1
rlabel alu0 86 19 86 19 6 n1
rlabel alu1 4 32 4 32 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 44 20 44 6 b
rlabel alu1 36 36 36 36 6 a1
rlabel polyct1 28 36 28 36 6 a1
rlabel alu1 36 52 36 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 52 6 52 6 6 vss
rlabel alu1 44 36 44 36 6 a1
rlabel alu1 60 44 60 44 6 a1
rlabel alu1 52 36 52 36 6 a1
rlabel alu1 60 52 60 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 52 74 52 74 6 vdd
rlabel alu1 76 44 76 44 6 a1
rlabel alu1 76 36 76 36 6 a2
rlabel alu1 68 44 68 44 6 a1
rlabel alu1 68 36 68 36 6 a2
rlabel alu1 68 52 68 52 6 z
rlabel alu1 76 56 76 56 6 z
rlabel alu1 84 28 84 28 6 a2
rlabel alu1 92 28 92 28 6 a2
rlabel alu1 84 44 84 44 6 a1
rlabel alu1 92 40 92 40 6 a1
<< end >>
