magic
tech scmos
timestamp 1199202475
<< ab >>
rect 0 0 112 72
<< nwell >>
rect -5 32 117 77
<< pwell >>
rect -5 -5 117 32
<< poly >>
rect 9 68 94 70
rect 9 58 11 68
rect 19 58 21 63
rect 29 58 31 63
rect 39 58 41 68
rect 50 60 52 64
rect 63 60 65 64
rect 73 60 75 64
rect 83 60 85 64
rect 92 61 94 68
rect 92 59 103 61
rect 101 56 103 59
rect 9 33 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 17 33 31 35
rect 39 33 41 38
rect 50 35 52 40
rect 63 37 65 40
rect 73 37 75 40
rect 63 35 75 37
rect 83 37 85 40
rect 83 35 97 37
rect 48 33 54 35
rect 17 31 19 33
rect 21 31 31 33
rect 48 31 50 33
rect 52 31 54 33
rect 17 29 35 31
rect 33 26 35 29
rect 45 29 54 31
rect 63 34 69 35
rect 63 32 65 34
rect 67 32 69 34
rect 63 30 69 32
rect 91 33 93 35
rect 95 33 97 35
rect 91 31 97 33
rect 101 31 103 40
rect 45 26 47 29
rect 66 26 68 30
rect 76 29 87 31
rect 76 26 78 29
rect 85 27 87 29
rect 101 29 110 31
rect 101 27 106 29
rect 108 27 110 29
rect 85 25 110 27
rect 96 22 98 25
rect 96 7 98 12
rect 33 2 35 6
rect 45 2 47 6
rect 66 2 68 6
rect 76 2 78 6
<< ndif >>
rect 24 17 33 26
rect 24 15 27 17
rect 29 15 33 17
rect 24 10 33 15
rect 24 8 27 10
rect 29 8 33 10
rect 24 6 33 8
rect 35 17 45 26
rect 35 15 38 17
rect 40 15 45 17
rect 35 6 45 15
rect 47 24 54 26
rect 47 22 50 24
rect 52 22 54 24
rect 47 17 54 22
rect 47 15 50 17
rect 52 15 54 17
rect 47 13 54 15
rect 47 6 52 13
rect 58 10 66 26
rect 58 8 61 10
rect 63 8 66 10
rect 58 6 66 8
rect 68 24 76 26
rect 68 22 71 24
rect 73 22 76 24
rect 68 6 76 22
rect 78 19 83 26
rect 89 20 96 22
rect 78 17 85 19
rect 78 15 81 17
rect 83 15 85 17
rect 89 18 91 20
rect 93 18 96 20
rect 89 16 96 18
rect 78 13 85 15
rect 78 6 83 13
rect 91 12 96 16
rect 98 12 107 22
rect 100 7 107 12
rect 100 5 102 7
rect 104 5 107 7
rect 100 3 107 5
<< pdif >>
rect 43 58 50 60
rect 4 51 9 58
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 42 19 58
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 56 29 58
rect 21 54 24 56
rect 26 54 29 56
rect 21 38 29 54
rect 31 42 39 58
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 56 45 58
rect 47 56 50 58
rect 41 40 50 56
rect 52 44 63 60
rect 52 42 58 44
rect 60 42 63 44
rect 52 40 63 42
rect 65 58 73 60
rect 65 56 68 58
rect 70 56 73 58
rect 65 40 73 56
rect 75 44 83 60
rect 75 42 78 44
rect 80 42 83 44
rect 75 40 83 42
rect 85 46 90 60
rect 94 54 101 56
rect 94 52 96 54
rect 98 52 101 54
rect 94 50 101 52
rect 85 44 92 46
rect 85 42 88 44
rect 90 42 92 44
rect 85 40 92 42
rect 96 40 101 50
rect 103 54 110 56
rect 103 52 106 54
rect 108 52 110 54
rect 103 46 110 52
rect 103 44 106 46
rect 108 44 110 46
rect 103 40 110 44
rect 41 38 46 40
<< alu1 >>
rect -2 67 114 72
rect -2 65 98 67
rect 100 65 105 67
rect 107 65 114 67
rect -2 64 114 65
rect 42 58 49 59
rect 42 56 45 58
rect 47 56 49 58
rect 42 55 49 56
rect 42 50 46 55
rect 2 49 46 50
rect 2 47 4 49
rect 6 47 46 49
rect 2 46 46 47
rect 2 42 7 46
rect 2 40 4 42
rect 6 40 7 42
rect 2 37 7 40
rect 18 33 22 35
rect 18 31 19 33
rect 21 31 22 33
rect 18 19 22 31
rect 10 13 22 19
rect 42 26 46 46
rect 85 44 92 45
rect 85 42 88 44
rect 90 42 92 44
rect 85 41 92 42
rect 57 34 70 35
rect 57 32 65 34
rect 67 32 70 34
rect 57 29 70 32
rect 42 24 53 26
rect 42 22 50 24
rect 52 22 53 24
rect 57 22 63 29
rect 85 35 89 41
rect 42 21 53 22
rect 82 31 89 35
rect 48 18 53 21
rect 82 18 86 31
rect 48 17 86 18
rect 48 15 50 17
rect 52 15 81 17
rect 83 15 86 17
rect 105 29 110 35
rect 105 27 106 29
rect 108 27 110 29
rect 105 19 110 27
rect 48 14 86 15
rect 98 13 110 19
rect -2 7 114 8
rect -2 5 5 7
rect 7 5 102 7
rect 104 5 114 7
rect -2 0 114 5
<< ptie >>
rect 3 7 9 24
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 96 67 109 69
rect 96 65 98 67
rect 100 65 105 67
rect 107 65 109 67
rect 96 63 109 65
<< nmos >>
rect 33 6 35 26
rect 45 6 47 26
rect 66 6 68 26
rect 76 6 78 26
rect 96 12 98 22
<< pmos >>
rect 9 38 11 58
rect 19 38 21 58
rect 29 38 31 58
rect 39 38 41 58
rect 50 40 52 60
rect 63 40 65 60
rect 73 40 75 60
rect 83 40 85 60
rect 101 40 103 56
<< polyct0 >>
rect 50 31 52 33
rect 93 33 95 35
<< polyct1 >>
rect 19 31 21 33
rect 65 32 67 34
rect 106 27 108 29
<< ndifct0 >>
rect 27 15 29 17
rect 27 8 29 10
rect 38 15 40 17
rect 61 8 63 10
rect 71 22 73 24
rect 91 18 93 20
<< ndifct1 >>
rect 50 22 52 24
rect 50 15 52 17
rect 81 15 83 17
rect 102 5 104 7
<< ntiect1 >>
rect 98 65 100 67
rect 105 65 107 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 14 40 16 42
rect 24 54 26 56
rect 34 40 36 42
rect 58 42 60 44
rect 68 56 70 58
rect 78 42 80 44
rect 96 52 98 54
rect 106 52 108 54
rect 106 44 108 46
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 45 56 47 58
rect 88 42 90 44
<< alu0 >>
rect 22 56 28 64
rect 22 54 24 56
rect 26 54 28 56
rect 22 53 28 54
rect 66 58 72 64
rect 66 56 68 58
rect 70 56 72 58
rect 66 55 72 56
rect 95 54 99 56
rect 95 52 96 54
rect 98 52 99 54
rect 12 42 38 43
rect 12 40 14 42
rect 16 40 34 42
rect 36 40 38 42
rect 12 39 38 40
rect 26 17 30 19
rect 26 15 27 17
rect 29 15 30 17
rect 26 10 30 15
rect 34 18 38 39
rect 49 48 99 52
rect 49 33 53 48
rect 56 44 82 45
rect 56 42 58 44
rect 60 42 78 44
rect 80 42 82 44
rect 56 41 82 42
rect 49 31 50 33
rect 52 31 53 33
rect 49 29 53 31
rect 74 25 78 41
rect 95 37 99 48
rect 105 54 109 64
rect 105 52 106 54
rect 108 52 109 54
rect 105 46 109 52
rect 105 44 106 46
rect 108 44 109 46
rect 105 42 109 44
rect 69 24 78 25
rect 69 22 71 24
rect 73 22 78 24
rect 69 21 78 22
rect 92 35 99 37
rect 92 33 93 35
rect 95 33 99 35
rect 92 26 96 33
rect 34 17 42 18
rect 34 15 38 17
rect 40 15 42 17
rect 34 14 42 15
rect 90 22 96 26
rect 90 20 94 22
rect 90 18 91 20
rect 93 18 94 20
rect 90 16 94 18
rect 26 8 27 10
rect 29 8 30 10
rect 59 10 65 11
rect 59 8 61 10
rect 63 8 65 10
<< labels >>
rlabel alu0 51 40 51 40 6 sn
rlabel alu0 36 28 36 28 6 a0n
rlabel alu0 25 41 25 41 6 a0n
rlabel alu0 73 23 73 23 6 a1n
rlabel alu0 69 43 69 43 6 a1n
rlabel alu0 92 21 92 21 6 sn
rlabel alu0 94 29 94 29 6 sn
rlabel alu0 97 44 97 44 6 sn
rlabel alu1 12 16 12 16 6 a0
rlabel alu1 20 24 20 24 6 a0
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 40 44 40 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 56 4 56 4 6 vss
rlabel alu1 76 16 76 16 6 z
rlabel alu1 68 16 68 16 6 z
rlabel alu1 60 16 60 16 6 z
rlabel alu1 60 28 60 28 6 a1
rlabel alu1 68 32 68 32 6 a1
rlabel alu1 56 68 56 68 6 vdd
rlabel alu1 100 16 100 16 6 s
rlabel alu1 84 28 84 28 6 z
rlabel alu1 108 24 108 24 6 s
<< end >>
