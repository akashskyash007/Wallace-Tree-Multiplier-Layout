magic
tech scmos
timestamp 1199543794
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 11 94 13 98
rect 55 94 57 98
rect 67 94 69 98
rect 35 85 37 89
rect 43 85 45 89
rect 11 73 13 76
rect 11 71 19 73
rect 11 69 15 71
rect 17 69 19 71
rect 11 67 19 69
rect 35 53 37 56
rect 31 51 37 53
rect 43 53 45 56
rect 43 51 51 53
rect 3 41 9 43
rect 31 41 33 51
rect 43 49 47 51
rect 49 49 51 51
rect 43 47 51 49
rect 3 39 5 41
rect 7 39 33 41
rect 3 37 9 39
rect 11 31 19 33
rect 11 29 15 31
rect 17 29 19 31
rect 11 27 19 29
rect 11 24 13 27
rect 31 25 33 39
rect 37 41 43 43
rect 55 41 57 55
rect 67 41 69 55
rect 37 39 39 41
rect 41 39 69 41
rect 37 37 43 39
rect 43 31 51 33
rect 43 29 47 31
rect 49 29 51 31
rect 43 27 51 29
rect 43 24 45 27
rect 55 25 57 39
rect 67 25 69 39
rect 11 10 13 14
rect 31 11 33 15
rect 43 10 45 14
rect 55 2 57 6
rect 67 2 69 6
<< ndif >>
rect 15 24 31 25
rect 3 21 11 24
rect 3 19 5 21
rect 7 19 11 21
rect 3 14 11 19
rect 13 15 31 24
rect 33 24 38 25
rect 50 24 55 25
rect 33 21 43 24
rect 33 19 37 21
rect 39 19 43 21
rect 33 15 43 19
rect 13 14 29 15
rect 15 11 29 14
rect 35 14 43 15
rect 45 14 55 24
rect 15 9 17 11
rect 19 9 25 11
rect 27 9 29 11
rect 47 11 55 14
rect 15 7 29 9
rect 47 9 49 11
rect 51 9 55 11
rect 47 6 55 9
rect 57 21 67 25
rect 57 19 61 21
rect 63 19 67 21
rect 57 6 67 19
rect 69 21 77 25
rect 69 19 73 21
rect 75 19 77 21
rect 69 11 77 19
rect 69 9 73 11
rect 75 9 77 11
rect 69 6 77 9
<< pdif >>
rect 3 81 11 94
rect 3 79 5 81
rect 7 79 11 81
rect 3 76 11 79
rect 13 91 21 94
rect 47 91 55 94
rect 13 89 17 91
rect 19 89 21 91
rect 47 89 49 91
rect 51 89 55 91
rect 13 76 21 89
rect 47 85 55 89
rect 27 81 35 85
rect 27 79 29 81
rect 31 79 35 81
rect 27 71 35 79
rect 27 69 29 71
rect 31 69 35 71
rect 27 61 35 69
rect 27 59 29 61
rect 31 59 35 61
rect 27 56 35 59
rect 37 56 43 85
rect 45 56 55 85
rect 50 55 55 56
rect 57 81 67 94
rect 57 79 61 81
rect 63 79 67 81
rect 57 71 67 79
rect 57 69 61 71
rect 63 69 67 71
rect 57 61 67 69
rect 57 59 61 61
rect 63 59 67 61
rect 57 55 67 59
rect 69 91 77 94
rect 69 89 73 91
rect 75 89 77 91
rect 69 81 77 89
rect 69 79 73 81
rect 75 79 77 81
rect 69 71 77 79
rect 69 69 73 71
rect 75 69 77 71
rect 69 61 77 69
rect 69 59 73 61
rect 75 59 77 61
rect 69 55 77 59
<< alu1 >>
rect -2 95 82 100
rect -2 93 29 95
rect 31 93 37 95
rect 39 93 82 95
rect -2 91 82 93
rect -2 89 17 91
rect 19 89 49 91
rect 51 89 73 91
rect 75 89 82 91
rect -2 88 82 89
rect 4 81 8 83
rect 4 79 5 81
rect 7 79 8 81
rect 4 41 8 79
rect 18 72 22 83
rect 13 71 22 72
rect 13 69 15 71
rect 17 69 22 71
rect 13 68 22 69
rect 4 39 5 41
rect 7 39 8 41
rect 4 21 8 39
rect 18 32 22 68
rect 28 81 32 83
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 60 32 61
rect 31 59 40 60
rect 28 56 40 59
rect 13 31 22 32
rect 13 29 15 31
rect 17 29 22 31
rect 13 28 22 29
rect 4 19 5 21
rect 7 19 8 21
rect 4 17 8 19
rect 18 17 22 28
rect 36 42 40 56
rect 48 52 52 83
rect 45 51 52 52
rect 45 49 47 51
rect 49 49 52 51
rect 45 48 52 49
rect 36 41 43 42
rect 36 39 39 41
rect 41 39 43 41
rect 36 38 43 39
rect 36 21 40 38
rect 48 32 52 48
rect 45 31 52 32
rect 45 29 47 31
rect 49 29 52 31
rect 45 28 52 29
rect 36 19 37 21
rect 39 19 40 21
rect 36 17 40 19
rect 48 17 52 28
rect 58 82 62 83
rect 58 81 65 82
rect 58 79 61 81
rect 63 79 65 81
rect 58 78 65 79
rect 72 81 76 88
rect 72 79 73 81
rect 75 79 76 81
rect 58 72 62 78
rect 58 71 65 72
rect 58 69 61 71
rect 63 69 65 71
rect 58 68 65 69
rect 72 71 76 79
rect 72 69 73 71
rect 75 69 76 71
rect 58 62 62 68
rect 58 61 65 62
rect 58 59 61 61
rect 63 59 65 61
rect 58 58 65 59
rect 72 61 76 69
rect 72 59 73 61
rect 75 59 76 61
rect 58 22 62 58
rect 72 57 76 59
rect 58 21 65 22
rect 58 19 61 21
rect 63 19 65 21
rect 58 18 65 19
rect 72 21 76 23
rect 72 19 73 21
rect 75 19 76 21
rect 58 17 62 18
rect 72 12 76 19
rect -2 11 82 12
rect -2 9 17 11
rect 19 9 25 11
rect 27 9 49 11
rect 51 9 73 11
rect 75 9 82 11
rect -2 0 82 9
<< ntie >>
rect 27 95 41 97
rect 27 93 29 95
rect 31 93 37 95
rect 39 93 41 95
rect 27 91 41 93
<< nmos >>
rect 11 14 13 24
rect 31 15 33 25
rect 43 14 45 24
rect 55 6 57 25
rect 67 6 69 25
<< pmos >>
rect 11 76 13 94
rect 35 56 37 85
rect 43 56 45 85
rect 55 55 57 94
rect 67 55 69 94
<< polyct1 >>
rect 15 69 17 71
rect 47 49 49 51
rect 5 39 7 41
rect 15 29 17 31
rect 39 39 41 41
rect 47 29 49 31
<< ndifct1 >>
rect 5 19 7 21
rect 37 19 39 21
rect 17 9 19 11
rect 25 9 27 11
rect 49 9 51 11
rect 61 19 63 21
rect 73 19 75 21
rect 73 9 75 11
<< ntiect1 >>
rect 29 93 31 95
rect 37 93 39 95
<< pdifct1 >>
rect 5 79 7 81
rect 17 89 19 91
rect 49 89 51 91
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
rect 61 79 63 81
rect 61 69 63 71
rect 61 59 63 61
rect 73 89 75 91
rect 73 79 75 81
rect 73 69 75 71
rect 73 59 75 61
<< labels >>
rlabel alu1 20 50 20 50 6 i0
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 50 50 50 50 6 i1
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 60 50 60 50 6 q
<< end >>
