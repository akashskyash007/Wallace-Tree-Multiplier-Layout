magic
tech scmos
timestamp 1199543486
<< ab >>
rect 0 0 120 100
<< nwell >>
rect -2 48 122 104
<< pwell >>
rect -2 -4 122 48
<< poly >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 79 95 81 98
rect 91 95 93 98
rect 103 95 105 98
rect 11 53 13 55
rect 23 53 25 55
rect 35 53 37 55
rect 47 53 49 55
rect 79 53 81 55
rect 91 53 93 55
rect 11 51 19 53
rect 23 51 29 53
rect 35 51 43 53
rect 17 43 19 51
rect 27 43 29 51
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 77 51 83 53
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 87 51 93 53
rect 87 49 89 51
rect 91 49 93 51
rect 87 47 93 49
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 17 29 19 37
rect 27 29 29 37
rect 37 29 39 47
rect 47 29 49 47
rect 15 27 19 29
rect 23 27 29 29
rect 35 27 39 29
rect 43 27 49 29
rect 79 29 81 47
rect 79 27 85 29
rect 15 25 17 27
rect 23 25 25 27
rect 35 25 37 27
rect 43 25 45 27
rect 83 25 85 27
rect 91 25 93 47
rect 103 43 105 55
rect 97 41 105 43
rect 97 39 99 41
rect 101 39 105 41
rect 97 37 105 39
rect 103 25 105 37
rect 15 2 17 5
rect 23 2 25 5
rect 35 2 37 5
rect 43 2 45 5
rect 83 2 85 5
rect 91 2 93 5
rect 103 2 105 5
<< ndif >>
rect 7 11 15 25
rect 7 9 9 11
rect 11 9 15 11
rect 7 5 15 9
rect 17 5 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 5 35 19
rect 37 5 43 25
rect 45 11 53 25
rect 75 21 83 25
rect 75 19 77 21
rect 79 19 83 21
rect 45 9 49 11
rect 51 9 53 11
rect 45 5 53 9
rect 75 5 83 19
rect 85 5 91 25
rect 93 11 103 25
rect 93 9 97 11
rect 99 9 103 11
rect 93 5 103 9
rect 105 21 113 25
rect 105 19 109 21
rect 111 19 113 21
rect 105 5 113 19
<< pdif >>
rect 3 81 11 95
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 71 23 95
rect 13 69 17 71
rect 19 69 23 71
rect 13 55 23 69
rect 25 81 35 95
rect 25 79 29 81
rect 31 79 35 81
rect 25 55 35 79
rect 37 71 47 95
rect 37 69 41 71
rect 43 69 47 71
rect 37 55 47 69
rect 49 81 57 95
rect 49 79 53 81
rect 55 79 57 81
rect 49 55 57 79
rect 71 91 79 95
rect 71 89 73 91
rect 75 89 79 91
rect 71 81 79 89
rect 71 79 73 81
rect 75 79 79 81
rect 71 55 79 79
rect 81 81 91 95
rect 81 79 85 81
rect 87 79 91 81
rect 81 55 91 79
rect 93 91 103 95
rect 93 89 97 91
rect 99 89 103 91
rect 93 81 103 89
rect 93 79 97 81
rect 99 79 103 81
rect 93 71 103 79
rect 93 69 97 71
rect 99 69 103 71
rect 93 55 103 69
rect 105 81 113 95
rect 105 79 109 81
rect 111 79 113 81
rect 105 71 113 79
rect 105 69 109 71
rect 111 69 113 71
rect 105 61 113 69
rect 105 59 109 61
rect 111 59 113 61
rect 105 55 113 59
<< alu1 >>
rect -2 91 122 100
rect -2 89 73 91
rect 75 89 97 91
rect 99 89 122 91
rect -2 88 122 89
rect 4 81 8 82
rect 28 81 32 82
rect 52 81 56 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 53 81
rect 55 79 56 81
rect 4 78 8 79
rect 28 78 32 79
rect 52 78 56 79
rect 72 81 76 88
rect 72 79 73 81
rect 75 79 76 81
rect 72 78 76 79
rect 84 81 88 82
rect 84 79 85 81
rect 87 79 88 81
rect 84 78 88 79
rect 96 81 100 88
rect 96 79 97 81
rect 99 79 100 81
rect 16 71 20 72
rect 16 70 17 71
rect 9 69 17 70
rect 19 69 20 71
rect 9 68 20 69
rect 9 21 11 68
rect 18 41 22 62
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 28 41 32 72
rect 40 71 44 72
rect 85 71 87 78
rect 40 69 41 71
rect 43 69 87 71
rect 96 71 100 79
rect 96 69 97 71
rect 99 69 100 71
rect 40 68 44 69
rect 96 68 100 69
rect 108 81 112 82
rect 108 79 109 81
rect 111 79 112 81
rect 108 71 112 79
rect 108 69 109 71
rect 111 69 112 71
rect 28 39 29 41
rect 31 39 32 41
rect 28 28 32 39
rect 38 51 42 62
rect 38 49 39 51
rect 41 49 42 51
rect 38 28 42 49
rect 48 51 52 62
rect 48 49 49 51
rect 51 49 52 51
rect 48 28 52 49
rect 78 51 82 62
rect 78 49 79 51
rect 81 49 82 51
rect 78 28 82 49
rect 88 51 92 62
rect 88 49 89 51
rect 91 49 92 51
rect 88 28 92 49
rect 108 61 112 69
rect 108 59 109 61
rect 111 59 112 61
rect 98 41 102 42
rect 98 39 99 41
rect 101 39 102 41
rect 98 38 102 39
rect 28 21 32 22
rect 76 21 80 22
rect 99 21 101 38
rect 9 19 29 21
rect 31 19 77 21
rect 79 19 101 21
rect 108 21 112 59
rect 108 19 109 21
rect 111 19 112 21
rect 28 18 32 19
rect 76 18 80 19
rect 108 18 112 19
rect -2 11 122 12
rect -2 9 9 11
rect 11 9 49 11
rect 51 9 97 11
rect 99 9 122 11
rect -2 7 63 9
rect 65 7 122 9
rect -2 0 122 7
<< ptie >>
rect 61 9 67 17
rect 61 7 63 9
rect 65 7 67 9
rect 61 5 67 7
<< nmos >>
rect 15 5 17 25
rect 23 5 25 25
rect 35 5 37 25
rect 43 5 45 25
rect 83 5 85 25
rect 91 5 93 25
rect 103 5 105 25
<< pmos >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 79 55 81 95
rect 91 55 93 95
rect 103 55 105 95
<< polyct1 >>
rect 39 49 41 51
rect 49 49 51 51
rect 79 49 81 51
rect 89 49 91 51
rect 19 39 21 41
rect 29 39 31 41
rect 99 39 101 41
<< ndifct1 >>
rect 9 9 11 11
rect 29 19 31 21
rect 77 19 79 21
rect 49 9 51 11
rect 97 9 99 11
rect 109 19 111 21
<< ptiect1 >>
rect 63 7 65 9
<< pdifct1 >>
rect 5 79 7 81
rect 17 69 19 71
rect 29 79 31 81
rect 41 69 43 71
rect 53 79 55 81
rect 73 89 75 91
rect 73 79 75 81
rect 85 79 87 81
rect 97 89 99 91
rect 97 79 99 81
rect 97 69 99 71
rect 109 79 111 81
rect 109 69 111 71
rect 109 59 111 61
<< labels >>
rlabel alu1 40 45 40 45 6 i3
rlabel alu1 20 45 20 45 6 i5
rlabel alu1 30 50 30 50 6 i4
rlabel alu1 60 6 60 6 6 vss
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 60 94 60 94 6 vdd
rlabel alu1 80 45 80 45 6 i1
rlabel alu1 90 45 90 45 6 i0
rlabel alu1 110 50 110 50 6 q
<< end >>
