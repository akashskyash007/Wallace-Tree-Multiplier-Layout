magic
tech scmos
timestamp 1199980696
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -8 40 72 97
<< pwell >>
rect -8 -9 72 40
<< poly >>
rect 5 84 14 86
rect 5 82 7 84
rect 9 82 14 84
rect 5 80 14 82
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 42 11 48
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 2 32 17 38
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
<< ndif >>
rect 2 11 9 29
rect 11 23 21 29
rect 11 21 15 23
rect 17 21 21 23
rect 11 16 21 21
rect 11 14 15 16
rect 17 14 21 16
rect 11 11 21 14
rect 23 16 30 29
rect 23 14 26 16
rect 28 14 30 16
rect 23 11 30 14
rect 34 24 41 29
rect 34 22 36 24
rect 38 22 41 24
rect 34 11 41 22
rect 43 16 53 29
rect 43 14 47 16
rect 49 14 53 16
rect 43 11 53 14
rect 55 26 62 29
rect 55 24 58 26
rect 60 24 62 26
rect 55 18 62 24
rect 55 16 58 18
rect 60 16 62 18
rect 55 11 62 16
<< pdif >>
rect 2 51 9 77
rect 11 74 21 77
rect 11 72 15 74
rect 17 72 21 74
rect 11 67 21 72
rect 11 65 15 67
rect 17 65 21 67
rect 11 51 21 65
rect 23 74 30 77
rect 23 72 26 74
rect 28 72 30 74
rect 23 66 30 72
rect 23 64 26 66
rect 28 64 30 66
rect 23 51 30 64
rect 34 74 41 77
rect 34 72 36 74
rect 38 72 41 74
rect 34 66 41 72
rect 34 64 36 66
rect 38 64 41 66
rect 34 51 41 64
rect 43 65 53 77
rect 43 63 47 65
rect 49 63 53 65
rect 43 57 53 63
rect 43 55 47 57
rect 49 55 53 57
rect 43 51 53 55
rect 55 74 62 77
rect 55 72 58 74
rect 60 72 62 74
rect 55 67 62 72
rect 55 65 58 67
rect 60 65 62 67
rect 55 51 62 65
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect 62 85 66 90
rect -2 83 -1 85
rect 1 84 31 85
rect 1 83 7 84
rect -2 82 7 83
rect 9 82 15 84
rect 17 83 31 84
rect 33 83 34 85
rect 17 82 34 83
rect -2 81 34 82
rect 57 83 63 85
rect 65 83 66 85
rect 57 81 66 83
rect 14 74 18 81
rect 14 72 15 74
rect 17 72 18 74
rect 14 67 18 72
rect 57 74 61 81
rect 57 72 58 74
rect 60 72 61 74
rect 57 67 61 72
rect 14 65 15 67
rect 17 65 18 67
rect 14 63 18 65
rect 46 65 50 67
rect 46 63 47 65
rect 49 63 50 65
rect 57 65 58 67
rect 60 65 61 67
rect 57 63 61 65
rect 22 46 26 59
rect 46 57 50 63
rect 46 55 47 57
rect 49 55 50 57
rect 22 44 23 46
rect 25 44 26 46
rect 22 36 26 44
rect 22 34 23 36
rect 25 34 26 36
rect 22 32 26 34
rect 38 46 42 51
rect 38 44 39 46
rect 41 44 42 46
rect 38 36 42 44
rect 38 34 39 36
rect 41 34 42 36
rect 38 29 42 34
rect 46 28 50 55
rect 54 46 58 59
rect 54 44 55 46
rect 57 44 58 46
rect 54 36 58 44
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 46 26 61 28
rect 14 24 40 25
rect 46 24 58 26
rect 60 24 61 26
rect 14 23 36 24
rect 14 21 15 23
rect 17 22 36 23
rect 38 22 40 24
rect 17 21 40 22
rect 14 16 18 21
rect 54 18 61 24
rect 14 14 15 16
rect 17 14 18 16
rect 14 7 18 14
rect 54 16 58 18
rect 60 16 61 18
rect 54 13 61 16
rect -2 6 34 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 4 15 6
rect 17 5 34 6
rect 17 4 31 5
rect 1 3 31 4
rect 33 3 34 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 5 66 7
rect 62 3 63 5
rect 65 3 66 5
rect 62 -2 66 3
<< alu2 >>
rect -2 85 66 90
rect -2 83 -1 85
rect 1 84 31 85
rect 1 83 15 84
rect -2 82 15 83
rect 17 83 31 84
rect 33 83 63 85
rect 65 83 66 85
rect 17 82 66 83
rect -2 80 66 82
rect -2 6 66 8
rect -2 5 15 6
rect -2 3 -1 5
rect 1 4 15 5
rect 17 5 66 6
rect 17 4 31 5
rect 1 3 31 4
rect 33 3 63 5
rect 65 3 66 5
rect -2 -2 66 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polyct1 >>
rect 7 82 9 84
rect 23 44 25 46
rect 39 44 41 46
rect 55 44 57 46
rect 23 34 25 36
rect 39 34 41 36
rect 55 34 57 36
rect 7 4 9 6
<< ndifct0 >>
rect 26 14 28 16
rect 47 14 49 16
<< ndifct1 >>
rect 15 21 17 23
rect 15 14 17 16
rect 36 22 38 24
rect 58 24 60 26
rect 58 16 60 18
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< pdifct0 >>
rect 26 72 28 74
rect 26 64 28 66
rect 36 72 38 74
rect 36 64 38 66
<< pdifct1 >>
rect 15 72 17 74
rect 15 65 17 67
rect 47 63 49 65
rect 47 55 49 57
rect 58 72 60 74
rect 58 65 60 67
<< alu0 >>
rect 24 74 40 75
rect 24 72 26 74
rect 28 72 36 74
rect 38 72 40 74
rect 24 71 40 72
rect 24 66 40 67
rect 24 64 26 66
rect 28 64 36 66
rect 38 64 40 66
rect 24 63 40 64
rect 24 16 51 17
rect 24 14 26 16
rect 28 14 47 16
rect 49 14 51 16
rect 24 13 51 14
<< via1 >>
rect -1 83 1 85
rect 15 82 17 84
rect 31 83 33 85
rect 63 83 65 85
rect -1 3 1 5
rect 15 4 17 6
rect 31 3 33 5
rect 63 3 65 5
<< labels >>
rlabel alu1 24 48 24 48 6 a1
rlabel alu1 40 40 40 40 6 a2
rlabel alu1 56 20 56 20 6 z
rlabel alu1 56 48 56 48 6 b
rlabel alu1 48 48 48 48 6 z
rlabel via1 32 4 32 4 6 vss
rlabel via1 32 84 32 84 6 vdd
<< end >>
