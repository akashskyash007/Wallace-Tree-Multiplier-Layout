magic
tech scmos
timestamp 1199203387
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< labels >>
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 74 28 74 6 vdd
<< end >>
