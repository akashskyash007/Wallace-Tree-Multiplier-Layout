magic
tech scmos
timestamp 1199203131
<< ab >>
rect 0 0 152 72
<< nwell >>
rect -5 32 157 77
<< pwell >>
rect -5 -5 157 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 46 66 48 70
rect 56 66 58 70
rect 63 66 65 70
rect 73 66 75 70
rect 80 66 82 70
rect 90 66 92 70
rect 97 66 99 70
rect 107 66 109 70
rect 114 66 116 70
rect 124 58 126 63
rect 131 58 133 63
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 46 35 48 38
rect 56 35 58 38
rect 9 33 31 35
rect 9 26 11 33
rect 18 31 20 33
rect 22 31 27 33
rect 29 31 31 33
rect 18 29 31 31
rect 36 33 42 35
rect 46 33 58 35
rect 63 35 65 38
rect 73 35 75 38
rect 63 33 75 35
rect 80 35 82 38
rect 90 35 92 38
rect 80 33 92 35
rect 97 35 99 38
rect 107 35 109 38
rect 114 35 116 38
rect 124 35 126 38
rect 131 35 133 38
rect 97 33 109 35
rect 36 31 38 33
rect 40 31 42 33
rect 36 29 42 31
rect 19 26 21 29
rect 29 26 31 29
rect 40 20 42 25
rect 50 24 52 33
rect 66 31 68 33
rect 70 31 72 33
rect 66 29 72 31
rect 80 31 82 33
rect 84 31 86 33
rect 80 29 86 31
rect 97 31 105 33
rect 107 31 109 33
rect 97 29 109 31
rect 113 33 126 35
rect 130 33 136 35
rect 113 31 115 33
rect 117 31 119 33
rect 113 29 119 31
rect 130 31 132 33
rect 134 31 136 33
rect 130 29 142 31
rect 60 24 62 29
rect 70 26 72 29
rect 83 26 85 29
rect 93 27 105 29
rect 70 8 72 12
rect 93 24 95 27
rect 103 24 105 27
rect 113 26 115 29
rect 130 26 132 29
rect 140 26 142 29
rect 9 2 11 7
rect 19 2 21 7
rect 29 4 31 7
rect 40 4 42 7
rect 29 2 42 4
rect 50 4 52 7
rect 60 4 62 7
rect 83 4 85 10
rect 130 11 132 16
rect 140 11 142 16
rect 50 2 85 4
rect 93 2 95 6
rect 103 2 105 6
rect 113 2 115 6
<< ndif >>
rect 4 18 9 26
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 4 7 9 12
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 7 19 22
rect 21 16 29 26
rect 21 14 24 16
rect 26 14 29 16
rect 21 7 29 14
rect 31 24 38 26
rect 31 22 34 24
rect 36 22 38 24
rect 31 20 38 22
rect 65 24 70 26
rect 45 20 50 24
rect 31 7 40 20
rect 42 18 50 20
rect 42 16 45 18
rect 47 16 50 18
rect 42 7 50 16
rect 52 11 60 24
rect 52 9 55 11
rect 57 9 60 11
rect 52 7 60 9
rect 62 21 70 24
rect 62 19 65 21
rect 67 19 70 21
rect 62 12 70 19
rect 72 16 83 26
rect 72 14 77 16
rect 79 14 83 16
rect 72 12 83 14
rect 62 7 67 12
rect 78 10 83 12
rect 85 24 90 26
rect 108 24 113 26
rect 85 21 93 24
rect 85 19 88 21
rect 90 19 93 21
rect 85 10 93 19
rect 88 6 93 10
rect 95 10 103 24
rect 95 8 98 10
rect 100 8 103 10
rect 95 6 103 8
rect 105 17 113 24
rect 105 15 108 17
rect 110 15 113 17
rect 105 6 113 15
rect 115 16 130 26
rect 132 21 140 26
rect 132 19 135 21
rect 137 19 140 21
rect 132 16 140 19
rect 142 20 149 26
rect 142 18 145 20
rect 147 18 149 20
rect 142 16 149 18
rect 115 10 128 16
rect 115 8 122 10
rect 124 8 128 10
rect 115 6 128 8
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 19 66
rect 11 62 14 64
rect 16 62 19 64
rect 11 57 19 62
rect 11 55 14 57
rect 16 55 19 57
rect 11 38 19 55
rect 21 56 29 66
rect 21 54 24 56
rect 26 54 29 56
rect 21 49 29 54
rect 21 47 24 49
rect 26 47 29 49
rect 21 38 29 47
rect 31 64 39 66
rect 31 62 34 64
rect 36 62 39 64
rect 31 57 39 62
rect 31 55 34 57
rect 36 55 39 57
rect 31 38 39 55
rect 41 38 46 66
rect 48 56 56 66
rect 48 54 51 56
rect 53 54 56 56
rect 48 49 56 54
rect 48 47 51 49
rect 53 47 56 49
rect 48 38 56 47
rect 58 38 63 66
rect 65 64 73 66
rect 65 62 68 64
rect 70 62 73 64
rect 65 57 73 62
rect 65 55 68 57
rect 70 55 73 57
rect 65 38 73 55
rect 75 38 80 66
rect 82 56 90 66
rect 82 54 85 56
rect 87 54 90 56
rect 82 49 90 54
rect 82 47 85 49
rect 87 47 90 49
rect 82 38 90 47
rect 92 38 97 66
rect 99 64 107 66
rect 99 62 102 64
rect 104 62 107 64
rect 99 57 107 62
rect 99 55 102 57
rect 104 55 107 57
rect 99 38 107 55
rect 109 38 114 66
rect 116 58 121 66
rect 116 56 124 58
rect 116 54 119 56
rect 121 54 124 56
rect 116 49 124 54
rect 116 47 119 49
rect 121 47 124 49
rect 116 38 124 47
rect 126 38 131 58
rect 133 56 140 58
rect 133 54 136 56
rect 138 54 140 56
rect 133 49 140 54
rect 133 47 136 49
rect 138 47 140 49
rect 133 38 140 47
<< alu1 >>
rect -2 67 154 72
rect -2 65 143 67
rect 145 65 154 67
rect -2 64 154 65
rect 50 56 54 59
rect 50 54 51 56
rect 53 54 54 56
rect 82 56 88 59
rect 82 54 85 56
rect 87 54 88 56
rect 50 50 54 54
rect 82 50 88 54
rect 2 49 127 50
rect 2 47 4 49
rect 6 47 24 49
rect 26 47 51 49
rect 53 47 85 49
rect 87 47 119 49
rect 121 47 127 49
rect 2 46 127 47
rect 2 42 6 46
rect 2 40 4 42
rect 2 26 6 40
rect 25 38 39 42
rect 68 38 135 42
rect 25 34 31 38
rect 68 34 72 38
rect 17 33 31 34
rect 17 31 20 33
rect 22 31 27 33
rect 29 31 31 33
rect 17 30 31 31
rect 36 33 72 34
rect 36 31 38 33
rect 40 31 68 33
rect 70 31 72 33
rect 36 30 72 31
rect 80 33 99 34
rect 80 31 82 33
rect 84 31 99 33
rect 80 30 99 31
rect 113 33 119 34
rect 113 31 115 33
rect 117 31 119 33
rect 95 26 99 30
rect 113 26 119 31
rect 130 33 135 38
rect 130 31 132 33
rect 134 31 135 33
rect 130 29 135 31
rect 2 24 39 26
rect 2 22 14 24
rect 16 22 34 24
rect 36 22 39 24
rect 2 21 39 22
rect 95 22 119 26
rect -2 7 154 8
rect -2 5 134 7
rect 136 5 145 7
rect 147 5 154 7
rect -2 0 154 5
<< ptie >>
rect 132 7 149 9
rect 132 5 134 7
rect 136 5 145 7
rect 147 5 149 7
rect 132 3 149 5
<< ntie >>
rect 139 67 149 69
rect 139 65 143 67
rect 145 65 149 67
rect 139 63 149 65
<< nmos >>
rect 9 7 11 26
rect 19 7 21 26
rect 29 7 31 26
rect 40 7 42 20
rect 50 7 52 24
rect 60 7 62 24
rect 70 12 72 26
rect 83 10 85 26
rect 93 6 95 24
rect 103 6 105 24
rect 113 6 115 26
rect 130 16 132 26
rect 140 16 142 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 46 38 48 66
rect 56 38 58 66
rect 63 38 65 66
rect 73 38 75 66
rect 80 38 82 66
rect 90 38 92 66
rect 97 38 99 66
rect 107 38 109 66
rect 114 38 116 66
rect 124 38 126 58
rect 131 38 133 58
<< polyct0 >>
rect 105 31 107 33
<< polyct1 >>
rect 20 31 22 33
rect 27 31 29 33
rect 38 31 40 33
rect 68 31 70 33
rect 82 31 84 33
rect 115 31 117 33
rect 132 31 134 33
<< ndifct0 >>
rect 4 14 6 16
rect 24 14 26 16
rect 45 16 47 18
rect 55 9 57 11
rect 65 19 67 21
rect 77 14 79 16
rect 88 19 90 21
rect 98 8 100 10
rect 108 15 110 17
rect 135 19 137 21
rect 145 18 147 20
rect 122 8 124 10
<< ndifct1 >>
rect 14 22 16 24
rect 34 22 36 24
<< ntiect1 >>
rect 143 65 145 67
<< ptiect1 >>
rect 134 5 136 7
rect 145 5 147 7
<< pdifct0 >>
rect 14 62 16 64
rect 14 55 16 57
rect 24 54 26 56
rect 34 62 36 64
rect 34 55 36 57
rect 68 62 70 64
rect 68 55 70 57
rect 102 62 104 64
rect 102 55 104 57
rect 119 54 121 56
rect 136 54 138 56
rect 136 47 138 49
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 24 47 26 49
rect 51 54 53 56
rect 51 47 53 49
rect 85 54 87 56
rect 85 47 87 49
rect 119 47 121 49
<< alu0 >>
rect 12 62 14 64
rect 16 62 18 64
rect 12 57 18 62
rect 32 62 34 64
rect 36 62 38 64
rect 12 55 14 57
rect 16 55 18 57
rect 12 54 18 55
rect 23 56 27 58
rect 23 54 24 56
rect 26 54 27 56
rect 32 57 38 62
rect 66 62 68 64
rect 70 62 72 64
rect 32 55 34 57
rect 36 55 38 57
rect 32 54 38 55
rect 66 57 72 62
rect 100 62 102 64
rect 104 62 106 64
rect 66 55 68 57
rect 70 55 72 57
rect 66 54 72 55
rect 100 57 106 62
rect 100 55 102 57
rect 104 55 106 57
rect 100 54 106 55
rect 118 56 123 58
rect 118 54 119 56
rect 121 54 123 56
rect 23 50 27 54
rect 118 50 123 54
rect 134 56 140 64
rect 134 54 136 56
rect 138 54 140 56
rect 134 49 140 54
rect 134 47 136 49
rect 138 47 140 49
rect 134 46 140 47
rect 6 38 7 46
rect 103 33 109 38
rect 103 31 105 33
rect 107 31 109 33
rect 103 30 109 31
rect 44 21 91 25
rect 44 18 48 21
rect 44 17 45 18
rect 2 16 45 17
rect 47 16 48 18
rect 64 19 65 21
rect 67 19 68 21
rect 64 17 68 19
rect 87 19 88 21
rect 90 19 91 21
rect 87 18 91 19
rect 134 21 138 23
rect 134 19 135 21
rect 137 19 138 21
rect 134 18 138 19
rect 87 17 138 18
rect 2 14 4 16
rect 6 14 24 16
rect 26 14 48 16
rect 2 13 48 14
rect 75 16 81 17
rect 75 14 77 16
rect 79 14 81 16
rect 87 15 108 17
rect 110 15 138 17
rect 87 14 138 15
rect 144 20 148 22
rect 144 18 145 20
rect 147 18 148 20
rect 54 11 58 13
rect 54 9 55 11
rect 57 9 58 11
rect 54 8 58 9
rect 75 8 81 14
rect 96 10 102 11
rect 96 8 98 10
rect 100 8 102 10
rect 120 10 126 11
rect 120 8 122 10
rect 124 8 126 10
rect 144 8 148 18
<< labels >>
rlabel ndifct0 25 15 25 15 6 n1
rlabel alu0 46 19 46 19 6 n1
rlabel alu0 89 19 89 19 6 n1
rlabel alu0 67 23 67 23 6 n1
rlabel alu0 112 16 112 16 6 n1
rlabel alu0 136 18 136 18 6 n1
rlabel alu1 20 24 20 24 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 32 20 32 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 36 24 36 24 6 z
rlabel alu1 52 32 52 32 6 a1
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 28 36 28 36 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 76 4 76 4 6 vss
rlabel alu1 84 32 84 32 6 a2
rlabel alu1 68 32 68 32 6 a1
rlabel alu1 60 32 60 32 6 a1
rlabel alu1 84 40 84 40 6 a1
rlabel alu1 76 40 76 40 6 a1
rlabel alu1 60 48 60 48 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 76 48 76 48 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 76 68 76 68 6 vdd
rlabel alu1 108 24 108 24 6 a2
rlabel alu1 100 24 100 24 6 a2
rlabel alu1 116 28 116 28 6 a2
rlabel alu1 92 32 92 32 6 a2
rlabel alu1 92 40 92 40 6 a1
rlabel alu1 116 40 116 40 6 a1
rlabel alu1 108 40 108 40 6 a1
rlabel alu1 100 40 100 40 6 a1
rlabel alu1 92 48 92 48 6 z
rlabel alu1 116 48 116 48 6 z
rlabel alu1 108 48 108 48 6 z
rlabel alu1 100 48 100 48 6 z
rlabel alu1 124 40 124 40 6 a1
rlabel alu1 132 36 132 36 6 a1
rlabel alu1 124 48 124 48 6 z
<< end >>
