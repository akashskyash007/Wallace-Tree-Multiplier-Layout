magic
tech scmos
timestamp 1199980722
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -8 40 104 97
<< pwell >>
rect -8 -9 104 40
<< poly >>
rect 5 84 14 86
rect 5 82 7 84
rect 9 82 14 84
rect 5 80 14 82
rect 18 84 27 86
rect 18 82 23 84
rect 25 82 27 84
rect 18 80 27 82
rect 37 80 46 86
rect 50 80 59 86
rect 69 84 78 86
rect 69 82 71 84
rect 73 82 78 84
rect 69 80 78 82
rect 82 80 91 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 42 11 48
rect 15 42 30 48
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 66 46 75 48
rect 66 44 71 46
rect 73 44 75 46
rect 66 42 75 44
rect 79 46 94 48
rect 79 44 87 46
rect 89 44 94 46
rect 79 42 94 44
rect 2 32 17 38
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 66 36 81 38
rect 66 34 71 36
rect 73 34 81 36
rect 66 32 81 34
rect 85 36 94 38
rect 85 34 87 36
rect 89 34 94 36
rect 85 32 94 34
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
rect 69 2 78 8
rect 82 2 91 8
<< ndif >>
rect 2 11 9 29
rect 11 23 21 29
rect 11 21 15 23
rect 17 21 21 23
rect 11 16 21 21
rect 11 14 15 16
rect 17 14 21 16
rect 11 11 21 14
rect 23 24 30 29
rect 23 22 26 24
rect 28 22 30 24
rect 23 17 30 22
rect 23 15 26 17
rect 28 15 30 17
rect 23 11 30 15
rect 34 16 41 29
rect 34 14 36 16
rect 38 14 41 16
rect 34 11 41 14
rect 43 11 53 29
rect 55 25 62 29
rect 55 23 58 25
rect 60 23 62 25
rect 55 17 62 23
rect 55 15 58 17
rect 60 15 62 17
rect 55 11 62 15
rect 66 25 73 29
rect 66 23 68 25
rect 70 23 73 25
rect 66 17 73 23
rect 66 15 68 17
rect 70 15 73 17
rect 66 11 73 15
rect 75 27 85 29
rect 75 25 79 27
rect 81 25 85 27
rect 75 20 85 25
rect 75 18 79 20
rect 81 18 85 20
rect 75 11 85 18
rect 87 23 94 29
rect 87 21 90 23
rect 92 21 94 23
rect 87 16 94 21
rect 87 14 90 16
rect 92 14 94 16
rect 87 11 94 14
<< pdif >>
rect 2 51 9 77
rect 11 51 21 77
rect 23 51 30 77
rect 34 70 41 77
rect 34 68 36 70
rect 38 68 41 70
rect 34 51 41 68
rect 43 55 53 77
rect 43 53 47 55
rect 49 53 53 55
rect 43 51 53 53
rect 55 63 62 77
rect 55 61 58 63
rect 60 61 62 63
rect 55 51 62 61
rect 66 70 73 77
rect 66 68 68 70
rect 70 68 73 70
rect 66 55 73 68
rect 66 53 68 55
rect 70 53 73 55
rect 66 51 73 53
rect 75 73 85 77
rect 75 71 79 73
rect 81 71 85 73
rect 75 51 85 71
rect 87 71 94 77
rect 87 69 90 71
rect 92 69 94 71
rect 87 64 94 69
rect 87 62 90 64
rect 92 62 94 64
rect 87 51 94 62
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 84 31 85
rect 1 83 7 84
rect -2 82 7 83
rect 9 82 23 84
rect 25 83 31 84
rect 33 83 34 85
rect 25 82 34 83
rect -2 81 34 82
rect 62 85 66 90
rect 94 85 98 90
rect 62 83 63 85
rect 65 83 66 85
rect 62 81 66 83
rect 22 36 26 76
rect 78 83 95 85
rect 97 83 98 85
rect 78 81 98 83
rect 78 73 82 81
rect 78 71 79 73
rect 81 71 82 73
rect 22 34 23 36
rect 25 34 26 36
rect 22 32 26 34
rect 78 69 82 71
rect 46 55 50 57
rect 46 53 47 55
rect 49 53 50 55
rect 14 23 18 25
rect 14 21 15 23
rect 17 21 18 23
rect 14 16 18 21
rect 14 14 15 16
rect 17 14 18 16
rect 14 7 18 14
rect 46 26 50 53
rect 86 46 90 51
rect 86 44 87 46
rect 89 44 90 46
rect 86 36 90 44
rect 86 34 87 36
rect 89 34 90 36
rect 86 29 90 34
rect 46 25 72 26
rect 46 23 58 25
rect 60 23 68 25
rect 70 23 72 25
rect 46 22 72 23
rect 46 18 50 22
rect 35 16 39 18
rect 35 14 36 16
rect 38 14 39 16
rect 46 17 72 18
rect 46 15 58 17
rect 60 15 68 17
rect 70 15 72 17
rect 89 23 93 25
rect 89 21 90 23
rect 92 21 93 23
rect 89 16 93 21
rect 46 14 72 15
rect 89 14 90 16
rect 92 14 93 16
rect 35 7 39 14
rect 89 7 93 14
rect -2 6 39 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 5 39 6
rect 9 4 31 5
rect 1 3 31 4
rect 33 3 39 5
rect 57 5 66 7
rect 57 3 63 5
rect 65 3 66 5
rect 89 5 98 7
rect 89 3 95 5
rect 97 3 98 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 -2 66 3
rect 94 -2 98 3
<< alu2 >>
rect -2 85 98 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 95 85
rect 97 83 98 85
rect -2 80 98 83
rect -2 5 98 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 95 5
rect 97 3 98 5
rect -2 -2 98 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
rect 93 5 99 7
rect 93 3 95 5
rect 97 3 99 5
rect 93 0 99 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
rect 93 85 99 88
rect 93 83 95 85
rect 97 83 99 85
rect 93 81 99 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polyct0 >>
rect 71 82 73 84
rect 39 44 41 46
rect 55 44 57 46
rect 71 44 73 46
rect 39 34 41 36
rect 55 34 57 36
rect 71 34 73 36
<< polyct1 >>
rect 7 82 9 84
rect 23 82 25 84
rect 87 44 89 46
rect 23 34 25 36
rect 87 34 89 36
rect 7 4 9 6
<< ndifct0 >>
rect 26 22 28 24
rect 26 15 28 17
rect 79 25 81 27
rect 79 18 81 20
<< ndifct1 >>
rect 15 21 17 23
rect 15 14 17 16
rect 36 14 38 16
rect 58 23 60 25
rect 58 15 60 17
rect 68 23 70 25
rect 68 15 70 17
rect 90 21 92 23
rect 90 14 92 16
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< pdifct0 >>
rect 36 68 38 70
rect 58 61 60 63
rect 68 68 70 70
rect 68 53 70 55
rect 90 69 92 71
rect 90 62 92 64
<< pdifct1 >>
rect 47 53 49 55
rect 79 71 81 73
<< alu0 >>
rect 69 84 75 85
rect 69 82 71 84
rect 73 82 75 84
rect 69 78 75 82
rect 22 76 75 78
rect 26 74 75 76
rect 30 70 72 71
rect 30 68 36 70
rect 38 68 68 70
rect 70 68 72 70
rect 89 71 93 73
rect 89 69 90 71
rect 92 69 93 71
rect 30 67 72 68
rect 30 26 34 67
rect 89 64 93 69
rect 38 63 90 64
rect 38 61 58 63
rect 60 62 90 63
rect 92 62 93 64
rect 60 61 93 62
rect 38 60 93 61
rect 38 46 42 60
rect 38 44 39 46
rect 41 44 42 46
rect 38 36 42 44
rect 38 34 39 36
rect 41 34 42 36
rect 38 32 42 34
rect 25 24 34 26
rect 25 22 26 24
rect 28 22 34 24
rect 54 55 72 56
rect 54 53 68 55
rect 70 53 72 55
rect 54 52 72 53
rect 54 46 58 52
rect 54 44 55 46
rect 57 44 58 46
rect 54 36 58 44
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 70 46 74 48
rect 70 44 71 46
rect 73 44 74 46
rect 70 36 74 44
rect 70 34 71 36
rect 73 34 74 36
rect 70 32 74 34
rect 78 27 82 60
rect 78 25 79 27
rect 81 25 82 27
rect 25 17 29 22
rect 78 20 82 25
rect 78 18 79 20
rect 81 18 82 20
rect 25 15 26 17
rect 28 15 29 17
rect 25 13 29 15
rect 78 16 82 18
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< labels >>
rlabel alu1 24 56 24 56 6 b
rlabel alu1 64 16 64 16 6 z
rlabel alu1 56 16 56 16 6 z
rlabel alu1 56 24 56 24 6 z
rlabel alu1 64 24 64 24 6 z
rlabel alu1 48 36 48 36 6 z
rlabel alu1 88 40 88 40 6 a
rlabel alu2 48 4 48 4 6 vss
rlabel alu2 48 84 48 84 6 vdd
<< end >>
