magic
tech scmos
timestamp 1199541540
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -2 48 52 104
<< pwell >>
rect -2 -4 52 48
<< poly >>
rect 35 95 37 98
rect 11 85 13 88
rect 23 85 25 88
rect 11 63 13 65
rect 7 61 13 63
rect 7 59 9 61
rect 11 59 13 61
rect 7 57 13 59
rect 23 53 25 65
rect 23 51 31 53
rect 23 49 27 51
rect 29 49 31 51
rect 23 47 31 49
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 35 41 37 55
rect 17 39 19 41
rect 21 39 37 41
rect 17 37 23 39
rect 11 35 13 37
rect 23 31 31 33
rect 23 29 27 31
rect 29 29 31 31
rect 23 27 31 29
rect 23 25 25 27
rect 35 25 37 39
rect 11 12 13 15
rect 23 2 25 5
rect 35 2 37 5
<< ndif >>
rect 3 21 11 35
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 25 21 35
rect 13 15 23 25
rect 15 5 23 15
rect 25 11 35 25
rect 25 9 29 11
rect 31 9 35 11
rect 25 5 35 9
rect 37 21 45 25
rect 37 19 41 21
rect 43 19 45 21
rect 37 5 45 19
<< pdif >>
rect 3 91 9 93
rect 3 89 5 91
rect 7 89 9 91
rect 3 85 9 89
rect 27 91 35 95
rect 27 89 29 91
rect 31 89 35 91
rect 27 85 35 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 65 11 79
rect 13 81 23 85
rect 13 79 17 81
rect 19 79 23 81
rect 13 65 23 79
rect 25 65 35 85
rect 27 55 35 65
rect 37 81 45 95
rect 37 79 41 81
rect 43 79 45 81
rect 37 71 45 79
rect 37 69 41 71
rect 43 69 45 71
rect 37 61 45 69
rect 37 59 41 61
rect 43 59 45 61
rect 37 55 45 59
<< alu1 >>
rect -2 91 52 100
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 52 91
rect -2 88 52 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 78 8 79
rect 16 81 20 82
rect 16 79 17 81
rect 19 79 20 81
rect 16 78 20 79
rect 8 61 12 72
rect 8 59 9 61
rect 11 59 12 61
rect 8 41 12 59
rect 8 39 9 41
rect 11 39 12 41
rect 8 28 12 39
rect 18 42 20 78
rect 28 52 32 82
rect 26 51 32 52
rect 26 49 27 51
rect 29 49 32 51
rect 26 48 32 49
rect 18 41 22 42
rect 18 39 19 41
rect 21 39 22 41
rect 18 38 22 39
rect 4 21 8 22
rect 18 21 20 38
rect 28 32 32 48
rect 26 31 32 32
rect 26 29 27 31
rect 29 29 32 31
rect 26 28 32 29
rect 4 19 5 21
rect 7 19 20 21
rect 4 18 8 19
rect 28 18 32 28
rect 38 81 44 82
rect 38 79 41 81
rect 43 79 44 81
rect 38 78 44 79
rect 38 72 42 78
rect 38 71 44 72
rect 38 69 41 71
rect 43 69 44 71
rect 38 68 44 69
rect 38 62 42 68
rect 38 61 44 62
rect 38 59 41 61
rect 43 59 44 61
rect 38 58 44 59
rect 38 22 42 58
rect 38 21 44 22
rect 38 19 41 21
rect 43 19 44 21
rect 38 18 44 19
rect -2 11 52 12
rect -2 9 29 11
rect 31 9 52 11
rect -2 0 52 9
<< nmos >>
rect 11 15 13 35
rect 23 5 25 25
rect 35 5 37 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 55 37 95
<< polyct1 >>
rect 9 59 11 61
rect 27 49 29 51
rect 9 39 11 41
rect 19 39 21 41
rect 27 29 29 31
<< ndifct1 >>
rect 5 19 7 21
rect 29 9 31 11
rect 41 19 43 21
<< pdifct1 >>
rect 5 89 7 91
rect 29 89 31 91
rect 5 79 7 81
rect 17 79 19 81
rect 41 79 43 81
rect 41 69 43 71
rect 41 59 43 61
<< labels >>
rlabel alu1 10 50 10 50 6 i0
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 50 30 50 6 i1
rlabel alu1 25 94 25 94 6 vdd
rlabel alu1 40 50 40 50 6 q
<< end >>
