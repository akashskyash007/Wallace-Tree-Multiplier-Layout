magic
tech scmos
timestamp 1199203489
<< ab >>
rect 0 0 168 72
<< nwell >>
rect -5 32 173 77
<< pwell >>
rect -5 -5 173 32
<< poly >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 50 66 52 70
rect 60 66 62 70
rect 67 66 69 70
rect 77 66 79 70
rect 87 66 89 70
rect 117 66 119 70
rect 127 66 129 70
rect 137 66 139 70
rect 147 66 149 70
rect 97 57 99 61
rect 107 57 109 61
rect 157 57 159 61
rect 9 35 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 33 35 35 38
rect 43 35 45 38
rect 5 33 11 35
rect 5 31 7 33
rect 9 31 11 33
rect 5 29 11 31
rect 15 33 28 35
rect 32 33 45 35
rect 50 35 52 38
rect 60 35 62 38
rect 67 35 69 38
rect 77 35 79 38
rect 87 35 89 38
rect 97 35 99 38
rect 50 33 62 35
rect 66 33 72 35
rect 15 18 17 33
rect 32 31 34 33
rect 36 31 38 33
rect 32 29 38 31
rect 26 25 28 29
rect 36 25 38 29
rect 46 25 48 29
rect 56 25 58 33
rect 66 31 68 33
rect 70 31 72 33
rect 66 29 72 31
rect 76 33 99 35
rect 66 25 68 29
rect 76 25 78 33
rect 88 31 95 33
rect 97 31 99 33
rect 88 29 99 31
rect 107 35 109 38
rect 117 35 119 38
rect 127 35 129 38
rect 137 35 139 38
rect 147 35 149 38
rect 157 35 159 38
rect 107 33 129 35
rect 107 31 123 33
rect 125 31 129 33
rect 107 29 129 31
rect 133 33 159 35
rect 133 31 135 33
rect 137 31 139 33
rect 133 29 139 31
rect 88 25 90 29
rect 109 26 111 29
rect 119 26 121 29
rect 11 16 17 18
rect 11 14 13 16
rect 15 14 17 16
rect 11 12 17 14
rect 15 4 17 12
rect 26 11 28 14
rect 36 11 38 14
rect 26 9 38 11
rect 46 4 48 7
rect 56 4 58 7
rect 66 4 68 9
rect 15 2 58 4
rect 76 2 78 6
rect 88 2 90 6
rect 109 2 111 7
rect 119 2 121 7
<< ndif >>
rect 19 23 26 25
rect 19 21 21 23
rect 23 21 26 23
rect 19 19 26 21
rect 21 14 26 19
rect 28 18 36 25
rect 28 16 31 18
rect 33 16 36 18
rect 28 14 36 16
rect 38 23 46 25
rect 38 21 41 23
rect 43 21 46 23
rect 38 14 46 21
rect 41 7 46 14
rect 48 23 56 25
rect 48 21 51 23
rect 53 21 56 23
rect 48 7 56 21
rect 58 23 66 25
rect 58 21 61 23
rect 63 21 66 23
rect 58 9 66 21
rect 68 16 76 25
rect 68 14 71 16
rect 73 14 76 16
rect 68 9 76 14
rect 58 7 63 9
rect 71 6 76 9
rect 78 7 88 25
rect 78 6 82 7
rect 80 5 82 6
rect 84 6 88 7
rect 90 18 95 25
rect 90 16 97 18
rect 90 14 93 16
rect 95 14 97 16
rect 90 12 97 14
rect 90 6 95 12
rect 101 7 109 26
rect 111 24 119 26
rect 111 22 114 24
rect 116 22 119 24
rect 111 7 119 22
rect 121 7 129 26
rect 84 5 86 6
rect 80 3 86 5
rect 101 5 103 7
rect 105 5 107 7
rect 101 3 107 5
rect 123 5 125 7
rect 127 5 129 7
rect 123 3 129 5
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 38 16 66
rect 18 64 26 66
rect 18 62 21 64
rect 23 62 26 64
rect 18 38 26 62
rect 28 38 33 66
rect 35 57 43 66
rect 35 55 38 57
rect 40 55 43 57
rect 35 42 43 55
rect 35 40 38 42
rect 40 40 43 42
rect 35 38 43 40
rect 45 38 50 66
rect 52 64 60 66
rect 52 62 55 64
rect 57 62 60 64
rect 52 38 60 62
rect 62 38 67 66
rect 69 57 77 66
rect 69 55 72 57
rect 74 55 77 57
rect 69 42 77 55
rect 69 40 72 42
rect 74 40 77 42
rect 69 38 77 40
rect 79 49 87 66
rect 79 47 82 49
rect 84 47 87 49
rect 79 42 87 47
rect 79 40 82 42
rect 84 40 87 42
rect 79 38 87 40
rect 89 57 94 66
rect 112 57 117 66
rect 89 55 97 57
rect 89 53 92 55
rect 94 53 97 55
rect 89 38 97 53
rect 99 49 107 57
rect 99 47 102 49
rect 104 47 107 49
rect 99 42 107 47
rect 99 40 102 42
rect 104 40 107 42
rect 99 38 107 40
rect 109 55 117 57
rect 109 53 112 55
rect 114 53 117 55
rect 109 38 117 53
rect 119 56 127 66
rect 119 54 122 56
rect 124 54 127 56
rect 119 49 127 54
rect 119 47 122 49
rect 124 47 127 49
rect 119 38 127 47
rect 129 64 137 66
rect 129 62 132 64
rect 134 62 137 64
rect 129 57 137 62
rect 129 55 132 57
rect 134 55 137 57
rect 129 38 137 55
rect 139 49 147 66
rect 139 47 142 49
rect 144 47 147 49
rect 139 42 147 47
rect 139 40 142 42
rect 144 40 147 42
rect 139 38 147 40
rect 149 57 154 66
rect 149 55 157 57
rect 149 53 152 55
rect 154 53 157 55
rect 149 38 157 53
rect 159 51 164 57
rect 159 49 166 51
rect 159 47 162 49
rect 164 47 166 49
rect 159 42 166 47
rect 159 40 162 42
rect 164 40 166 42
rect 159 38 166 40
<< alu1 >>
rect -2 67 170 72
rect -2 65 102 67
rect 104 65 161 67
rect 163 65 170 67
rect -2 64 170 65
rect 17 57 95 58
rect 17 55 38 57
rect 40 55 72 57
rect 74 55 95 57
rect 17 54 92 55
rect 17 50 23 54
rect 91 53 92 54
rect 94 53 95 55
rect 91 51 95 53
rect 2 49 23 50
rect 2 47 4 49
rect 6 47 23 49
rect 2 46 23 47
rect 2 42 7 46
rect 2 40 4 42
rect 6 40 7 42
rect 2 37 7 40
rect 113 38 135 42
rect 113 34 117 38
rect 131 34 135 38
rect 93 33 117 34
rect 93 31 95 33
rect 97 31 117 33
rect 93 30 117 31
rect 121 33 127 34
rect 121 31 123 33
rect 125 31 127 33
rect 121 26 127 31
rect 131 33 139 34
rect 131 31 135 33
rect 137 31 139 33
rect 131 30 139 31
rect 121 22 135 26
rect -2 7 170 8
rect -2 5 5 7
rect 7 5 82 7
rect 84 5 103 7
rect 105 5 125 7
rect 127 5 153 7
rect 155 5 161 7
rect 163 5 170 7
rect -2 0 170 5
<< ptie >>
rect 3 7 9 24
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 151 7 165 9
rect 151 5 153 7
rect 155 5 161 7
rect 163 5 165 7
rect 151 3 165 5
<< ntie >>
rect 98 67 108 69
rect 98 65 102 67
rect 104 65 108 67
rect 159 67 165 69
rect 98 63 108 65
rect 159 65 161 67
rect 163 65 165 67
rect 159 63 165 65
<< nmos >>
rect 26 14 28 25
rect 36 14 38 25
rect 46 7 48 25
rect 56 7 58 25
rect 66 9 68 25
rect 76 6 78 25
rect 88 6 90 25
rect 109 7 111 26
rect 119 7 121 26
<< pmos >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 38 45 66
rect 50 38 52 66
rect 60 38 62 66
rect 67 38 69 66
rect 77 38 79 66
rect 87 38 89 66
rect 97 38 99 57
rect 107 38 109 57
rect 117 38 119 66
rect 127 38 129 66
rect 137 38 139 66
rect 147 38 149 66
rect 157 38 159 57
<< polyct0 >>
rect 7 31 9 33
rect 34 31 36 33
rect 68 31 70 33
rect 13 14 15 16
<< polyct1 >>
rect 95 31 97 33
rect 123 31 125 33
rect 135 31 137 33
<< ndifct0 >>
rect 21 21 23 23
rect 31 16 33 18
rect 41 21 43 23
rect 51 21 53 23
rect 61 21 63 23
rect 71 14 73 16
rect 93 14 95 16
rect 114 22 116 24
<< ndifct1 >>
rect 82 5 84 7
rect 103 5 105 7
rect 125 5 127 7
<< ntiect1 >>
rect 102 65 104 67
rect 161 65 163 67
<< ptiect1 >>
rect 5 5 7 7
rect 153 5 155 7
rect 161 5 163 7
<< pdifct0 >>
rect 21 62 23 64
rect 38 40 40 42
rect 55 62 57 64
rect 72 40 74 42
rect 82 47 84 49
rect 82 40 84 42
rect 102 47 104 49
rect 102 40 104 42
rect 112 53 114 55
rect 122 54 124 56
rect 122 47 124 49
rect 132 62 134 64
rect 132 55 134 57
rect 142 47 144 49
rect 142 40 144 42
rect 152 53 154 55
rect 162 47 164 49
rect 162 40 164 42
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 38 55 40 57
rect 72 55 74 57
rect 92 53 94 55
<< alu0 >>
rect 19 62 21 64
rect 23 62 25 64
rect 19 61 25 62
rect 53 62 55 64
rect 57 62 59 64
rect 53 61 59 62
rect 110 55 116 64
rect 131 62 132 64
rect 134 62 135 64
rect 110 53 112 55
rect 114 53 116 55
rect 110 52 116 53
rect 121 56 125 58
rect 121 54 122 56
rect 124 54 125 56
rect 28 49 86 50
rect 28 47 82 49
rect 84 47 86 49
rect 28 46 86 47
rect 28 34 32 46
rect 36 42 45 43
rect 36 40 38 42
rect 40 40 45 42
rect 36 39 45 40
rect 5 33 38 34
rect 5 31 7 33
rect 9 31 34 33
rect 36 31 38 33
rect 5 30 38 31
rect 41 26 45 39
rect 19 23 45 26
rect 19 21 21 23
rect 23 22 41 23
rect 23 21 25 22
rect 19 20 25 21
rect 39 21 41 22
rect 43 21 45 23
rect 39 20 45 21
rect 49 24 53 46
rect 59 42 76 43
rect 59 40 72 42
rect 74 40 76 42
rect 59 39 76 40
rect 81 42 86 46
rect 101 49 105 51
rect 121 49 125 54
rect 131 57 135 62
rect 131 55 132 57
rect 134 55 135 57
rect 131 53 135 55
rect 151 55 155 64
rect 151 53 152 55
rect 154 53 155 55
rect 151 51 155 53
rect 101 47 102 49
rect 104 47 122 49
rect 124 47 125 49
rect 101 45 125 47
rect 141 49 145 51
rect 141 47 142 49
rect 144 47 145 49
rect 101 42 105 45
rect 141 42 145 47
rect 161 49 165 51
rect 161 47 162 49
rect 164 47 165 49
rect 161 42 165 47
rect 81 40 82 42
rect 84 40 102 42
rect 104 40 105 42
rect 59 24 63 39
rect 81 38 105 40
rect 141 40 142 42
rect 144 40 162 42
rect 164 40 165 42
rect 141 38 165 40
rect 81 34 85 38
rect 66 33 85 34
rect 66 31 68 33
rect 70 31 85 33
rect 66 30 85 31
rect 81 25 85 30
rect 81 24 118 25
rect 49 23 55 24
rect 49 21 51 23
rect 53 21 55 23
rect 49 20 55 21
rect 59 23 65 24
rect 59 21 61 23
rect 63 21 65 23
rect 81 22 114 24
rect 116 22 118 24
rect 81 21 118 22
rect 59 20 65 21
rect 29 18 35 19
rect 29 17 31 18
rect 11 16 31 17
rect 33 17 35 18
rect 143 17 147 38
rect 33 16 147 17
rect 11 14 13 16
rect 15 14 71 16
rect 73 14 93 16
rect 95 14 147 16
rect 11 13 147 14
<< labels >>
rlabel alu0 21 32 21 32 6 an
rlabel alu0 51 35 51 35 6 an
rlabel alu0 99 23 99 23 6 an
rlabel alu0 75 32 75 32 6 an
rlabel alu0 103 44 103 44 6 an
rlabel alu0 83 35 83 35 6 an
rlabel alu0 79 15 79 15 6 bn
rlabel alu0 163 44 163 44 6 bn
rlabel alu0 143 44 143 44 6 bn
rlabel alu0 123 51 123 51 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 60 56 60 56 6 z
rlabel alu1 52 56 52 56 6 z
rlabel alu1 76 56 76 56 6 z
rlabel alu1 68 56 68 56 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 84 4 84 4 6 vss
rlabel alu1 100 32 100 32 6 b
rlabel alu1 108 32 108 32 6 b
rlabel alu1 124 28 124 28 6 a
rlabel alu1 116 40 116 40 6 b
rlabel alu1 124 40 124 40 6 b
rlabel alu1 92 56 92 56 6 z
rlabel alu1 84 56 84 56 6 z
rlabel alu1 84 68 84 68 6 vdd
rlabel alu1 132 24 132 24 6 a
rlabel alu1 132 40 132 40 6 b
<< end >>
