magic
tech scmos
timestamp 1199542932
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -5 48 105 105
<< pwell >>
rect -5 -5 105 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 75 94 77 98
rect 87 94 89 98
rect 11 53 13 56
rect 23 53 25 56
rect 35 53 37 56
rect 47 53 49 56
rect 75 53 77 56
rect 87 53 89 56
rect 11 51 19 53
rect 23 51 29 53
rect 35 51 43 53
rect 17 43 19 51
rect 27 43 29 51
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 75 51 81 53
rect 75 49 77 51
rect 79 49 81 51
rect 75 47 81 49
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 17 29 19 37
rect 27 29 29 37
rect 37 29 39 47
rect 47 29 49 47
rect 15 27 19 29
rect 23 27 29 29
rect 35 27 39 29
rect 43 27 49 29
rect 15 24 17 27
rect 23 24 25 27
rect 35 24 37 27
rect 43 24 45 27
rect 79 25 81 47
rect 87 51 93 53
rect 87 49 89 51
rect 91 49 93 51
rect 87 47 93 49
rect 87 25 89 47
rect 15 2 17 6
rect 23 2 25 6
rect 35 2 37 6
rect 43 2 45 6
rect 79 2 81 6
rect 87 2 89 6
<< ndif >>
rect 7 11 15 24
rect 7 9 9 11
rect 11 9 15 11
rect 7 6 15 9
rect 17 6 23 24
rect 25 21 35 24
rect 25 19 29 21
rect 31 19 35 21
rect 25 6 35 19
rect 37 6 43 24
rect 45 11 53 24
rect 71 21 79 25
rect 71 19 73 21
rect 75 19 79 21
rect 45 9 49 11
rect 51 9 53 11
rect 45 6 53 9
rect 71 6 79 19
rect 81 6 87 25
rect 89 21 97 25
rect 89 19 93 21
rect 95 19 97 21
rect 89 11 97 19
rect 89 9 93 11
rect 95 9 97 11
rect 89 6 97 9
<< pdif >>
rect 3 81 11 94
rect 3 79 5 81
rect 7 79 11 81
rect 3 56 11 79
rect 13 71 23 94
rect 13 69 17 71
rect 19 69 23 71
rect 13 56 23 69
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 56 35 79
rect 37 71 47 94
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 49 81 57 94
rect 49 79 53 81
rect 55 79 57 81
rect 49 56 57 79
rect 67 81 75 94
rect 67 79 69 81
rect 71 79 75 81
rect 67 56 75 79
rect 77 81 87 94
rect 77 79 81 81
rect 83 79 87 81
rect 77 56 87 79
rect 89 91 97 94
rect 89 89 93 91
rect 95 89 97 91
rect 89 81 97 89
rect 89 79 93 81
rect 95 79 97 81
rect 89 71 97 79
rect 89 69 93 71
rect 95 69 97 71
rect 89 56 97 69
<< alu1 >>
rect -2 91 102 100
rect -2 89 93 91
rect 95 89 102 91
rect -2 88 102 89
rect 3 81 57 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 79 53 81
rect 55 79 57 81
rect 3 78 57 79
rect 68 81 72 88
rect 68 79 69 81
rect 71 79 72 81
rect 68 77 72 79
rect 80 81 84 83
rect 80 79 81 81
rect 83 79 84 81
rect 8 72 12 73
rect 8 71 21 72
rect 8 69 17 71
rect 19 69 21 71
rect 8 68 21 69
rect 8 22 12 68
rect 18 41 22 63
rect 18 39 19 41
rect 21 39 22 41
rect 18 27 22 39
rect 28 41 32 73
rect 80 72 84 79
rect 39 71 84 72
rect 39 69 41 71
rect 43 69 84 71
rect 39 68 84 69
rect 92 81 96 88
rect 92 79 93 81
rect 95 79 96 81
rect 92 71 96 79
rect 92 69 93 71
rect 95 69 96 71
rect 92 67 96 69
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 51 42 63
rect 38 49 39 51
rect 41 49 42 51
rect 38 27 42 49
rect 48 51 52 63
rect 78 52 82 63
rect 48 49 49 51
rect 51 49 52 51
rect 48 27 52 49
rect 75 51 82 52
rect 75 49 77 51
rect 79 49 82 51
rect 75 48 82 49
rect 78 27 82 48
rect 88 51 92 63
rect 88 49 89 51
rect 91 49 92 51
rect 88 27 92 49
rect 8 21 77 22
rect 8 19 29 21
rect 31 19 73 21
rect 75 19 77 21
rect 8 18 77 19
rect 92 21 96 23
rect 92 19 93 21
rect 95 19 96 21
rect 8 17 12 18
rect 92 12 96 19
rect -2 11 102 12
rect -2 9 9 11
rect 11 9 49 11
rect 51 9 93 11
rect 95 9 102 11
rect -2 7 61 9
rect 63 7 102 9
rect -2 0 102 7
<< ptie >>
rect 59 9 65 16
rect 59 7 61 9
rect 63 7 65 9
rect 59 5 65 7
<< nmos >>
rect 15 6 17 24
rect 23 6 25 24
rect 35 6 37 24
rect 43 6 45 24
rect 79 6 81 25
rect 87 6 89 25
<< pmos >>
rect 11 56 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 47 56 49 94
rect 75 56 77 94
rect 87 56 89 94
<< polyct1 >>
rect 39 49 41 51
rect 49 49 51 51
rect 77 49 79 51
rect 19 39 21 41
rect 29 39 31 41
rect 89 49 91 51
<< ndifct1 >>
rect 9 9 11 11
rect 29 19 31 21
rect 73 19 75 21
rect 49 9 51 11
rect 93 19 95 21
rect 93 9 95 11
<< ptiect1 >>
rect 61 7 63 9
<< pdifct1 >>
rect 5 79 7 81
rect 17 69 19 71
rect 29 79 31 81
rect 41 69 43 71
rect 53 79 55 81
rect 69 79 71 81
rect 81 79 83 81
rect 93 89 95 91
rect 93 79 95 81
rect 93 69 95 71
<< labels >>
rlabel alu1 20 20 20 20 6 nq
rlabel alu1 10 45 10 45 6 nq
rlabel alu1 20 45 20 45 6 i5
rlabel ndifct1 30 20 30 20 6 nq
rlabel alu1 40 20 40 20 6 nq
rlabel alu1 40 45 40 45 6 i3
rlabel alu1 30 50 30 50 6 i4
rlabel alu1 50 20 50 20 6 nq
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 60 20 60 20 6 nq
rlabel alu1 70 20 70 20 6 nq
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 50 94 50 94 6 vdd
rlabel alu1 80 45 80 45 6 i1
rlabel alu1 90 45 90 45 6 i0
<< end >>
