magic
tech scmos
timestamp 1199469740
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 33 94 35 98
rect 45 94 47 98
rect 57 94 59 98
rect 21 83 23 88
rect 57 63 59 66
rect 55 61 61 63
rect 55 59 57 61
rect 59 59 61 61
rect 55 57 61 59
rect 21 52 23 55
rect 33 52 35 55
rect 17 50 23 52
rect 17 48 19 50
rect 21 48 23 50
rect 13 46 23 48
rect 27 50 35 52
rect 27 48 29 50
rect 31 48 35 50
rect 45 52 47 55
rect 45 50 53 52
rect 45 48 49 50
rect 51 48 53 50
rect 27 46 39 48
rect 13 31 15 46
rect 37 39 39 46
rect 45 46 53 48
rect 45 39 47 46
rect 57 39 59 57
rect 13 12 15 17
rect 57 20 59 25
rect 37 2 39 6
rect 45 2 47 6
<< ndif >>
rect 32 33 37 39
rect 29 31 37 33
rect 5 29 13 31
rect 5 27 7 29
rect 9 27 13 29
rect 5 21 13 27
rect 5 19 7 21
rect 9 19 13 21
rect 5 17 13 19
rect 15 21 23 31
rect 15 19 19 21
rect 21 19 23 21
rect 15 17 23 19
rect 29 29 31 31
rect 33 29 37 31
rect 29 21 37 29
rect 29 19 31 21
rect 33 19 37 21
rect 29 17 37 19
rect 32 6 37 17
rect 39 6 45 39
rect 47 31 57 39
rect 47 29 51 31
rect 53 29 57 31
rect 47 25 57 29
rect 59 37 67 39
rect 59 35 63 37
rect 65 35 67 37
rect 59 29 67 35
rect 59 27 63 29
rect 65 27 67 29
rect 59 25 67 27
rect 47 21 55 25
rect 47 19 51 21
rect 53 19 55 21
rect 47 11 55 19
rect 47 9 51 11
rect 53 9 55 11
rect 47 6 55 9
<< pdif >>
rect 25 91 33 94
rect 25 89 27 91
rect 29 89 33 91
rect 25 83 33 89
rect 16 71 21 83
rect 13 69 21 71
rect 13 67 15 69
rect 17 67 21 69
rect 13 61 21 67
rect 13 59 15 61
rect 17 59 21 61
rect 13 57 21 59
rect 16 55 21 57
rect 23 81 33 83
rect 23 79 27 81
rect 29 79 33 81
rect 23 71 33 79
rect 23 69 27 71
rect 29 69 33 71
rect 23 55 33 69
rect 35 71 45 94
rect 35 69 39 71
rect 41 69 45 71
rect 35 61 45 69
rect 35 59 39 61
rect 41 59 45 61
rect 35 55 45 59
rect 47 91 57 94
rect 47 89 51 91
rect 53 89 57 91
rect 47 66 57 89
rect 59 73 64 94
rect 59 71 67 73
rect 59 69 63 71
rect 65 69 67 71
rect 59 66 67 69
rect 47 55 52 66
<< alu1 >>
rect -2 95 72 100
rect -2 93 5 95
rect 7 93 15 95
rect 17 93 72 95
rect -2 91 72 93
rect -2 89 27 91
rect 29 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 26 81 30 88
rect 26 79 27 81
rect 29 79 30 81
rect 26 71 30 79
rect 48 78 63 83
rect 14 69 18 71
rect 14 67 15 69
rect 17 67 18 69
rect 26 69 27 71
rect 29 69 30 71
rect 26 67 30 69
rect 38 71 42 73
rect 38 69 39 71
rect 41 69 42 71
rect 14 62 18 67
rect 6 61 32 62
rect 6 59 15 61
rect 17 59 32 61
rect 6 58 32 59
rect 6 29 10 58
rect 6 27 7 29
rect 9 27 10 29
rect 18 50 22 53
rect 18 48 19 50
rect 21 48 22 50
rect 18 42 22 48
rect 28 50 32 58
rect 28 48 29 50
rect 31 48 32 50
rect 28 46 32 48
rect 38 61 42 69
rect 38 59 39 61
rect 41 59 42 61
rect 18 38 33 42
rect 18 27 22 38
rect 38 33 42 59
rect 48 63 52 78
rect 61 71 68 73
rect 61 69 63 71
rect 65 69 68 71
rect 61 67 68 69
rect 48 61 60 63
rect 48 59 57 61
rect 59 59 60 61
rect 48 57 60 59
rect 64 51 68 67
rect 47 50 68 51
rect 47 48 49 50
rect 51 48 68 50
rect 47 47 68 48
rect 62 37 66 47
rect 62 35 63 37
rect 65 35 66 37
rect 28 31 42 33
rect 28 29 31 31
rect 33 29 42 31
rect 28 27 42 29
rect 50 31 54 33
rect 50 29 51 31
rect 53 29 54 31
rect 6 21 10 27
rect 6 19 7 21
rect 9 19 10 21
rect 6 17 10 19
rect 18 21 22 23
rect 18 19 19 21
rect 21 19 22 21
rect 18 12 22 19
rect 28 21 34 27
rect 28 19 31 21
rect 33 19 34 21
rect 28 17 34 19
rect 50 21 54 29
rect 62 29 66 35
rect 62 27 63 29
rect 65 27 66 29
rect 62 25 66 27
rect 50 19 51 21
rect 53 19 54 21
rect 50 12 54 19
rect -2 11 72 12
rect -2 9 51 11
rect 53 9 72 11
rect -2 7 72 9
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 72 7
rect -2 0 72 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 3 95 19 97
rect 3 93 5 95
rect 7 93 15 95
rect 17 93 19 95
rect 3 91 19 93
<< nmos >>
rect 13 17 15 31
rect 37 6 39 39
rect 45 6 47 39
rect 57 25 59 39
<< pmos >>
rect 21 55 23 83
rect 33 55 35 94
rect 45 55 47 94
rect 57 66 59 94
<< polyct1 >>
rect 57 59 59 61
rect 19 48 21 50
rect 29 48 31 50
rect 49 48 51 50
<< ndifct1 >>
rect 7 27 9 29
rect 7 19 9 21
rect 19 19 21 21
rect 31 29 33 31
rect 31 19 33 21
rect 51 29 53 31
rect 63 35 65 37
rect 63 27 65 29
rect 51 19 53 21
rect 51 9 53 11
<< ntiect1 >>
rect 5 93 7 95
rect 15 93 17 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 27 89 29 91
rect 15 67 17 69
rect 15 59 17 61
rect 27 79 29 81
rect 27 69 29 71
rect 39 69 41 71
rect 39 59 41 61
rect 51 89 53 91
rect 63 69 65 71
<< labels >>
rlabel ndifct1 8 20 8 20 6 bn
rlabel ndifct1 8 28 8 28 6 bn
rlabel pdifct1 16 68 16 68 6 bn
rlabel pdifct1 16 60 16 60 6 bn
rlabel ndifct1 64 28 64 28 6 an
rlabel ndifct1 64 36 64 36 6 an
rlabel polyct1 50 49 50 49 6 an
rlabel pdifct1 64 70 64 70 6 an
rlabel alu1 30 25 30 25 6 z
rlabel alu1 20 40 20 40 6 b
rlabel alu1 30 40 30 40 6 b
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 50 40 50 6 z
rlabel alu1 50 70 50 70 6 a
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 80 60 80 6 a
<< end >>
