magic
tech scmos
timestamp 1199202503
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 26 70 28 74
rect 36 70 38 74
rect 43 70 45 74
rect 56 57 62 59
rect 56 55 58 57
rect 60 55 62 57
rect 9 34 11 52
rect 19 44 21 54
rect 16 42 22 44
rect 16 40 18 42
rect 20 40 22 42
rect 16 38 22 40
rect 26 39 28 54
rect 36 49 38 54
rect 33 47 39 49
rect 33 45 35 47
rect 37 45 39 47
rect 33 43 39 45
rect 43 39 45 54
rect 53 53 62 55
rect 53 50 55 53
rect 8 32 14 34
rect 8 30 10 32
rect 12 30 14 32
rect 8 28 14 30
rect 9 25 11 28
rect 19 24 21 38
rect 26 37 38 39
rect 26 31 32 33
rect 26 29 28 31
rect 30 29 32 31
rect 26 27 32 29
rect 26 24 28 27
rect 36 24 38 37
rect 43 37 49 39
rect 43 35 45 37
rect 47 35 49 37
rect 43 33 49 35
rect 43 24 45 33
rect 53 24 55 42
rect 9 11 11 16
rect 19 11 21 16
rect 26 11 28 16
rect 36 8 38 16
rect 43 12 45 16
rect 53 8 55 18
rect 36 6 55 8
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 4 16 9 19
rect 11 24 16 25
rect 11 20 19 24
rect 11 18 14 20
rect 16 18 19 20
rect 11 16 19 18
rect 21 16 26 24
rect 28 20 36 24
rect 28 18 31 20
rect 33 18 36 20
rect 28 16 36 18
rect 38 16 43 24
rect 45 22 53 24
rect 45 20 48 22
rect 50 20 53 22
rect 45 18 53 20
rect 55 22 62 24
rect 55 20 58 22
rect 60 20 62 22
rect 55 18 62 20
rect 45 16 51 18
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 57 9 59
rect 4 52 9 57
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 54 19 66
rect 21 54 26 70
rect 28 58 36 70
rect 28 56 31 58
rect 33 56 36 58
rect 28 54 36 56
rect 38 54 43 70
rect 45 68 52 70
rect 45 66 48 68
rect 50 66 52 68
rect 45 58 52 66
rect 45 54 51 58
rect 11 52 16 54
rect 47 50 51 54
rect 47 42 53 50
rect 55 48 60 50
rect 55 46 62 48
rect 55 44 58 46
rect 60 44 62 46
rect 55 42 62 44
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 61 15 62
rect 2 59 4 61
rect 6 59 15 61
rect 2 58 15 59
rect 2 25 6 58
rect 57 57 62 63
rect 57 55 58 57
rect 60 55 62 57
rect 57 54 62 55
rect 49 50 62 54
rect 18 42 30 47
rect 20 41 30 42
rect 20 40 22 41
rect 18 33 22 40
rect 42 37 48 39
rect 42 35 45 37
rect 47 35 48 37
rect 42 30 48 35
rect 42 26 55 30
rect 2 23 7 25
rect 2 21 4 23
rect 6 21 7 23
rect 2 19 7 21
rect 2 17 6 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 16 11 25
rect 19 16 21 24
rect 26 16 28 24
rect 36 16 38 24
rect 43 16 45 24
rect 53 18 55 24
<< pmos >>
rect 9 52 11 70
rect 19 54 21 70
rect 26 54 28 70
rect 36 54 38 70
rect 43 54 45 70
rect 53 42 55 50
<< polyct0 >>
rect 35 45 37 47
rect 10 30 12 32
rect 28 29 30 31
<< polyct1 >>
rect 58 55 60 57
rect 18 40 20 42
rect 45 35 47 37
<< ndifct0 >>
rect 14 18 16 20
rect 31 18 33 20
rect 48 20 50 22
rect 58 20 60 22
<< ndifct1 >>
rect 4 21 6 23
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 14 66 16 68
rect 31 56 33 58
rect 48 66 50 68
rect 58 44 60 46
<< pdifct1 >>
rect 4 59 6 61
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 65 18 66
rect 47 66 48 68
rect 50 66 51 68
rect 47 64 51 66
rect 22 58 35 59
rect 22 56 31 58
rect 33 56 35 58
rect 22 55 35 56
rect 10 51 26 55
rect 10 34 14 51
rect 34 47 38 49
rect 17 38 18 44
rect 34 45 35 47
rect 37 46 62 47
rect 37 45 58 46
rect 34 44 58 45
rect 60 44 62 46
rect 34 43 62 44
rect 9 32 14 34
rect 34 33 38 43
rect 9 30 10 32
rect 12 30 14 32
rect 27 31 38 33
rect 9 28 24 30
rect 10 26 24 28
rect 27 29 28 31
rect 30 29 38 31
rect 27 27 38 29
rect 13 20 17 22
rect 13 18 14 20
rect 16 18 17 20
rect 13 12 17 18
rect 20 21 24 26
rect 58 23 62 43
rect 46 22 52 23
rect 20 20 35 21
rect 20 18 31 20
rect 33 18 35 20
rect 20 17 35 18
rect 46 20 48 22
rect 50 20 52 22
rect 46 12 52 20
rect 56 22 62 23
rect 56 20 58 22
rect 60 20 62 22
rect 56 19 62 20
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 27 19 27 19 6 zn
rlabel alu0 32 30 32 30 6 sn
rlabel alu0 36 38 36 38 6 sn
rlabel alu0 28 57 28 57 6 zn
rlabel alu0 60 33 60 33 6 sn
rlabel alu0 48 45 48 45 6 sn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 44 28 44 6 a0
rlabel alu1 20 40 20 40 6 a0
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 36 44 36 6 a1
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 a1
rlabel alu1 52 52 52 52 6 s
rlabel alu1 60 60 60 60 6 s
<< end >>
