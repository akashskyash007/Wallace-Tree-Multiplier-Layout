magic
tech scmos
timestamp 1199980718
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -8 40 104 97
<< pwell >>
rect -8 -9 104 40
<< poly >>
rect 5 84 14 86
rect 5 82 7 84
rect 9 82 14 84
rect 5 80 14 82
rect 18 84 27 86
rect 18 82 23 84
rect 25 82 27 84
rect 18 80 27 82
rect 37 80 46 86
rect 50 80 59 86
rect 69 84 78 86
rect 69 82 71 84
rect 73 82 78 84
rect 69 80 78 82
rect 82 80 91 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 42 11 48
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 66 42 75 48
rect 79 46 94 48
rect 79 44 87 46
rect 89 44 94 46
rect 79 42 94 44
rect 2 32 17 38
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 66 32 81 38
rect 85 36 94 38
rect 85 34 87 36
rect 89 34 94 36
rect 85 32 94 34
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 2 27 8
rect 37 2 46 8
rect 50 6 59 8
rect 50 4 52 6
rect 54 4 59 6
rect 50 2 59 4
rect 69 6 78 8
rect 69 4 71 6
rect 73 4 78 6
rect 69 2 78 4
rect 82 2 91 8
<< ndif >>
rect 2 11 9 29
rect 11 23 21 29
rect 11 21 15 23
rect 17 21 21 23
rect 11 16 21 21
rect 11 14 15 16
rect 17 14 21 16
rect 11 11 21 14
rect 23 25 30 29
rect 23 23 26 25
rect 28 23 30 25
rect 23 17 30 23
rect 23 15 26 17
rect 28 15 30 17
rect 23 11 30 15
rect 34 25 41 29
rect 34 23 36 25
rect 38 23 41 25
rect 34 17 41 23
rect 34 15 36 17
rect 38 15 41 17
rect 34 11 41 15
rect 43 25 53 29
rect 43 23 47 25
rect 49 23 53 25
rect 43 17 53 23
rect 43 15 47 17
rect 49 15 53 17
rect 43 11 53 15
rect 55 24 62 29
rect 55 22 58 24
rect 60 22 62 24
rect 55 17 62 22
rect 55 15 58 17
rect 60 15 62 17
rect 55 11 62 15
rect 66 11 73 29
rect 75 17 85 29
rect 75 15 79 17
rect 81 15 85 17
rect 75 11 85 15
rect 87 24 94 29
rect 87 22 90 24
rect 92 22 94 24
rect 87 17 94 22
rect 87 15 90 17
rect 92 15 94 17
rect 87 11 94 15
<< pdif >>
rect 2 51 9 77
rect 11 74 21 77
rect 11 72 15 74
rect 17 72 21 74
rect 11 67 21 72
rect 11 65 15 67
rect 17 65 21 67
rect 11 51 21 65
rect 23 62 30 77
rect 23 60 26 62
rect 28 60 30 62
rect 23 55 30 60
rect 23 53 26 55
rect 28 53 30 55
rect 23 51 30 53
rect 34 70 41 77
rect 34 68 36 70
rect 38 68 41 70
rect 34 51 41 68
rect 43 51 53 77
rect 55 55 62 77
rect 55 53 58 55
rect 60 53 62 55
rect 55 51 62 53
rect 66 55 73 77
rect 66 53 68 55
rect 70 53 73 55
rect 66 51 73 53
rect 75 62 85 77
rect 75 60 79 62
rect 81 60 85 62
rect 75 55 85 60
rect 75 53 79 55
rect 81 53 85 55
rect 75 51 85 53
rect 87 73 94 77
rect 87 71 90 73
rect 92 71 94 73
rect 87 66 94 71
rect 87 64 90 66
rect 92 64 94 66
rect 87 51 94 64
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 84 18 85
rect 1 83 7 84
rect -2 82 7 83
rect 9 82 18 84
rect -2 81 18 82
rect 14 74 18 81
rect 30 83 31 85
rect 33 83 34 85
rect 30 81 34 83
rect 62 85 66 90
rect 94 85 98 90
rect 62 83 63 85
rect 65 83 66 85
rect 62 81 66 83
rect 89 83 95 85
rect 97 83 98 85
rect 89 81 98 83
rect 14 72 15 74
rect 17 72 18 74
rect 14 71 18 72
rect 89 73 93 81
rect 89 71 90 73
rect 92 71 93 73
rect 14 70 40 71
rect 14 68 36 70
rect 38 68 40 70
rect 14 67 40 68
rect 14 65 15 67
rect 17 65 18 67
rect 14 63 18 65
rect 89 66 93 71
rect 89 64 90 66
rect 92 64 93 66
rect 14 48 18 59
rect 89 62 93 64
rect 14 46 26 48
rect 14 44 23 46
rect 25 44 26 46
rect 22 36 26 44
rect 22 34 23 36
rect 25 34 26 36
rect 22 29 26 34
rect 46 55 72 56
rect 46 53 58 55
rect 60 53 68 55
rect 70 53 72 55
rect 46 52 72 53
rect 14 23 18 25
rect 14 21 15 23
rect 17 21 18 23
rect 46 25 50 52
rect 86 46 90 51
rect 86 44 87 46
rect 89 44 90 46
rect 86 36 90 44
rect 86 34 87 36
rect 89 34 90 36
rect 86 29 90 34
rect 46 23 47 25
rect 49 23 50 25
rect 14 16 18 21
rect 14 14 15 16
rect 17 14 18 16
rect 14 7 18 14
rect 46 17 50 23
rect 46 15 47 17
rect 49 15 50 17
rect 46 13 50 15
rect 78 17 82 19
rect 78 15 79 17
rect 81 15 82 17
rect 78 7 82 15
rect -2 6 34 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 5 34 6
rect 9 4 31 5
rect 1 3 31 4
rect 33 3 34 5
rect 62 6 98 7
rect 62 5 71 6
rect 62 3 63 5
rect 65 4 71 5
rect 73 5 98 6
rect 73 4 95 5
rect 65 3 95 4
rect 97 3 98 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 -2 66 3
rect 94 -2 98 3
<< alu2 >>
rect -2 85 98 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 95 85
rect 97 83 98 85
rect -2 80 98 83
rect -2 5 98 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 95 5
rect 97 3 98 5
rect -2 -2 98 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
rect 93 5 99 7
rect 93 3 95 5
rect 97 3 99 5
rect 93 0 99 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
rect 93 85 99 88
rect 93 83 95 85
rect 97 83 99 85
rect 93 81 99 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polyct0 >>
rect 23 82 25 84
rect 71 82 73 84
rect 39 44 41 46
rect 55 44 57 46
rect 39 34 41 36
rect 55 34 57 36
rect 52 4 54 6
<< polyct1 >>
rect 7 82 9 84
rect 23 44 25 46
rect 87 44 89 46
rect 23 34 25 36
rect 87 34 89 36
rect 7 4 9 6
rect 71 4 73 6
<< ndifct0 >>
rect 26 23 28 25
rect 26 15 28 17
rect 36 23 38 25
rect 36 15 38 17
rect 58 22 60 24
rect 58 15 60 17
rect 90 22 92 24
rect 90 15 92 17
<< ndifct1 >>
rect 15 21 17 23
rect 15 14 17 16
rect 47 23 49 25
rect 47 15 49 17
rect 79 15 81 17
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< pdifct0 >>
rect 26 60 28 62
rect 26 53 28 55
rect 79 60 81 62
rect 79 53 81 55
<< pdifct1 >>
rect 15 72 17 74
rect 15 65 17 67
rect 36 68 38 70
rect 58 53 60 55
rect 68 53 70 55
rect 90 71 92 73
rect 90 64 92 66
<< alu0 >>
rect 21 84 27 85
rect 21 82 23 84
rect 25 82 27 84
rect 21 78 27 82
rect 69 84 75 85
rect 69 82 71 84
rect 73 82 75 84
rect 69 78 75 82
rect 21 74 75 78
rect 25 62 29 64
rect 25 60 26 62
rect 28 60 29 62
rect 25 55 29 60
rect 38 62 82 64
rect 38 60 79 62
rect 81 60 82 62
rect 25 53 26 55
rect 28 53 34 55
rect 25 51 34 53
rect 30 26 34 51
rect 38 46 42 60
rect 38 44 39 46
rect 41 44 42 46
rect 38 36 42 44
rect 38 34 39 36
rect 41 34 42 36
rect 38 32 42 34
rect 78 55 82 60
rect 78 53 79 55
rect 81 53 82 55
rect 24 25 40 26
rect 24 23 26 25
rect 28 23 36 25
rect 38 23 40 25
rect 24 22 40 23
rect 54 46 58 48
rect 54 44 55 46
rect 57 44 58 46
rect 54 36 58 44
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 78 26 82 53
rect 30 18 34 22
rect 24 17 42 18
rect 24 15 26 17
rect 28 15 36 17
rect 38 15 42 17
rect 24 14 42 15
rect 38 7 42 14
rect 57 24 93 26
rect 57 22 58 24
rect 60 22 90 24
rect 92 22 93 24
rect 57 17 61 22
rect 57 15 58 17
rect 60 15 61 17
rect 57 13 61 15
rect 89 17 93 22
rect 89 15 90 17
rect 92 15 93 17
rect 89 13 93 15
rect 38 6 56 7
rect 38 4 52 6
rect 54 4 56 6
rect 38 3 56 4
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< labels >>
rlabel alu1 16 52 16 52 6 b
rlabel alu1 24 36 24 36 6 b
rlabel alu1 48 32 48 32 6 z
rlabel alu1 88 40 88 40 6 a
rlabel alu2 48 4 48 4 6 vss
rlabel alu2 48 84 48 84 6 vdd
<< end >>
