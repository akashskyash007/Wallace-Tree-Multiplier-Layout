magic
tech scmos
timestamp 1199202469
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 19 68 53 70
rect 9 60 11 65
rect 19 60 21 68
rect 29 60 31 64
rect 40 60 42 64
rect 51 56 53 68
rect 51 42 53 46
rect 50 40 56 42
rect 50 38 52 40
rect 54 38 56 40
rect 9 35 11 38
rect 2 33 12 35
rect 19 33 21 38
rect 29 35 31 38
rect 25 33 32 35
rect 2 31 4 33
rect 6 31 12 33
rect 2 29 12 31
rect 10 26 12 29
rect 25 31 28 33
rect 30 31 32 33
rect 25 29 32 31
rect 40 32 42 38
rect 50 36 56 38
rect 40 30 46 32
rect 25 27 27 29
rect 21 25 27 27
rect 40 28 42 30
rect 44 28 46 30
rect 40 26 46 28
rect 53 26 55 36
rect 21 21 23 25
rect 31 21 33 25
rect 41 23 43 26
rect 10 11 12 15
rect 21 5 23 10
rect 31 4 33 10
rect 41 8 43 12
rect 53 4 55 19
rect 31 2 55 4
<< ndif >>
rect 2 19 10 26
rect 2 17 4 19
rect 6 17 10 19
rect 2 15 10 17
rect 12 21 17 26
rect 48 23 53 26
rect 36 21 41 23
rect 12 18 21 21
rect 12 16 16 18
rect 18 16 21 18
rect 12 15 21 16
rect 14 14 21 15
rect 16 10 21 14
rect 23 19 31 21
rect 23 17 26 19
rect 28 17 31 19
rect 23 10 31 17
rect 33 19 41 21
rect 33 17 36 19
rect 38 17 41 19
rect 33 12 41 17
rect 43 19 53 23
rect 55 24 62 26
rect 55 22 58 24
rect 60 22 62 24
rect 55 19 62 22
rect 43 12 51 19
rect 33 10 38 12
rect 45 10 51 12
rect 45 8 47 10
rect 49 8 51 10
rect 45 6 51 8
<< pdif >>
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 38 9 56
rect 11 42 19 60
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 57 29 60
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 42 40 60
rect 31 40 35 42
rect 37 40 40 42
rect 31 38 40 40
rect 42 58 49 60
rect 42 56 45 58
rect 47 56 49 58
rect 42 46 51 56
rect 53 52 58 56
rect 53 50 60 52
rect 53 48 56 50
rect 58 48 60 50
rect 53 46 60 48
rect 42 38 48 46
<< alu1 >>
rect -2 67 66 72
rect -2 65 57 67
rect 59 65 66 67
rect -2 64 66 65
rect 10 51 14 59
rect 2 47 14 51
rect 20 57 31 58
rect 20 55 24 57
rect 26 55 31 57
rect 20 54 31 55
rect 2 33 7 47
rect 2 31 4 33
rect 6 31 7 33
rect 2 29 7 31
rect 20 35 24 54
rect 18 29 24 35
rect 20 26 24 29
rect 20 22 31 26
rect 25 19 31 22
rect 25 17 26 19
rect 28 17 31 19
rect 25 14 31 17
rect 41 40 55 42
rect 41 38 52 40
rect 54 38 55 40
rect 50 36 55 38
rect 41 30 46 32
rect 41 28 42 30
rect 44 28 46 30
rect 50 29 54 36
rect 41 26 46 28
rect 42 18 46 26
rect 42 14 55 18
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 55 67 61 69
rect 55 65 57 67
rect 59 65 61 67
rect 55 63 61 65
<< nmos >>
rect 10 15 12 26
rect 21 10 23 21
rect 31 10 33 21
rect 41 12 43 23
rect 53 19 55 26
<< pmos >>
rect 9 38 11 60
rect 19 38 21 60
rect 29 38 31 60
rect 40 38 42 60
rect 51 46 53 56
<< polyct0 >>
rect 28 31 30 33
<< polyct1 >>
rect 52 38 54 40
rect 4 31 6 33
rect 42 28 44 30
<< ndifct0 >>
rect 4 17 6 19
rect 16 16 18 18
rect 36 17 38 19
rect 58 22 60 24
rect 47 8 49 10
<< ndifct1 >>
rect 26 17 28 19
<< ntiect1 >>
rect 57 65 59 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 4 56 6 58
rect 14 40 16 42
rect 35 40 37 42
rect 45 56 47 58
rect 56 48 58 50
<< pdifct1 >>
rect 24 55 26 57
<< alu0 >>
rect 3 58 7 64
rect 3 56 4 58
rect 6 56 7 58
rect 3 54 7 56
rect 43 58 49 64
rect 43 56 45 58
rect 47 56 49 58
rect 43 55 49 56
rect 11 42 17 44
rect 11 40 14 42
rect 16 40 17 42
rect 11 38 17 40
rect 3 19 7 21
rect 3 17 4 19
rect 6 17 7 19
rect 3 8 7 17
rect 11 19 15 38
rect 27 50 62 51
rect 27 48 56 50
rect 58 48 62 50
rect 27 47 62 48
rect 27 33 31 47
rect 27 31 28 33
rect 30 31 31 33
rect 27 29 31 31
rect 34 42 38 44
rect 34 40 35 42
rect 37 40 38 42
rect 11 18 20 19
rect 11 16 16 18
rect 18 16 20 18
rect 11 15 20 16
rect 34 21 38 40
rect 34 19 39 21
rect 34 17 36 19
rect 38 17 39 19
rect 34 15 39 17
rect 58 25 62 47
rect 56 24 62 25
rect 56 22 58 24
rect 60 22 62 24
rect 56 21 62 22
rect 45 10 51 11
rect 45 8 47 10
rect 49 8 51 10
<< labels >>
rlabel alu0 15 17 15 17 6 a0n
rlabel alu0 14 41 14 41 6 a0n
rlabel alu0 36 29 36 29 6 a1n
rlabel alu0 29 40 29 40 6 sn
rlabel alu0 44 49 44 49 6 sn
rlabel alu0 60 36 60 36 6 sn
rlabel alu1 4 40 4 40 6 a0
rlabel alu1 12 56 12 56 6 a0
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 32 20 32 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 44 24 44 24 6 a1
rlabel alu1 44 40 44 40 6 s
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 16 52 16 6 a1
rlabel alu1 52 36 52 36 6 s
<< end >>
