magic
tech scmos
timestamp 1199542018
<< ab >>
rect 0 0 160 100
<< nwell >>
rect -5 48 165 105
<< pwell >>
rect -5 -5 165 48
<< poly >>
rect 13 94 15 98
rect 145 94 147 98
rect 25 83 27 87
rect 37 84 39 88
rect 73 78 75 82
rect 85 78 87 82
rect 61 72 63 76
rect 13 41 15 55
rect 25 53 27 65
rect 37 63 39 66
rect 37 61 43 63
rect 37 59 39 61
rect 41 59 43 61
rect 37 57 43 59
rect 97 77 99 81
rect 109 77 111 81
rect 121 78 123 82
rect 19 51 27 53
rect 61 53 63 56
rect 73 53 75 56
rect 61 51 75 53
rect 85 53 87 56
rect 85 51 93 53
rect 19 49 21 51
rect 23 49 27 51
rect 19 47 27 49
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 87 49 89 51
rect 91 49 93 51
rect 87 47 93 49
rect 27 41 33 43
rect 13 39 29 41
rect 31 39 33 41
rect 13 25 15 39
rect 27 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 53 41 59 43
rect 97 41 99 55
rect 109 43 111 55
rect 121 53 123 56
rect 117 51 123 53
rect 117 49 119 51
rect 121 49 123 51
rect 117 47 123 49
rect 145 43 147 55
rect 53 39 55 41
rect 57 39 99 41
rect 53 37 59 39
rect 19 31 27 33
rect 19 29 21 31
rect 23 29 27 31
rect 37 29 39 37
rect 87 33 93 35
rect 67 31 73 33
rect 87 31 89 33
rect 91 31 93 33
rect 67 29 69 31
rect 71 29 73 31
rect 85 29 93 31
rect 19 27 27 29
rect 25 24 27 27
rect 61 27 75 29
rect 61 24 63 27
rect 73 24 75 27
rect 85 26 87 29
rect 97 27 99 39
rect 107 41 113 43
rect 127 41 133 43
rect 107 39 109 41
rect 111 39 129 41
rect 131 39 133 41
rect 107 37 113 39
rect 127 37 133 39
rect 137 41 147 43
rect 137 39 139 41
rect 141 39 147 41
rect 137 37 147 39
rect 117 31 123 33
rect 117 29 119 31
rect 121 29 123 31
rect 109 27 123 29
rect 25 11 27 15
rect 37 11 39 15
rect 61 12 63 16
rect 109 24 111 27
rect 121 24 123 27
rect 145 25 147 37
rect 73 11 75 15
rect 85 11 87 15
rect 97 11 99 15
rect 109 11 111 15
rect 121 12 123 16
rect 13 2 15 6
rect 145 2 147 6
<< ndif >>
rect 5 21 13 25
rect 5 19 7 21
rect 9 19 13 21
rect 5 6 13 19
rect 15 24 20 25
rect 29 24 37 29
rect 15 15 25 24
rect 27 15 37 24
rect 39 21 47 29
rect 92 26 97 27
rect 77 24 85 26
rect 39 19 43 21
rect 45 19 47 21
rect 39 15 47 19
rect 53 21 61 24
rect 53 19 55 21
rect 57 19 61 21
rect 53 17 61 19
rect 56 16 61 17
rect 63 16 73 24
rect 15 11 23 15
rect 65 15 73 16
rect 75 15 85 24
rect 87 23 97 26
rect 87 21 91 23
rect 93 21 97 23
rect 87 15 97 21
rect 99 24 107 27
rect 125 31 133 33
rect 125 29 129 31
rect 131 29 133 31
rect 125 27 133 29
rect 125 24 131 27
rect 99 15 109 24
rect 111 16 121 24
rect 123 16 131 24
rect 140 21 145 25
rect 111 15 119 16
rect 65 11 71 15
rect 113 11 119 15
rect 15 9 19 11
rect 21 9 23 11
rect 65 9 67 11
rect 69 9 71 11
rect 113 9 115 11
rect 117 9 119 11
rect 15 6 23 9
rect 65 7 71 9
rect 113 7 119 9
rect 137 11 145 21
rect 137 9 139 11
rect 141 9 145 11
rect 137 6 145 9
rect 147 21 155 25
rect 147 19 151 21
rect 153 19 155 21
rect 147 6 155 19
<< pdif >>
rect 5 81 13 94
rect 5 79 7 81
rect 9 79 13 81
rect 5 71 13 79
rect 5 69 7 71
rect 9 69 13 71
rect 5 61 13 69
rect 5 59 7 61
rect 9 59 13 61
rect 5 55 13 59
rect 15 91 23 94
rect 15 89 19 91
rect 21 89 23 91
rect 15 83 23 89
rect 41 91 47 93
rect 41 89 43 91
rect 45 89 47 91
rect 41 84 47 89
rect 65 91 71 93
rect 113 91 119 93
rect 65 89 67 91
rect 69 89 71 91
rect 29 83 37 84
rect 15 65 25 83
rect 27 71 37 83
rect 27 69 31 71
rect 33 69 37 71
rect 27 66 37 69
rect 39 66 47 84
rect 65 78 71 89
rect 113 89 115 91
rect 117 89 119 91
rect 65 72 73 78
rect 27 65 32 66
rect 15 55 23 65
rect 53 61 61 72
rect 53 59 55 61
rect 57 59 61 61
rect 53 56 61 59
rect 63 56 73 72
rect 75 71 85 78
rect 75 69 79 71
rect 81 69 85 71
rect 75 56 85 69
rect 87 77 95 78
rect 113 78 119 89
rect 137 91 145 94
rect 137 89 139 91
rect 141 89 145 91
rect 137 81 145 89
rect 137 79 139 81
rect 141 79 145 81
rect 113 77 121 78
rect 87 61 97 77
rect 87 59 91 61
rect 93 59 97 61
rect 87 56 97 59
rect 92 55 97 56
rect 99 71 109 77
rect 99 69 103 71
rect 105 69 109 71
rect 99 61 109 69
rect 99 59 103 61
rect 105 59 109 61
rect 99 55 109 59
rect 111 56 121 77
rect 123 61 131 78
rect 137 71 145 79
rect 137 69 139 71
rect 141 69 145 71
rect 137 67 145 69
rect 123 59 133 61
rect 123 57 129 59
rect 131 57 133 59
rect 123 56 133 57
rect 111 55 116 56
rect 127 55 133 56
rect 140 55 145 67
rect 147 81 155 94
rect 147 79 151 81
rect 153 79 155 81
rect 147 71 155 79
rect 147 69 151 71
rect 153 69 155 71
rect 147 61 155 69
rect 147 59 151 61
rect 153 59 155 61
rect 147 55 155 59
<< alu1 >>
rect -2 95 162 100
rect -2 93 55 95
rect 57 93 79 95
rect 81 93 91 95
rect 93 93 103 95
rect 105 93 127 95
rect 129 93 162 95
rect -2 91 162 93
rect -2 89 19 91
rect 21 89 43 91
rect 45 89 67 91
rect 69 89 115 91
rect 117 89 139 91
rect 141 89 162 91
rect -2 88 162 89
rect 8 82 12 83
rect 5 81 12 82
rect 5 79 7 81
rect 9 79 12 81
rect 5 78 12 79
rect 8 72 12 78
rect 5 71 12 72
rect 5 69 7 71
rect 9 69 12 71
rect 5 68 12 69
rect 8 62 12 68
rect 5 61 12 62
rect 5 59 7 61
rect 9 59 12 61
rect 5 58 12 59
rect 8 22 12 58
rect 5 21 12 22
rect 5 19 7 21
rect 9 19 12 21
rect 5 18 12 19
rect 8 17 12 18
rect 18 82 22 83
rect 18 78 122 82
rect 18 52 22 78
rect 68 72 72 73
rect 102 72 106 73
rect 29 71 35 72
rect 29 69 31 71
rect 33 69 35 71
rect 29 68 35 69
rect 40 68 72 72
rect 77 71 106 72
rect 77 69 79 71
rect 81 69 103 71
rect 105 69 106 71
rect 77 68 106 69
rect 18 51 25 52
rect 18 49 21 51
rect 23 49 25 51
rect 18 48 25 49
rect 18 32 22 48
rect 29 42 33 68
rect 40 63 44 68
rect 27 41 33 42
rect 27 39 29 41
rect 31 39 33 41
rect 27 38 33 39
rect 18 31 25 32
rect 18 29 21 31
rect 23 29 25 31
rect 18 28 25 29
rect 18 17 22 28
rect 29 22 33 38
rect 38 61 44 63
rect 38 59 39 61
rect 41 59 44 61
rect 38 58 44 59
rect 54 61 58 63
rect 54 59 55 61
rect 57 59 58 61
rect 38 41 42 58
rect 38 39 39 41
rect 41 39 42 41
rect 38 37 42 39
rect 54 41 58 59
rect 54 39 55 41
rect 57 39 58 41
rect 29 21 47 22
rect 29 19 43 21
rect 45 19 47 21
rect 29 18 47 19
rect 54 21 58 39
rect 54 19 55 21
rect 57 19 58 21
rect 54 17 58 19
rect 68 51 72 68
rect 68 49 69 51
rect 71 49 72 51
rect 68 31 72 49
rect 68 29 69 31
rect 71 29 72 31
rect 68 17 72 29
rect 78 61 95 62
rect 78 59 91 61
rect 93 59 95 61
rect 78 58 95 59
rect 102 61 106 68
rect 102 59 103 61
rect 105 59 106 61
rect 78 22 82 58
rect 102 57 106 59
rect 118 52 122 78
rect 138 81 142 88
rect 138 79 139 81
rect 141 79 142 81
rect 138 71 142 79
rect 138 69 139 71
rect 141 69 142 71
rect 138 67 142 69
rect 148 82 152 83
rect 148 81 155 82
rect 148 79 151 81
rect 153 79 155 81
rect 148 78 155 79
rect 148 72 152 78
rect 148 71 155 72
rect 148 69 151 71
rect 153 69 155 71
rect 148 68 155 69
rect 148 62 152 68
rect 148 61 155 62
rect 87 51 122 52
rect 87 49 89 51
rect 91 49 119 51
rect 121 49 122 51
rect 87 48 122 49
rect 98 41 113 42
rect 98 39 109 41
rect 111 39 113 41
rect 98 38 113 39
rect 98 34 102 38
rect 87 33 102 34
rect 87 31 89 33
rect 91 31 102 33
rect 87 30 102 31
rect 118 31 122 48
rect 118 29 119 31
rect 121 29 122 31
rect 118 27 122 29
rect 128 59 132 61
rect 128 57 129 59
rect 131 57 132 59
rect 128 41 132 57
rect 148 59 151 61
rect 153 59 155 61
rect 148 58 155 59
rect 128 39 129 41
rect 131 39 132 41
rect 128 31 132 39
rect 128 29 129 31
rect 131 29 132 31
rect 128 27 132 29
rect 138 41 142 43
rect 138 39 139 41
rect 141 39 142 41
rect 89 23 95 24
rect 89 22 91 23
rect 78 21 91 22
rect 93 22 95 23
rect 138 22 142 39
rect 93 21 142 22
rect 78 18 142 21
rect 148 22 152 58
rect 148 21 155 22
rect 148 19 151 21
rect 153 19 155 21
rect 148 18 155 19
rect 148 17 152 18
rect -2 11 162 12
rect -2 9 19 11
rect 21 9 67 11
rect 69 9 115 11
rect 117 9 139 11
rect 141 9 162 11
rect -2 7 162 9
rect -2 5 31 7
rect 33 5 43 7
rect 45 5 55 7
rect 57 5 79 7
rect 81 5 91 7
rect 93 5 103 7
rect 105 5 162 7
rect -2 0 162 5
<< ptie >>
rect 29 7 59 9
rect 77 7 107 9
rect 29 5 31 7
rect 33 5 43 7
rect 45 5 55 7
rect 57 5 59 7
rect 29 3 59 5
rect 77 5 79 7
rect 81 5 91 7
rect 93 5 103 7
rect 105 5 107 7
rect 77 3 107 5
<< ntie >>
rect 53 95 59 97
rect 53 93 55 95
rect 57 93 59 95
rect 77 95 107 97
rect 77 93 79 95
rect 81 93 91 95
rect 93 93 103 95
rect 105 93 107 95
rect 125 95 131 97
rect 125 93 127 95
rect 129 93 131 95
rect 53 86 59 93
rect 77 91 107 93
rect 125 86 131 93
<< nmos >>
rect 13 6 15 25
rect 25 15 27 24
rect 37 15 39 29
rect 61 16 63 24
rect 73 15 75 24
rect 85 15 87 26
rect 97 15 99 27
rect 109 15 111 24
rect 121 16 123 24
rect 145 6 147 25
<< pmos >>
rect 13 55 15 94
rect 25 65 27 83
rect 37 66 39 84
rect 61 56 63 72
rect 73 56 75 78
rect 85 56 87 78
rect 97 55 99 77
rect 109 55 111 77
rect 121 56 123 78
rect 145 55 147 94
<< polyct1 >>
rect 39 59 41 61
rect 21 49 23 51
rect 69 49 71 51
rect 89 49 91 51
rect 29 39 31 41
rect 39 39 41 41
rect 119 49 121 51
rect 55 39 57 41
rect 21 29 23 31
rect 89 31 91 33
rect 69 29 71 31
rect 109 39 111 41
rect 129 39 131 41
rect 139 39 141 41
rect 119 29 121 31
<< ndifct1 >>
rect 7 19 9 21
rect 43 19 45 21
rect 55 19 57 21
rect 91 21 93 23
rect 129 29 131 31
rect 19 9 21 11
rect 67 9 69 11
rect 115 9 117 11
rect 139 9 141 11
rect 151 19 153 21
<< ntiect1 >>
rect 55 93 57 95
rect 79 93 81 95
rect 91 93 93 95
rect 103 93 105 95
rect 127 93 129 95
<< ptiect1 >>
rect 31 5 33 7
rect 43 5 45 7
rect 55 5 57 7
rect 79 5 81 7
rect 91 5 93 7
rect 103 5 105 7
<< pdifct1 >>
rect 7 79 9 81
rect 7 69 9 71
rect 7 59 9 61
rect 19 89 21 91
rect 43 89 45 91
rect 67 89 69 91
rect 31 69 33 71
rect 115 89 117 91
rect 55 59 57 61
rect 79 69 81 71
rect 139 89 141 91
rect 139 79 141 81
rect 91 59 93 61
rect 103 69 105 71
rect 103 59 105 61
rect 139 69 141 71
rect 129 57 131 59
rect 151 79 153 81
rect 151 69 153 71
rect 151 59 153 61
<< labels >>
rlabel alu1 10 50 10 50 6 cout
rlabel alu1 20 50 20 50 6 a
rlabel polyct1 40 40 40 40 6 b
rlabel alu1 70 45 70 45 6 b
rlabel alu1 40 50 40 50 6 b
rlabel polyct1 40 60 40 60 6 b
rlabel alu1 50 70 50 70 6 b
rlabel alu1 60 70 60 70 6 b
rlabel ptiect1 80 6 80 6 6 vss
rlabel ntiect1 80 94 80 94 6 vdd
rlabel alu1 150 50 150 50 6 sout
<< end >>
