magic
tech scmos
timestamp 1199202079
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 24 39
rect 9 35 13 37
rect 15 35 20 37
rect 22 35 24 37
rect 9 33 24 35
rect 29 37 41 39
rect 29 35 37 37
rect 39 35 41 37
rect 29 33 41 35
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 33
rect 9 11 11 16
rect 19 11 21 16
rect 39 15 41 20
rect 29 7 31 12
<< ndif >>
rect 2 20 9 30
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 16 19 19
rect 21 20 29 30
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 23 12 29 16
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 20 39 26
rect 41 24 48 30
rect 41 22 44 24
rect 46 22 48 24
rect 41 20 48 22
rect 31 12 36 20
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 53 39 70
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 68 48 70
rect 41 66 44 68
rect 46 66 48 68
rect 41 61 48 66
rect 41 59 44 61
rect 46 59 48 61
rect 41 42 48 59
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 55 17 59
rect 2 54 17 55
rect 2 52 14 54
rect 16 52 23 54
rect 2 50 23 52
rect 2 30 6 50
rect 42 38 46 55
rect 33 37 46 38
rect 33 35 37 37
rect 39 35 46 37
rect 33 34 46 35
rect 2 28 17 30
rect 2 26 14 28
rect 16 26 17 28
rect 2 25 17 26
rect 13 21 17 25
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 12 31 30
rect 39 20 41 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
<< polyct0 >>
rect 13 35 15 37
rect 20 35 22 37
<< polyct1 >>
rect 37 35 39 37
<< ndifct0 >>
rect 4 18 6 20
rect 24 18 26 20
rect 34 26 36 28
rect 44 22 46 24
<< ndifct1 >>
rect 14 26 16 28
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 24 66 26 68
rect 24 59 26 61
rect 34 51 36 53
rect 34 44 36 46
rect 44 66 46 68
rect 44 59 46 61
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 23 66 24 68
rect 26 66 27 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 23 61 27 66
rect 23 59 24 61
rect 26 59 27 61
rect 23 57 27 59
rect 42 66 44 68
rect 46 66 48 68
rect 42 61 48 66
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 33 53 37 55
rect 33 51 34 53
rect 36 51 37 53
rect 33 46 37 51
rect 23 44 34 46
rect 36 44 37 46
rect 23 42 37 44
rect 23 38 27 42
rect 11 37 27 38
rect 11 35 13 37
rect 15 35 20 37
rect 22 35 27 37
rect 11 34 27 35
rect 23 29 27 34
rect 23 28 38 29
rect 23 26 34 28
rect 36 26 38 28
rect 23 25 38 26
rect 43 24 47 26
rect 43 22 44 24
rect 46 22 47 24
rect 2 20 8 21
rect 2 18 4 20
rect 6 18 8 20
rect 2 12 8 18
rect 22 20 28 21
rect 22 18 24 20
rect 26 18 28 20
rect 22 12 28 18
rect 43 12 47 22
<< labels >>
rlabel alu0 19 36 19 36 6 an
rlabel alu0 30 27 30 27 6 an
rlabel alu0 35 48 35 48 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 36 36 36 6 a
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 48 44 48 6 a
<< end >>
