magic
tech scmos
timestamp 1199201640
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 61 11 65
rect 19 63 21 68
rect 29 63 31 68
rect 9 39 11 43
rect 19 39 21 50
rect 29 47 31 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 28 11 33
rect 22 28 24 33
rect 29 28 31 41
rect 9 15 11 19
rect 22 12 24 17
rect 29 12 31 17
<< ndif >>
rect 4 25 9 28
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 19 22 28
rect 13 17 22 19
rect 24 17 29 28
rect 31 23 36 28
rect 31 21 38 23
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
rect 13 11 20 17
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 13 61 19 63
rect 4 56 9 61
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 59 19 61
rect 11 57 14 59
rect 16 57 19 59
rect 11 50 19 57
rect 21 61 29 63
rect 21 59 24 61
rect 26 59 29 61
rect 21 54 29 59
rect 21 52 24 54
rect 26 52 29 54
rect 21 50 29 52
rect 31 61 38 63
rect 31 59 34 61
rect 36 59 38 61
rect 31 50 38 59
rect 11 43 17 50
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 54 7 56
rect 2 52 4 54
rect 6 52 7 54
rect 2 47 7 52
rect 2 45 4 47
rect 6 45 7 47
rect 2 43 7 45
rect 2 23 6 43
rect 34 46 38 55
rect 25 45 38 46
rect 25 43 31 45
rect 33 43 38 45
rect 25 42 38 43
rect 17 37 31 38
rect 17 35 21 37
rect 23 35 31 37
rect 17 34 31 35
rect 2 21 4 23
rect 6 21 14 23
rect 2 17 14 21
rect 26 25 31 34
rect -2 11 42 12
rect -2 9 15 11
rect 17 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 19 11 28
rect 22 17 24 28
rect 29 17 31 28
<< pmos >>
rect 9 43 11 61
rect 19 50 21 63
rect 29 50 31 63
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 21 35 23 37
<< ndifct0 >>
rect 34 19 36 21
<< ndifct1 >>
rect 4 21 6 23
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 57 16 59
rect 24 59 26 61
rect 24 52 26 54
rect 34 59 36 61
<< pdifct1 >>
rect 4 52 6 54
rect 4 45 6 47
<< alu0 >>
rect 12 59 18 68
rect 12 57 14 59
rect 16 57 18 59
rect 12 56 18 57
rect 23 61 27 63
rect 23 59 24 61
rect 26 59 27 61
rect 23 54 27 59
rect 32 61 38 68
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 23 53 24 54
rect 10 52 24 53
rect 26 52 27 54
rect 10 49 27 52
rect 10 37 14 49
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 10 26 22 30
rect 6 23 7 25
rect 18 22 22 26
rect 18 21 38 22
rect 18 19 34 21
rect 36 19 38 21
rect 18 18 38 19
<< labels >>
rlabel alu0 12 39 12 39 6 zn
rlabel alu0 25 56 25 56 6 zn
rlabel alu0 28 20 28 20 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 52 36 52 6 b
<< end >>
