magic
tech scmos
timestamp 1199202811
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 10 72 62 74
rect 10 63 12 72
rect 20 63 22 68
rect 30 63 32 68
rect 40 63 42 68
rect 50 63 52 68
rect 60 63 62 72
rect 10 35 12 43
rect 20 39 22 43
rect 30 39 32 43
rect 40 39 42 43
rect 50 39 52 43
rect 60 39 62 43
rect 20 37 26 39
rect 20 35 22 37
rect 24 35 26 37
rect 10 33 16 35
rect 20 33 26 35
rect 30 37 42 39
rect 30 35 35 37
rect 37 35 42 37
rect 30 33 42 35
rect 46 37 52 39
rect 46 35 48 37
rect 50 35 52 37
rect 46 33 52 35
rect 56 37 63 39
rect 56 35 59 37
rect 61 35 63 37
rect 56 33 63 35
rect 14 30 16 33
rect 22 30 24 33
rect 30 30 32 33
rect 40 30 42 33
rect 48 30 50 33
rect 56 30 58 33
rect 14 6 16 10
rect 22 6 24 10
rect 30 6 32 10
rect 40 6 42 10
rect 48 6 50 10
rect 56 6 58 10
<< ndif >>
rect 6 14 14 30
rect 6 12 9 14
rect 11 12 14 14
rect 6 10 14 12
rect 16 10 22 30
rect 24 10 30 30
rect 32 21 40 30
rect 32 19 35 21
rect 37 19 40 21
rect 32 10 40 19
rect 42 10 48 30
rect 50 10 56 30
rect 58 21 66 30
rect 58 19 61 21
rect 63 19 66 21
rect 58 14 66 19
rect 58 12 61 14
rect 63 12 66 14
rect 58 10 66 12
<< pdif >>
rect 2 61 10 63
rect 2 59 4 61
rect 6 59 10 61
rect 2 54 10 59
rect 2 52 4 54
rect 6 52 10 54
rect 2 43 10 52
rect 12 61 20 63
rect 12 59 15 61
rect 17 59 20 61
rect 12 54 20 59
rect 12 52 15 54
rect 17 52 20 54
rect 12 43 20 52
rect 22 61 30 63
rect 22 59 25 61
rect 27 59 30 61
rect 22 43 30 59
rect 32 61 40 63
rect 32 59 35 61
rect 37 59 40 61
rect 32 54 40 59
rect 32 52 35 54
rect 37 52 40 54
rect 32 43 40 52
rect 42 61 50 63
rect 42 59 45 61
rect 47 59 50 61
rect 42 43 50 59
rect 52 61 60 63
rect 52 59 55 61
rect 57 59 60 61
rect 52 54 60 59
rect 52 52 55 54
rect 57 52 60 54
rect 52 43 60 52
rect 62 61 70 63
rect 62 59 66 61
rect 68 59 70 61
rect 62 43 70 59
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 14 61 18 63
rect 14 59 15 61
rect 17 59 18 61
rect 14 55 18 59
rect 34 61 38 63
rect 34 59 35 61
rect 37 59 38 61
rect 10 54 18 55
rect 34 54 38 59
rect 54 61 58 63
rect 54 59 55 61
rect 57 59 58 61
rect 54 54 58 59
rect 10 52 15 54
rect 17 52 35 54
rect 37 52 55 54
rect 57 52 58 54
rect 10 50 58 52
rect 10 22 14 50
rect 22 42 52 46
rect 22 39 26 42
rect 18 37 26 39
rect 18 35 22 37
rect 24 35 26 37
rect 18 33 26 35
rect 33 37 39 38
rect 33 35 35 37
rect 37 35 39 37
rect 33 30 39 35
rect 46 37 52 42
rect 66 39 70 55
rect 46 35 48 37
rect 50 35 52 37
rect 46 34 52 35
rect 58 37 70 39
rect 58 35 59 37
rect 61 35 70 37
rect 58 33 70 35
rect 33 26 47 30
rect 10 21 39 22
rect 10 19 35 21
rect 37 19 39 21
rect 10 18 39 19
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 14 10 16 30
rect 22 10 24 30
rect 30 10 32 30
rect 40 10 42 30
rect 48 10 50 30
rect 56 10 58 30
<< pmos >>
rect 10 43 12 63
rect 20 43 22 63
rect 30 43 32 63
rect 40 43 42 63
rect 50 43 52 63
rect 60 43 62 63
<< polyct1 >>
rect 22 35 24 37
rect 35 35 37 37
rect 48 35 50 37
rect 59 35 61 37
<< ndifct0 >>
rect 9 12 11 14
rect 61 19 63 21
rect 61 12 63 14
<< ndifct1 >>
rect 35 19 37 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 59 6 61
rect 4 52 6 54
rect 25 59 27 61
rect 45 59 47 61
rect 66 59 68 61
<< pdifct1 >>
rect 15 59 17 61
rect 15 52 17 54
rect 35 59 37 61
rect 35 52 37 54
rect 55 59 57 61
rect 55 52 57 54
<< alu0 >>
rect 3 61 7 68
rect 3 59 4 61
rect 6 59 7 61
rect 3 54 7 59
rect 23 61 29 68
rect 23 59 25 61
rect 27 59 29 61
rect 23 58 29 59
rect 3 52 4 54
rect 6 52 7 54
rect 3 50 7 52
rect 43 61 49 68
rect 43 59 45 61
rect 47 59 49 61
rect 43 58 49 59
rect 64 61 70 68
rect 64 59 66 61
rect 68 59 70 61
rect 64 58 70 59
rect 59 21 65 22
rect 59 19 61 21
rect 63 19 65 21
rect 7 14 13 15
rect 7 12 9 14
rect 11 12 13 14
rect 59 14 65 19
rect 59 12 61 14
rect 63 12 65 14
<< labels >>
rlabel alu1 12 40 12 40 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 36 20 36 6 b
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel ndifct1 36 20 36 20 6 z
rlabel alu1 36 32 36 32 6 c
rlabel alu1 44 28 44 28 6 c
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 44 36 44 6 b
rlabel alu1 36 56 36 56 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel polyct1 60 36 60 36 6 a
rlabel alu1 68 44 68 44 6 a
<< end >>
