magic
tech scmos
timestamp 1199202364
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 58 51 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 41 39
rect 22 35 37 37
rect 39 35 41 37
rect 22 33 41 35
rect 49 39 51 42
rect 49 37 55 39
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 22 30 24 33
rect 32 30 34 33
rect 22 9 24 14
rect 32 9 34 14
<< ndif >>
rect 14 26 22 30
rect 14 24 17 26
rect 19 24 22 26
rect 14 18 22 24
rect 14 16 17 18
rect 19 16 22 18
rect 14 14 22 16
rect 24 28 32 30
rect 24 26 27 28
rect 29 26 32 28
rect 24 21 32 26
rect 24 19 27 21
rect 29 19 32 21
rect 24 14 32 19
rect 34 26 42 30
rect 34 24 37 26
rect 39 24 42 26
rect 34 18 42 24
rect 34 16 37 18
rect 39 16 42 18
rect 34 14 42 16
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 53 39 70
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 58 47 70
rect 41 56 49 58
rect 41 54 44 56
rect 46 54 49 56
rect 41 42 49 54
rect 51 55 56 58
rect 51 53 58 55
rect 51 51 54 53
rect 56 51 58 53
rect 51 46 58 51
rect 51 44 54 46
rect 56 44 58 46
rect 51 42 58 44
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 33 53 38 55
rect 33 51 34 53
rect 36 51 38 53
rect 53 53 62 55
rect 33 46 38 51
rect 53 51 54 53
rect 56 51 62 53
rect 53 49 62 51
rect 53 46 57 49
rect 9 44 14 46
rect 16 44 34 46
rect 36 44 54 46
rect 56 44 57 46
rect 9 42 57 44
rect 26 28 30 42
rect 35 37 55 38
rect 35 35 37 37
rect 39 35 51 37
rect 53 35 55 37
rect 35 34 55 35
rect 26 26 27 28
rect 29 26 30 28
rect 26 21 30 26
rect 26 19 27 21
rect 29 19 30 21
rect 26 17 30 19
rect 49 26 55 34
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 22 14 24 30
rect 32 14 34 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 58
<< polyct1 >>
rect 37 35 39 37
rect 51 35 53 37
<< ndifct0 >>
rect 17 24 19 26
rect 17 16 19 18
rect 37 24 39 26
rect 37 16 39 18
<< ndifct1 >>
rect 27 26 29 28
rect 27 19 29 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 51 16 53
rect 24 66 26 68
rect 24 59 26 61
rect 44 54 46 56
<< pdifct1 >>
rect 14 44 16 46
rect 34 51 36 53
rect 34 44 36 46
rect 54 51 56 53
rect 54 44 56 46
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 43 56 47 68
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 13 46 17 51
rect 43 54 44 56
rect 46 54 47 56
rect 43 52 47 54
rect 16 26 20 28
rect 16 24 17 26
rect 19 24 20 26
rect 16 18 20 24
rect 16 16 17 18
rect 19 16 20 18
rect 36 26 40 28
rect 36 24 37 26
rect 39 24 40 26
rect 36 18 40 24
rect 16 12 20 16
rect 36 16 37 18
rect 39 16 40 18
rect 36 12 40 16
<< labels >>
rlabel alu1 12 44 12 44 6 z
rlabel alu1 28 32 28 32 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 36 44 36 6 a
rlabel alu1 44 44 44 44 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 32 52 32 6 a
rlabel alu1 52 44 52 44 6 z
rlabel alu1 60 52 60 52 6 z
<< end >>
