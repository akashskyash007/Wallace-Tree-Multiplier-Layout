magic
tech scmos
timestamp 1199202946
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 12 61 14 65
rect 19 61 21 66
rect 12 43 14 46
rect 9 41 15 43
rect 9 39 11 41
rect 13 39 15 41
rect 9 37 15 39
rect 19 40 21 46
rect 19 38 25 40
rect 10 26 12 37
rect 19 36 21 38
rect 23 36 25 38
rect 19 34 25 36
rect 20 26 22 34
rect 10 15 12 19
rect 20 15 22 19
<< ndif >>
rect 2 23 10 26
rect 2 21 4 23
rect 6 21 10 23
rect 2 19 10 21
rect 12 24 20 26
rect 12 22 15 24
rect 17 22 20 24
rect 12 19 20 22
rect 22 23 30 26
rect 22 21 26 23
rect 28 21 30 23
rect 22 19 30 21
<< pdif >>
rect 5 59 12 61
rect 5 57 7 59
rect 9 57 12 59
rect 5 55 12 57
rect 7 46 12 55
rect 14 46 19 61
rect 21 59 30 61
rect 21 57 26 59
rect 28 57 30 59
rect 21 46 30 57
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 60 6 63
rect 2 59 11 60
rect 2 57 7 59
rect 9 57 11 59
rect 2 56 11 57
rect 2 33 6 56
rect 18 47 22 55
rect 10 43 22 47
rect 10 41 14 43
rect 10 39 11 41
rect 13 39 14 41
rect 26 39 30 47
rect 10 37 14 39
rect 18 38 30 39
rect 18 36 21 38
rect 23 36 30 38
rect 18 33 30 36
rect 2 29 14 33
rect 10 25 14 29
rect 10 24 19 25
rect 10 22 15 24
rect 17 22 19 24
rect 10 21 19 22
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 10 19 12 26
rect 20 19 22 26
<< pmos >>
rect 12 46 14 61
rect 19 46 21 61
<< polyct1 >>
rect 11 39 13 41
rect 21 36 23 38
<< ndifct0 >>
rect 4 21 6 23
rect 26 21 28 23
<< ndifct1 >>
rect 15 22 17 24
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 26 57 28 59
<< pdifct1 >>
rect 7 57 9 59
<< alu0 >>
rect 25 59 29 68
rect 25 57 26 59
rect 28 57 29 59
rect 25 55 29 57
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 25 23 29 25
rect 25 21 26 23
rect 28 21 29 23
rect 3 12 7 21
rect 25 12 29 21
<< labels >>
rlabel alu1 4 48 4 48 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 44 12 44 6 b
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 20 52 20 52 6 b
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 40 28 40 6 a
<< end >>
