magic
tech scmos
timestamp 1199202664
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 10 61 12 66
rect 20 61 22 65
rect 10 40 12 43
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 20 36 22 43
rect 9 34 15 36
rect 19 34 30 36
rect 12 27 14 34
rect 19 32 26 34
rect 28 32 30 34
rect 19 30 30 32
rect 19 27 21 30
rect 12 15 14 19
rect 19 14 21 19
<< ndif >>
rect 5 25 12 27
rect 5 23 7 25
rect 9 23 12 25
rect 5 21 12 23
rect 7 19 12 21
rect 14 19 19 27
rect 21 19 30 27
rect 23 17 26 19
rect 28 17 30 19
rect 23 15 30 17
<< pdif >>
rect 2 61 8 63
rect 2 59 4 61
rect 6 59 10 61
rect 2 43 10 59
rect 12 59 20 61
rect 12 57 15 59
rect 17 57 20 59
rect 12 52 20 57
rect 12 50 15 52
rect 17 50 20 52
rect 12 43 20 50
rect 22 59 30 61
rect 22 57 26 59
rect 28 57 30 59
rect 22 52 30 57
rect 22 50 26 52
rect 28 50 30 52
rect 22 43 30 50
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 50 15 54
rect 2 26 6 50
rect 17 43 23 46
rect 10 39 23 43
rect 10 38 14 39
rect 10 36 11 38
rect 13 36 14 38
rect 10 33 14 36
rect 24 34 30 35
rect 24 32 26 34
rect 28 32 30 34
rect 24 31 30 32
rect 2 25 11 26
rect 2 23 7 25
rect 9 23 11 25
rect 2 22 11 23
rect 18 25 30 31
rect 18 17 22 25
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 12 19 14 27
rect 19 19 21 27
<< pmos >>
rect 10 43 12 61
rect 20 43 22 61
<< polyct1 >>
rect 11 36 13 38
rect 26 32 28 34
<< ndifct0 >>
rect 26 17 28 19
<< ndifct1 >>
rect 7 23 9 25
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 59 6 61
rect 15 57 17 59
rect 15 50 17 52
rect 26 57 28 59
rect 26 50 28 52
<< alu0 >>
rect 2 61 8 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 59 19 60
rect 13 57 15 59
rect 17 57 19 59
rect 13 54 19 57
rect 15 52 19 54
rect 17 50 19 52
rect 6 49 19 50
rect 24 59 30 68
rect 24 57 26 59
rect 28 57 30 59
rect 24 52 30 57
rect 24 50 26 52
rect 28 50 30 52
rect 24 49 30 50
rect 25 19 29 21
rect 25 17 26 19
rect 28 17 29 19
rect 25 12 29 17
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 36 12 36 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 24 20 24 6 a
rlabel alu1 20 44 20 44 6 b
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 28 28 28 6 a
<< end >>
