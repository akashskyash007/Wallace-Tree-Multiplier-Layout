magic
tech scmos
timestamp 1199543359
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -2 48 82 104
<< pwell >>
rect -2 -4 82 48
<< poly >>
rect 19 95 21 98
rect 27 95 29 98
rect 35 95 37 98
rect 43 95 45 98
rect 55 95 57 98
rect 67 95 69 98
rect 19 53 21 55
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 11 47 23 49
rect 11 25 13 47
rect 27 43 29 55
rect 35 53 37 55
rect 43 53 45 55
rect 55 53 57 55
rect 67 53 69 55
rect 35 51 39 53
rect 43 51 49 53
rect 55 51 69 53
rect 37 43 39 51
rect 47 43 49 51
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 23 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 23 25 25 37
rect 37 29 39 37
rect 47 29 49 37
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 33 27 39 29
rect 45 27 49 29
rect 55 27 69 29
rect 33 25 35 27
rect 45 25 47 27
rect 55 25 57 27
rect 67 25 69 27
rect 11 12 13 15
rect 23 12 25 15
rect 33 12 35 15
rect 45 12 47 15
rect 55 2 57 5
rect 67 2 69 5
<< ndif >>
rect 3 15 11 25
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 15 23 19
rect 25 15 33 25
rect 35 21 45 25
rect 35 19 39 21
rect 41 19 45 21
rect 35 15 45 19
rect 47 15 55 25
rect 3 11 9 15
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 27 9 31 15
rect 49 9 55 15
rect 27 7 33 9
rect 27 5 29 7
rect 31 5 33 7
rect 27 3 33 5
rect 47 7 55 9
rect 47 5 49 7
rect 51 5 55 7
rect 57 21 67 25
rect 57 19 61 21
rect 63 19 67 21
rect 57 5 67 19
rect 69 11 77 25
rect 69 9 73 11
rect 75 9 77 11
rect 69 5 77 9
rect 47 3 53 5
<< pdif >>
rect 11 85 19 95
rect 7 81 19 85
rect 7 79 9 81
rect 11 79 19 81
rect 7 71 19 79
rect 7 69 9 71
rect 11 69 19 71
rect 7 61 19 69
rect 7 59 9 61
rect 11 59 19 61
rect 7 55 19 59
rect 21 55 27 95
rect 29 55 35 95
rect 37 55 43 95
rect 45 91 55 95
rect 45 89 49 91
rect 51 89 55 91
rect 45 55 55 89
rect 57 81 67 95
rect 57 79 61 81
rect 63 79 67 81
rect 57 71 67 79
rect 57 69 61 71
rect 63 69 67 71
rect 57 61 67 69
rect 57 59 61 61
rect 63 59 67 61
rect 57 55 67 59
rect 69 91 77 95
rect 69 89 73 91
rect 75 89 77 91
rect 69 81 77 89
rect 69 79 73 81
rect 75 79 77 81
rect 69 71 77 79
rect 69 69 73 71
rect 75 69 77 71
rect 69 55 77 69
<< alu1 >>
rect -2 91 82 100
rect -2 89 49 91
rect 51 89 73 91
rect 75 89 82 91
rect -2 88 82 89
rect 8 81 12 82
rect 8 79 9 81
rect 11 79 12 81
rect 8 78 12 79
rect 9 72 11 78
rect 8 71 12 72
rect 8 69 9 71
rect 11 69 12 71
rect 8 68 12 69
rect 9 62 11 68
rect 8 61 12 62
rect 8 59 9 61
rect 11 59 12 61
rect 8 58 12 59
rect 9 22 11 58
rect 18 51 22 82
rect 18 49 19 51
rect 21 49 22 51
rect 18 28 22 49
rect 28 41 32 82
rect 28 39 29 41
rect 31 39 32 41
rect 28 28 32 39
rect 38 41 42 82
rect 38 39 39 41
rect 41 39 42 41
rect 38 28 42 39
rect 48 41 52 82
rect 58 81 64 82
rect 58 79 61 81
rect 63 79 64 81
rect 58 78 64 79
rect 72 81 76 88
rect 72 79 73 81
rect 75 79 76 81
rect 58 72 62 78
rect 58 71 64 72
rect 58 69 61 71
rect 63 69 64 71
rect 58 68 64 69
rect 72 71 76 79
rect 72 69 73 71
rect 75 69 76 71
rect 72 68 76 69
rect 58 62 62 68
rect 58 61 72 62
rect 58 59 61 61
rect 63 59 72 61
rect 58 58 72 59
rect 58 51 62 52
rect 58 49 59 51
rect 61 49 62 51
rect 58 48 62 49
rect 48 39 49 41
rect 51 39 52 41
rect 48 38 52 39
rect 59 32 61 48
rect 58 31 62 32
rect 49 29 59 31
rect 61 29 62 31
rect 49 22 51 29
rect 58 28 62 29
rect 68 22 72 58
rect 9 21 20 22
rect 38 21 51 22
rect 9 19 17 21
rect 19 19 39 21
rect 41 19 51 21
rect 9 18 20 19
rect 38 18 51 19
rect 60 21 72 22
rect 60 19 61 21
rect 63 19 72 21
rect 60 18 72 19
rect -2 11 82 12
rect -2 9 5 11
rect 7 9 73 11
rect 75 9 82 11
rect -2 7 82 9
rect -2 5 29 7
rect 31 5 49 7
rect 51 5 82 7
rect -2 0 82 5
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 33 15 35 25
rect 45 15 47 25
rect 55 5 57 25
rect 67 5 69 25
<< pmos >>
rect 19 55 21 95
rect 27 55 29 95
rect 35 55 37 95
rect 43 55 45 95
rect 55 55 57 95
rect 67 55 69 95
<< polyct1 >>
rect 19 49 21 51
rect 59 49 61 51
rect 29 39 31 41
rect 39 39 41 41
rect 49 39 51 41
rect 59 29 61 31
<< ndifct1 >>
rect 17 19 19 21
rect 39 19 41 21
rect 5 9 7 11
rect 29 5 31 7
rect 49 5 51 7
rect 61 19 63 21
rect 73 9 75 11
<< pdifct1 >>
rect 9 79 11 81
rect 9 69 11 71
rect 9 59 11 61
rect 49 89 51 91
rect 61 79 63 81
rect 61 69 63 71
rect 61 59 63 61
rect 73 89 75 91
rect 73 79 75 81
rect 73 69 75 71
<< labels >>
rlabel alu1 30 55 30 55 6 i0
rlabel alu1 20 55 20 55 6 i1
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 40 55 40 55 6 i2
rlabel alu1 50 60 50 60 6 i3
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 70 40 70 40 6 q
rlabel alu1 60 70 60 70 6 q
<< end >>
