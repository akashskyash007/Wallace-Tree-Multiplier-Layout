magic
tech scmos
timestamp 1635158097
<< ab >>
rect -39 5 1 77
rect -22 -67 2 5
rect 5 -67 45 77
rect 49 -67 73 77
<< nwell >>
rect -44 37 78 82
rect -27 -72 78 -27
<< pwell >>
rect -44 10 78 37
rect -27 -27 78 10
<< poly >>
rect -17 71 -15 75
rect -10 71 -8 75
rect -30 61 -28 66
rect 14 62 16 66
rect 24 64 26 69
rect 34 64 36 69
rect -30 40 -28 43
rect -17 40 -15 50
rect -10 47 -8 50
rect -10 45 -4 47
rect -10 43 -8 45
rect -6 43 -4 45
rect 58 61 60 66
rect -10 41 -4 43
rect -30 38 -24 40
rect -30 36 -28 38
rect -26 36 -24 38
rect -30 34 -24 36
rect -20 38 -14 40
rect -20 36 -18 38
rect -16 36 -14 38
rect -20 34 -14 36
rect -30 31 -28 34
rect -20 31 -18 34
rect -10 31 -8 41
rect 14 40 16 44
rect 24 40 26 51
rect 34 48 36 51
rect 34 46 40 48
rect 34 44 36 46
rect 38 44 40 46
rect 34 42 40 44
rect 14 38 20 40
rect 14 36 16 38
rect 18 36 20 38
rect 14 34 20 36
rect 24 38 30 40
rect 24 36 26 38
rect 28 36 30 38
rect 24 34 30 36
rect 14 29 16 34
rect 27 29 29 34
rect 34 29 36 42
rect 58 40 60 43
rect 58 38 64 40
rect 58 36 60 38
rect 62 36 64 38
rect 58 34 64 36
rect 58 31 60 34
rect -30 17 -28 22
rect -20 20 -18 25
rect -10 20 -8 25
rect 14 16 16 20
rect 27 13 29 18
rect 34 13 36 18
rect 58 17 60 22
rect -9 -12 -7 -7
rect 14 -10 16 -6
rect 27 -8 29 -3
rect 34 -8 36 -3
rect 58 -12 60 -7
rect -9 -24 -7 -21
rect -13 -26 -7 -24
rect -13 -28 -11 -26
rect -9 -28 -7 -26
rect -13 -30 -7 -28
rect -9 -33 -7 -30
rect 14 -24 16 -19
rect 27 -24 29 -19
rect 14 -26 20 -24
rect 14 -28 16 -26
rect 18 -28 20 -26
rect 14 -30 20 -28
rect 24 -26 30 -24
rect 24 -28 26 -26
rect 28 -28 30 -26
rect 24 -30 30 -28
rect 14 -34 16 -30
rect -9 -56 -7 -51
rect 24 -41 26 -30
rect 34 -32 36 -19
rect 58 -24 60 -21
rect 58 -26 64 -24
rect 58 -28 60 -26
rect 62 -28 64 -26
rect 58 -30 64 -28
rect 34 -34 40 -32
rect 58 -33 60 -30
rect 34 -36 36 -34
rect 38 -36 40 -34
rect 34 -38 40 -36
rect 34 -41 36 -38
rect 14 -56 16 -52
rect 24 -59 26 -54
rect 34 -59 36 -54
rect 58 -56 60 -51
<< ndif >>
rect -37 29 -30 31
rect -37 27 -35 29
rect -33 27 -30 29
rect -37 25 -30 27
rect -35 22 -30 25
rect -28 25 -20 31
rect -18 29 -10 31
rect -18 27 -15 29
rect -13 27 -10 29
rect -18 25 -10 27
rect -8 25 -1 31
rect 51 29 58 31
rect 9 26 14 29
rect -28 22 -22 25
rect -26 18 -22 22
rect -6 18 -1 25
rect 7 24 14 26
rect 7 22 9 24
rect 11 22 14 24
rect 7 20 14 22
rect 16 20 27 29
rect -26 16 -20 18
rect -26 14 -24 16
rect -22 14 -20 16
rect -26 12 -20 14
rect -7 16 -1 18
rect 18 18 27 20
rect 29 18 34 29
rect 36 24 41 29
rect 51 27 53 29
rect 55 27 58 29
rect 51 25 58 27
rect 36 22 43 24
rect 53 22 58 25
rect 60 26 71 31
rect 60 24 67 26
rect 69 24 71 26
rect 60 22 71 24
rect 36 20 39 22
rect 41 20 43 22
rect 36 18 43 20
rect -7 14 -5 16
rect -3 14 -1 16
rect -7 12 -1 14
rect 18 12 25 18
rect 18 10 20 12
rect 22 10 25 12
rect 18 8 25 10
rect 18 0 25 2
rect 18 -2 20 0
rect 22 -2 25 0
rect 18 -8 25 -2
rect 18 -10 27 -8
rect 7 -12 14 -10
rect -20 -14 -9 -12
rect -20 -16 -18 -14
rect -16 -16 -9 -14
rect -20 -21 -9 -16
rect -7 -15 -2 -12
rect 7 -14 9 -12
rect 11 -14 14 -12
rect -7 -17 0 -15
rect 7 -16 14 -14
rect -7 -19 -4 -17
rect -2 -19 0 -17
rect 9 -19 14 -16
rect 16 -19 27 -10
rect 29 -19 34 -8
rect 36 -10 43 -8
rect 36 -12 39 -10
rect 41 -12 43 -10
rect 36 -14 43 -12
rect 36 -19 41 -14
rect 53 -15 58 -12
rect 51 -17 58 -15
rect 51 -19 53 -17
rect 55 -19 58 -17
rect -7 -21 0 -19
rect 51 -21 58 -19
rect 60 -14 71 -12
rect 60 -16 67 -14
rect 69 -16 71 -14
rect 60 -21 71 -16
<< pdif >>
rect -26 69 -17 71
rect -26 67 -24 69
rect -22 67 -17 69
rect -26 61 -17 67
rect -37 59 -30 61
rect -37 57 -35 59
rect -33 57 -30 59
rect -37 52 -30 57
rect -37 50 -35 52
rect -33 50 -30 52
rect -37 48 -30 50
rect -35 43 -30 48
rect -28 50 -17 61
rect -15 50 -10 71
rect -8 64 -3 71
rect -8 62 -1 64
rect 18 62 24 64
rect -8 60 -5 62
rect -3 60 -1 62
rect -8 58 -1 60
rect -8 50 -3 58
rect 9 57 14 62
rect 7 55 14 57
rect 7 53 9 55
rect 11 53 14 55
rect -28 43 -20 50
rect 7 48 14 53
rect 7 46 9 48
rect 11 46 14 48
rect 7 44 14 46
rect 16 60 24 62
rect 16 58 19 60
rect 21 58 24 60
rect 16 51 24 58
rect 26 62 34 64
rect 26 60 29 62
rect 31 60 34 62
rect 26 55 34 60
rect 26 53 29 55
rect 31 53 34 55
rect 26 51 34 53
rect 36 62 43 64
rect 36 60 39 62
rect 41 60 43 62
rect 62 62 69 64
rect 62 61 64 62
rect 36 51 43 60
rect 53 56 58 61
rect 51 54 58 56
rect 51 52 53 54
rect 55 52 58 54
rect 16 44 22 51
rect 51 47 58 52
rect 51 45 53 47
rect 55 45 58 47
rect 51 43 58 45
rect 60 60 64 61
rect 66 60 69 62
rect 60 43 69 60
rect -18 -50 -9 -33
rect -18 -52 -15 -50
rect -13 -51 -9 -50
rect -7 -35 0 -33
rect -7 -37 -4 -35
rect -2 -37 0 -35
rect -7 -42 0 -37
rect -7 -44 -4 -42
rect -2 -44 0 -42
rect -7 -46 0 -44
rect 7 -36 14 -34
rect 7 -38 9 -36
rect 11 -38 14 -36
rect 7 -43 14 -38
rect 7 -45 9 -43
rect 11 -45 14 -43
rect -7 -51 -2 -46
rect 7 -47 14 -45
rect -13 -52 -11 -51
rect -18 -54 -11 -52
rect 9 -52 14 -47
rect 16 -41 22 -34
rect 51 -35 58 -33
rect 51 -37 53 -35
rect 55 -37 58 -35
rect 16 -48 24 -41
rect 16 -50 19 -48
rect 21 -50 24 -48
rect 16 -52 24 -50
rect 18 -54 24 -52
rect 26 -43 34 -41
rect 26 -45 29 -43
rect 31 -45 34 -43
rect 26 -50 34 -45
rect 26 -52 29 -50
rect 31 -52 34 -50
rect 26 -54 34 -52
rect 36 -50 43 -41
rect 51 -42 58 -37
rect 51 -44 53 -42
rect 55 -44 58 -42
rect 51 -46 58 -44
rect 36 -52 39 -50
rect 41 -52 43 -50
rect 53 -51 58 -46
rect 60 -50 69 -33
rect 60 -51 64 -50
rect 36 -54 43 -52
rect 62 -52 64 -51
rect 66 -52 69 -50
rect 62 -54 69 -52
<< alu1 >>
rect -41 76 75 77
rect -41 74 -40 76
rect -38 74 75 76
rect -41 72 75 74
rect -41 70 -34 72
rect -32 70 10 72
rect 12 70 54 72
rect 56 70 66 72
rect 68 70 75 72
rect -41 69 75 70
rect -37 63 -33 64
rect -37 59 -24 63
rect -37 57 -35 59
rect -37 52 -33 57
rect -37 50 -35 52
rect -37 35 -33 50
rect 7 56 12 57
rect -5 55 12 56
rect -5 53 9 55
rect 11 53 12 55
rect -5 52 12 53
rect -37 33 -36 35
rect -34 33 -33 35
rect -37 31 -33 33
rect -5 47 -1 52
rect -22 45 -1 47
rect -22 43 -8 45
rect -6 43 -1 45
rect 7 48 12 52
rect 7 46 9 48
rect 11 46 12 48
rect 7 44 12 46
rect 39 52 43 56
rect 51 54 63 56
rect 51 52 53 54
rect 55 52 63 54
rect 39 50 63 52
rect -37 29 -32 31
rect -37 27 -35 29
rect -33 27 -32 29
rect -37 25 -32 27
rect -22 38 0 39
rect -22 36 -18 38
rect -16 36 -3 38
rect -1 36 0 38
rect -22 35 0 36
rect -5 26 0 35
rect 7 24 11 44
rect 39 48 55 50
rect 39 47 43 48
rect 30 46 43 47
rect 30 44 36 46
rect 38 44 43 46
rect 30 43 43 44
rect 51 47 55 48
rect 51 45 53 47
rect 22 38 36 39
rect 22 36 26 38
rect 28 36 36 38
rect 22 35 36 36
rect 31 33 47 35
rect 31 31 43 33
rect 46 31 47 33
rect 7 22 9 24
rect 11 22 19 24
rect 7 18 19 22
rect 31 30 47 31
rect 31 26 36 30
rect 51 29 55 45
rect 59 38 71 40
rect 59 36 60 38
rect 62 37 71 38
rect 62 36 68 37
rect 59 35 68 36
rect 70 35 71 37
rect 59 34 71 35
rect 51 27 53 29
rect 51 18 55 27
rect 59 26 63 34
rect -41 12 75 13
rect -41 10 -34 12
rect -32 10 10 12
rect 12 10 20 12
rect 22 10 54 12
rect 56 10 66 12
rect 68 10 75 12
rect -41 5 75 10
rect -24 0 75 5
rect -24 -2 -17 0
rect -15 -2 -5 0
rect -3 -2 10 0
rect 12 -2 20 0
rect 22 -2 54 0
rect 56 -2 66 0
rect 68 -2 75 0
rect -24 -3 75 -2
rect -12 -17 -8 -16
rect -12 -19 -11 -17
rect -9 -19 -8 -17
rect -12 -24 -8 -19
rect -4 -17 0 -8
rect -2 -19 0 -17
rect -20 -26 -8 -24
rect -20 -28 -11 -26
rect -9 -28 -8 -26
rect -20 -30 -8 -28
rect -4 -35 0 -19
rect -2 -37 0 -35
rect -4 -40 0 -37
rect -12 -42 0 -40
rect -12 -44 -4 -42
rect -2 -44 0 -42
rect -12 -46 0 -44
rect 7 -9 19 -8
rect 7 -11 8 -9
rect 10 -11 19 -9
rect 7 -12 19 -11
rect 7 -14 9 -12
rect 11 -14 19 -12
rect 7 -34 11 -14
rect 31 -23 36 -16
rect 51 -17 55 -8
rect 59 -12 63 -11
rect 59 -14 60 -12
rect 62 -14 63 -12
rect 51 -19 53 -17
rect 51 -23 55 -19
rect 31 -25 55 -23
rect 7 -36 12 -34
rect 7 -38 9 -36
rect 11 -38 12 -36
rect 7 -43 12 -38
rect 7 -45 9 -43
rect 11 -45 12 -43
rect 22 -26 55 -25
rect 22 -28 26 -26
rect 28 -28 55 -26
rect 22 -29 55 -28
rect 30 -34 43 -33
rect 30 -36 36 -34
rect 38 -35 43 -34
rect 38 -36 40 -35
rect 30 -37 40 -36
rect 42 -37 43 -35
rect 7 -47 12 -45
rect 39 -46 43 -37
rect 51 -35 55 -29
rect 59 -24 63 -14
rect 59 -26 71 -24
rect 59 -28 60 -26
rect 62 -28 71 -26
rect 59 -30 71 -28
rect 51 -37 53 -35
rect 51 -40 55 -37
rect 51 -42 63 -40
rect 51 -44 53 -42
rect 55 -44 63 -42
rect 51 -46 63 -44
rect -24 -60 75 -59
rect -24 -62 -17 -60
rect -15 -62 -5 -60
rect -3 -62 10 -60
rect 12 -62 54 -60
rect 56 -62 66 -60
rect 68 -62 75 -60
rect -24 -64 -23 -62
rect -21 -64 75 -62
rect -24 -67 75 -64
<< alu2 >>
rect -48 76 -36 77
rect -48 74 -40 76
rect -38 74 -36 76
rect -48 72 -36 74
rect -48 -61 -44 72
rect -4 38 4 39
rect -4 36 -3 38
rect -1 36 4 38
rect -37 35 -33 36
rect -4 35 4 36
rect -37 33 -36 35
rect -34 33 -33 35
rect -37 -16 -33 33
rect 0 -8 4 35
rect 67 37 73 38
rect 67 35 68 37
rect 70 35 73 37
rect 42 33 47 34
rect 42 31 43 33
rect 46 31 47 33
rect 42 30 47 31
rect 42 26 48 30
rect 44 -4 48 26
rect 44 -8 63 -4
rect 0 -9 11 -8
rect 0 -11 8 -9
rect 10 -11 11 -9
rect 0 -16 11 -11
rect 59 -12 63 -8
rect 59 -14 60 -12
rect 62 -14 63 -12
rect 59 -15 63 -14
rect -37 -17 -8 -16
rect -37 -19 -11 -17
rect -9 -19 -8 -17
rect -37 -20 -8 -19
rect 67 -34 73 35
rect 39 -35 73 -34
rect 39 -37 40 -35
rect 42 -37 73 -35
rect 39 -40 73 -37
rect -48 -62 -20 -61
rect -48 -64 -23 -62
rect -21 -64 -20 -62
rect -48 -66 -20 -64
<< ptie >>
rect -36 12 -30 14
rect 8 12 14 14
rect -36 10 -34 12
rect -32 10 -30 12
rect -36 8 -30 10
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect 52 12 70 14
rect 52 10 54 12
rect 56 10 66 12
rect 68 10 70 12
rect 52 8 70 10
rect -19 0 -1 2
rect -19 -2 -17 0
rect -15 -2 -5 0
rect -3 -2 -1 0
rect -19 -4 -1 -2
rect 8 0 14 2
rect 8 -2 10 0
rect 12 -2 14 0
rect 8 -4 14 -2
rect 52 0 70 2
rect 52 -2 54 0
rect 56 -2 66 0
rect 68 -2 70 0
rect 52 -4 70 -2
<< ntie >>
rect -36 72 -30 74
rect -36 70 -34 72
rect -32 70 -30 72
rect 8 72 14 74
rect -36 68 -30 70
rect 8 70 10 72
rect 12 70 14 72
rect 8 68 14 70
rect 52 72 70 74
rect 52 70 54 72
rect 56 70 66 72
rect 68 70 70 72
rect 52 68 70 70
rect -19 -60 -1 -58
rect -19 -62 -17 -60
rect -15 -62 -5 -60
rect -3 -62 -1 -60
rect -19 -64 -1 -62
rect 8 -60 14 -58
rect 8 -62 10 -60
rect 12 -62 14 -60
rect 8 -64 14 -62
rect 52 -60 70 -58
rect 52 -62 54 -60
rect 56 -62 66 -60
rect 68 -62 70 -60
rect 52 -64 70 -62
<< nmos >>
rect -30 22 -28 31
rect -20 25 -18 31
rect -10 25 -8 31
rect 14 20 16 29
rect 27 18 29 29
rect 34 18 36 29
rect 58 22 60 31
rect -9 -21 -7 -12
rect 14 -19 16 -10
rect 27 -19 29 -8
rect 34 -19 36 -8
rect 58 -21 60 -12
<< pmos >>
rect -30 43 -28 61
rect -17 50 -15 71
rect -10 50 -8 71
rect 14 44 16 62
rect 24 51 26 64
rect 34 51 36 64
rect 58 43 60 61
rect -9 -51 -7 -33
rect 14 -52 16 -34
rect 24 -54 26 -41
rect 34 -54 36 -41
rect 58 -51 60 -33
<< polyct0 >>
rect -28 36 -26 38
rect 16 36 18 38
rect 16 -28 18 -26
<< polyct1 >>
rect -8 43 -6 45
rect -18 36 -16 38
rect 36 44 38 46
rect 26 36 28 38
rect 60 36 62 38
rect -11 -28 -9 -26
rect 26 -28 28 -26
rect 60 -28 62 -26
rect 36 -36 38 -34
<< ndifct0 >>
rect -15 27 -13 29
rect -24 14 -22 16
rect 67 24 69 26
rect 39 20 41 22
rect -5 14 -3 16
rect -18 -16 -16 -14
rect 39 -12 41 -10
rect 67 -16 69 -14
<< ndifct1 >>
rect -35 27 -33 29
rect 9 22 11 24
rect 53 27 55 29
rect 20 10 22 12
rect 20 -2 22 0
rect 9 -14 11 -12
rect -4 -19 -2 -17
rect 53 -19 55 -17
<< ntiect1 >>
rect -34 70 -32 72
rect 10 70 12 72
rect 54 70 56 72
rect 66 70 68 72
rect -17 -62 -15 -60
rect -5 -62 -3 -60
rect 10 -62 12 -60
rect 54 -62 56 -60
rect 66 -62 68 -60
<< ptiect1 >>
rect -34 10 -32 12
rect 10 10 12 12
rect 54 10 56 12
rect 66 10 68 12
rect -17 -2 -15 0
rect -5 -2 -3 0
rect 10 -2 12 0
rect 54 -2 56 0
rect 66 -2 68 0
<< pdifct0 >>
rect -24 67 -22 69
rect -5 60 -3 62
rect 19 58 21 60
rect 29 60 31 62
rect 29 53 31 55
rect 39 60 41 62
rect 64 60 66 62
rect -15 -52 -13 -50
rect 19 -50 21 -48
rect 29 -45 31 -43
rect 29 -52 31 -50
rect 39 -52 41 -50
rect 64 -52 66 -50
<< pdifct1 >>
rect -35 57 -33 59
rect -35 50 -33 52
rect 9 53 11 55
rect 9 46 11 48
rect 53 52 55 54
rect 53 45 55 47
rect -4 -37 -2 -35
rect -4 -44 -2 -42
rect 9 -38 11 -36
rect 9 -45 11 -43
rect 53 -37 55 -35
rect 53 -44 55 -42
<< alu0 >>
rect -26 67 -24 69
rect -22 67 -20 69
rect -26 66 -20 67
rect -18 62 -1 63
rect -18 60 -5 62
rect -3 60 -1 62
rect -18 59 -1 60
rect 17 60 23 69
rect -33 48 -32 59
rect -18 55 -14 59
rect 17 58 19 60
rect 21 58 23 60
rect 17 57 23 58
rect 28 62 32 64
rect 28 60 29 62
rect 31 60 32 62
rect -29 51 -14 55
rect 28 55 32 60
rect 37 62 43 69
rect 37 60 39 62
rect 41 60 43 62
rect 37 59 43 60
rect 62 62 68 69
rect 62 60 64 62
rect 66 60 68 62
rect 62 59 68 60
rect 28 54 29 55
rect -29 38 -25 51
rect 15 53 29 54
rect 31 53 32 55
rect 15 50 32 53
rect -10 42 -4 43
rect -29 36 -28 38
rect -26 36 -25 38
rect -29 30 -25 36
rect -29 29 -11 30
rect -29 27 -15 29
rect -13 27 -11 29
rect -29 26 -11 27
rect 15 38 19 50
rect 15 36 16 38
rect 18 36 19 38
rect 15 31 19 36
rect 15 27 27 31
rect 11 24 12 26
rect 23 23 27 27
rect 55 43 56 50
rect 23 22 43 23
rect 23 20 39 22
rect 41 20 43 22
rect 23 19 43 20
rect 55 25 56 31
rect 66 26 70 28
rect 66 24 67 26
rect 69 24 70 26
rect -26 16 -20 17
rect -26 14 -24 16
rect -22 14 -20 16
rect -26 13 -20 14
rect -7 16 -1 17
rect -7 14 -5 16
rect -3 14 -1 16
rect -7 13 -1 14
rect 66 13 70 24
rect -19 -14 -15 -3
rect -19 -16 -18 -14
rect -16 -16 -15 -14
rect -19 -18 -15 -16
rect -5 -21 -4 -15
rect -5 -40 -4 -33
rect 23 -10 43 -9
rect 23 -12 39 -10
rect 41 -12 43 -10
rect 23 -13 43 -12
rect 11 -16 12 -14
rect 23 -17 27 -13
rect 15 -21 27 -17
rect 15 -26 19 -21
rect 55 -21 56 -15
rect 15 -28 16 -26
rect 18 -28 19 -26
rect 15 -40 19 -28
rect 15 -43 32 -40
rect 15 -44 29 -43
rect 28 -45 29 -44
rect 31 -45 32 -43
rect 17 -48 23 -47
rect -17 -50 -11 -49
rect -17 -52 -15 -50
rect -13 -52 -11 -50
rect -17 -59 -11 -52
rect 17 -50 19 -48
rect 21 -50 23 -48
rect 17 -59 23 -50
rect 28 -50 32 -45
rect 66 -14 70 -3
rect 66 -16 67 -14
rect 69 -16 70 -14
rect 66 -18 70 -16
rect 55 -40 56 -33
rect 28 -52 29 -50
rect 31 -52 32 -50
rect 28 -54 32 -52
rect 37 -50 43 -49
rect 37 -52 39 -50
rect 41 -52 43 -50
rect 37 -59 43 -52
rect 62 -50 68 -49
rect 62 -52 64 -50
rect 66 -52 68 -50
rect 62 -59 68 -52
<< via1 >>
rect -40 74 -38 76
rect -36 33 -34 35
rect -3 36 -1 38
rect 43 31 46 33
rect 68 35 70 37
rect -11 -19 -9 -17
rect 8 -11 10 -9
rect 60 -14 62 -12
rect 40 -37 42 -35
rect -23 -64 -21 -62
<< labels >>
rlabel alu1 25 9 25 9 6 vss
rlabel alu1 25 37 25 37 6 a
rlabel alu1 33 33 33 33 6 a
rlabel alu1 25 73 25 73 6 vdd
rlabel alu1 41 53 41 53 1 binv
rlabel alu1 33 45 33 45 1 binv
rlabel alu0 17 40 17 40 1 tempand1
rlabel alu1 9 37 9 37 1 outand1
rlabel alu0 33 21 33 21 1 tempand1
rlabel alu1 17 21 17 21 1 outand1
rlabel alu0 30 57 30 57 1 tempand1
rlabel alu1 17 -11 17 -11 8 z
rlabel alu1 25 1 25 1 8 vss
rlabel alu1 33 -35 33 -35 8 b
rlabel alu1 25 -63 25 -63 8 vdd
rlabel alu1 41 -43 41 -43 8 b
rlabel alu0 33 -11 33 -11 1 tempand2
rlabel alu0 17 -30 17 -30 1 tempand2
rlabel alu0 30 -47 30 -47 1 tempand2
rlabel alu1 9 -27 9 -27 1 outand2
rlabel alu1 33 -23 33 -23 1 ainv
rlabel alu1 25 -27 25 -27 1 ainv
rlabel alu1 61 9 61 9 6 vss
rlabel alu1 61 73 61 73 6 vdd
rlabel alu1 61 1 61 1 8 vss
rlabel alu1 61 -23 61 -23 8 a
rlabel alu1 61 -63 61 -63 8 vdd
rlabel alu1 69 -27 69 -27 8 a
rlabel alu1 69 37 69 37 1 b
rlabel alu1 61 33 61 33 1 b
rlabel alu1 61 53 61 53 1 binv
rlabel alu1 53 37 53 37 1 binv
rlabel alu1 61 -43 61 -43 1 ainv
rlabel alu1 53 -27 53 -27 1 ainv
rlabel alu1 -19 9 -19 9 6 vss
rlabel alu1 -19 73 -19 73 6 vdd
rlabel alu1 -3 53 -3 53 1 outand1
rlabel alu1 -11 45 -11 45 1 outand1
rlabel alu1 -19 45 -19 45 1 outand1
rlabel alu0 -10 61 -10 61 1 tempor
rlabel alu0 -27 40 -27 40 1 tempor
rlabel alu0 -20 28 -20 28 1 tempor
rlabel alu1 -27 61 -27 61 1 outor
rlabel alu1 -35 45 -35 45 1 outor
rlabel alu1 -19 37 -19 37 1 outand2
rlabel alu1 -11 37 -11 37 1 outand2
rlabel alu1 -3 29 -3 29 1 outand2
rlabel alu1 -10 1 -10 1 2 vss
rlabel alu1 -10 -63 -10 -63 2 vdd
rlabel alu1 -18 -27 -18 -27 1 outor
rlabel alu1 -10 -23 -10 -23 1 outor
rlabel alu1 -10 -43 -10 -43 1 out
rlabel alu1 -2 -27 -2 -27 1 out
<< end >>
