magic
tech scmos
timestamp 1199202487
<< ab >>
rect 0 0 224 72
<< nwell >>
rect -5 32 229 77
<< pwell >>
rect -5 -5 229 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 59 67 81 69
rect 59 61 61 67
rect 69 64 71 67
rect 79 64 81 67
rect 139 68 205 70
rect 139 65 141 68
rect 49 59 61 61
rect 49 56 51 59
rect 59 56 61 59
rect 89 60 91 65
rect 99 63 141 65
rect 99 60 101 63
rect 109 60 111 63
rect 119 60 121 63
rect 129 60 131 63
rect 139 60 141 63
rect 149 60 151 64
rect 163 60 165 64
rect 173 60 175 64
rect 183 60 185 64
rect 193 60 195 64
rect 203 60 205 68
rect 213 54 215 59
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 33 41 35
rect 49 34 51 38
rect 59 34 61 38
rect 69 34 71 38
rect 79 35 81 38
rect 89 35 91 38
rect 9 31 11 33
rect 13 31 19 33
rect 21 31 41 33
rect 9 29 41 31
rect 79 33 91 35
rect 99 34 101 38
rect 109 34 111 38
rect 119 35 121 38
rect 79 31 85 33
rect 87 31 91 33
rect 19 26 21 29
rect 29 26 31 29
rect 39 26 41 29
rect 49 26 51 30
rect 59 26 61 30
rect 69 26 71 30
rect 79 29 91 31
rect 119 33 125 35
rect 129 33 131 38
rect 139 33 141 38
rect 149 35 151 38
rect 163 35 165 38
rect 173 35 175 38
rect 183 35 185 38
rect 193 35 195 38
rect 149 33 195 35
rect 203 35 205 38
rect 213 35 215 38
rect 119 31 121 33
rect 123 31 125 33
rect 79 26 81 29
rect 89 26 91 29
rect 99 26 101 30
rect 109 26 111 30
rect 119 29 125 31
rect 149 31 151 33
rect 153 31 159 33
rect 161 31 181 33
rect 149 29 181 31
rect 79 9 81 13
rect 89 10 91 13
rect 99 10 101 13
rect 109 10 111 13
rect 89 8 111 10
rect 19 3 21 8
rect 29 3 31 8
rect 39 3 41 8
rect 49 4 51 8
rect 59 4 61 8
rect 69 4 71 8
rect 120 4 122 29
rect 149 26 151 29
rect 159 26 161 29
rect 169 26 171 29
rect 179 26 181 29
rect 203 29 215 35
rect 203 26 205 29
rect 213 26 215 29
rect 49 2 122 4
rect 149 7 151 12
rect 159 7 161 12
rect 169 7 171 12
rect 179 7 181 12
rect 203 10 205 15
rect 213 11 215 15
<< ndif >>
rect 11 20 19 26
rect 11 18 14 20
rect 16 18 19 20
rect 11 12 19 18
rect 11 10 14 12
rect 16 10 19 12
rect 11 8 19 10
rect 21 24 29 26
rect 21 22 24 24
rect 26 22 29 24
rect 21 17 29 22
rect 21 15 24 17
rect 26 15 29 17
rect 21 8 29 15
rect 31 12 39 26
rect 31 10 34 12
rect 36 10 39 12
rect 31 8 39 10
rect 41 24 49 26
rect 41 22 44 24
rect 46 22 49 24
rect 41 17 49 22
rect 41 15 44 17
rect 46 15 49 17
rect 41 8 49 15
rect 51 24 59 26
rect 51 22 54 24
rect 56 22 59 24
rect 51 8 59 22
rect 61 16 69 26
rect 61 14 64 16
rect 66 14 69 16
rect 61 8 69 14
rect 71 24 79 26
rect 71 22 74 24
rect 76 22 79 24
rect 71 17 79 22
rect 71 15 74 17
rect 76 15 79 17
rect 71 13 79 15
rect 81 17 89 26
rect 81 15 84 17
rect 86 15 89 17
rect 81 13 89 15
rect 91 24 99 26
rect 91 22 94 24
rect 96 22 99 24
rect 91 13 99 22
rect 101 17 109 26
rect 101 15 104 17
rect 106 15 109 17
rect 101 13 109 15
rect 111 24 118 26
rect 111 22 114 24
rect 116 22 118 24
rect 111 20 118 22
rect 111 13 116 20
rect 71 8 76 13
rect 141 12 149 26
rect 151 24 159 26
rect 151 22 154 24
rect 156 22 159 24
rect 151 17 159 22
rect 151 15 154 17
rect 156 15 159 17
rect 151 12 159 15
rect 161 16 169 26
rect 161 14 164 16
rect 166 14 169 16
rect 161 12 169 14
rect 171 24 179 26
rect 171 22 174 24
rect 176 22 179 24
rect 171 17 179 22
rect 171 15 174 17
rect 176 15 179 17
rect 171 12 179 15
rect 181 24 189 26
rect 181 22 184 24
rect 186 22 189 24
rect 181 16 189 22
rect 181 14 184 16
rect 186 14 189 16
rect 195 19 203 26
rect 195 17 198 19
rect 200 17 203 19
rect 195 15 203 17
rect 205 24 213 26
rect 205 22 208 24
rect 210 22 213 24
rect 205 15 213 22
rect 215 19 222 26
rect 215 17 218 19
rect 220 17 222 19
rect 215 15 222 17
rect 181 12 189 14
rect 141 7 147 12
rect 141 5 143 7
rect 145 5 147 7
rect 141 3 147 5
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 19 66
rect 11 62 14 64
rect 16 62 19 64
rect 11 57 19 62
rect 11 55 14 57
rect 16 55 19 57
rect 11 38 19 55
rect 21 49 29 66
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 64 39 66
rect 31 62 34 64
rect 36 62 39 64
rect 31 57 39 62
rect 31 55 34 57
rect 36 55 39 57
rect 31 38 39 55
rect 41 56 46 66
rect 64 56 69 64
rect 41 49 49 56
rect 41 47 44 49
rect 46 47 49 49
rect 41 42 49 47
rect 41 40 44 42
rect 46 40 49 42
rect 41 38 49 40
rect 51 49 59 56
rect 51 47 54 49
rect 56 47 59 49
rect 51 42 59 47
rect 51 40 54 42
rect 56 40 59 42
rect 51 38 59 40
rect 61 54 69 56
rect 61 52 64 54
rect 66 52 69 54
rect 61 47 69 52
rect 61 45 64 47
rect 66 45 69 47
rect 61 38 69 45
rect 71 49 79 64
rect 71 47 74 49
rect 76 47 79 49
rect 71 42 79 47
rect 71 40 74 42
rect 76 40 79 42
rect 71 38 79 40
rect 81 60 86 64
rect 81 58 89 60
rect 81 56 84 58
rect 86 56 89 58
rect 81 38 89 56
rect 91 42 99 60
rect 91 40 94 42
rect 96 40 99 42
rect 91 38 99 40
rect 101 50 109 60
rect 101 48 104 50
rect 106 48 109 50
rect 101 38 109 48
rect 111 42 119 60
rect 111 40 114 42
rect 116 40 119 42
rect 111 38 119 40
rect 121 50 129 60
rect 121 48 124 50
rect 126 48 129 50
rect 121 38 129 48
rect 131 42 139 60
rect 131 40 134 42
rect 136 40 139 42
rect 131 38 139 40
rect 141 49 149 60
rect 141 47 144 49
rect 146 47 149 49
rect 141 42 149 47
rect 141 40 144 42
rect 146 40 149 42
rect 141 38 149 40
rect 151 58 163 60
rect 151 56 158 58
rect 160 56 163 58
rect 151 38 163 56
rect 165 42 173 60
rect 165 40 168 42
rect 170 40 173 42
rect 165 38 173 40
rect 175 58 183 60
rect 175 56 178 58
rect 180 56 183 58
rect 175 38 183 56
rect 185 42 193 60
rect 185 40 188 42
rect 190 40 193 42
rect 185 38 193 40
rect 195 58 203 60
rect 195 56 198 58
rect 200 56 203 58
rect 195 38 203 56
rect 205 54 210 60
rect 205 49 213 54
rect 205 47 208 49
rect 210 47 213 49
rect 205 42 213 47
rect 205 40 208 42
rect 210 40 213 42
rect 205 38 213 40
rect 215 52 222 54
rect 215 50 218 52
rect 220 50 222 52
rect 215 44 222 50
rect 215 42 218 44
rect 220 42 222 44
rect 215 38 222 42
<< alu1 >>
rect -2 67 226 72
rect -2 65 52 67
rect 54 65 217 67
rect 219 65 226 67
rect -2 64 226 65
rect 2 33 22 35
rect 2 31 11 33
rect 13 31 19 33
rect 21 31 22 33
rect 2 29 22 31
rect 2 13 6 29
rect 53 49 57 51
rect 53 47 54 49
rect 56 47 57 49
rect 53 42 57 47
rect 73 49 78 52
rect 73 47 74 49
rect 76 47 78 49
rect 53 40 54 42
rect 56 40 57 42
rect 53 26 57 40
rect 73 42 78 47
rect 73 40 74 42
rect 76 40 78 42
rect 73 26 78 40
rect 92 42 98 43
rect 112 42 118 43
rect 132 42 138 43
rect 92 40 94 42
rect 96 40 114 42
rect 116 40 134 42
rect 136 40 138 42
rect 92 38 138 40
rect 98 26 102 38
rect 119 33 135 34
rect 119 31 121 33
rect 123 31 135 33
rect 119 30 135 31
rect 53 24 119 26
rect 53 22 54 24
rect 56 22 74 24
rect 76 22 94 24
rect 96 22 114 24
rect 116 22 119 24
rect 129 22 135 30
rect 146 33 166 35
rect 146 31 151 33
rect 153 31 159 33
rect 161 31 166 33
rect 146 29 166 31
rect 53 20 57 22
rect 73 17 78 22
rect 92 21 98 22
rect 112 21 119 22
rect 146 21 150 29
rect 73 15 74 17
rect 76 15 78 17
rect 73 13 78 15
rect -2 7 226 8
rect -2 5 126 7
rect 128 5 133 7
rect 135 5 143 7
rect 145 5 209 7
rect 211 5 217 7
rect 219 5 226 7
rect -2 0 226 5
<< ptie >>
rect 124 7 137 9
rect 124 5 126 7
rect 128 5 133 7
rect 135 5 137 7
rect 124 3 137 5
rect 207 7 221 9
rect 207 5 209 7
rect 211 5 217 7
rect 219 5 221 7
rect 207 3 221 5
<< ntie >>
rect 50 67 56 69
rect 50 65 52 67
rect 54 65 56 67
rect 50 63 56 65
rect 215 67 221 69
rect 215 65 217 67
rect 219 65 221 67
rect 215 63 221 65
<< nmos >>
rect 19 8 21 26
rect 29 8 31 26
rect 39 8 41 26
rect 49 8 51 26
rect 59 8 61 26
rect 69 8 71 26
rect 79 13 81 26
rect 89 13 91 26
rect 99 13 101 26
rect 109 13 111 26
rect 149 12 151 26
rect 159 12 161 26
rect 169 12 171 26
rect 179 12 181 26
rect 203 15 205 26
rect 213 15 215 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 56
rect 59 38 61 56
rect 69 38 71 64
rect 79 38 81 64
rect 89 38 91 60
rect 99 38 101 60
rect 109 38 111 60
rect 119 38 121 60
rect 129 38 131 60
rect 139 38 141 60
rect 149 38 151 60
rect 163 38 165 60
rect 173 38 175 60
rect 183 38 185 60
rect 193 38 195 60
rect 203 38 205 60
rect 213 38 215 54
<< polyct0 >>
rect 85 31 87 33
<< polyct1 >>
rect 11 31 13 33
rect 19 31 21 33
rect 121 31 123 33
rect 151 31 153 33
rect 159 31 161 33
<< ndifct0 >>
rect 14 18 16 20
rect 14 10 16 12
rect 24 22 26 24
rect 24 15 26 17
rect 34 10 36 12
rect 44 22 46 24
rect 44 15 46 17
rect 64 14 66 16
rect 84 15 86 17
rect 104 15 106 17
rect 154 22 156 24
rect 154 15 156 17
rect 164 14 166 16
rect 174 22 176 24
rect 174 15 176 17
rect 184 22 186 24
rect 184 14 186 16
rect 198 17 200 19
rect 208 22 210 24
rect 218 17 220 19
<< ndifct1 >>
rect 54 22 56 24
rect 74 22 76 24
rect 74 15 76 17
rect 94 22 96 24
rect 114 22 116 24
rect 143 5 145 7
<< ntiect1 >>
rect 52 65 54 67
rect 217 65 219 67
<< ptiect1 >>
rect 126 5 128 7
rect 133 5 135 7
rect 209 5 211 7
rect 217 5 219 7
<< pdifct0 >>
rect 4 47 6 49
rect 4 40 6 42
rect 14 62 16 64
rect 14 55 16 57
rect 24 47 26 49
rect 24 40 26 42
rect 34 62 36 64
rect 34 55 36 57
rect 44 47 46 49
rect 44 40 46 42
rect 64 52 66 54
rect 64 45 66 47
rect 84 56 86 58
rect 104 48 106 50
rect 124 48 126 50
rect 144 47 146 49
rect 144 40 146 42
rect 158 56 160 58
rect 168 40 170 42
rect 178 56 180 58
rect 188 40 190 42
rect 198 56 200 58
rect 208 47 210 49
rect 208 40 210 42
rect 218 50 220 52
rect 218 42 220 44
<< pdifct1 >>
rect 54 47 56 49
rect 54 40 56 42
rect 74 47 76 49
rect 74 40 76 42
rect 94 40 96 42
rect 114 40 116 42
rect 134 40 136 42
<< alu0 >>
rect 13 62 14 64
rect 16 62 17 64
rect 13 57 17 62
rect 13 55 14 57
rect 16 55 17 57
rect 13 53 17 55
rect 33 62 34 64
rect 36 62 37 64
rect 33 57 37 62
rect 33 55 34 57
rect 36 55 37 57
rect 33 53 37 55
rect 43 58 88 59
rect 43 56 84 58
rect 86 56 88 58
rect 43 55 88 56
rect 93 55 154 59
rect 3 49 7 51
rect 3 47 4 49
rect 6 47 7 49
rect 3 42 7 47
rect 23 49 27 51
rect 23 47 24 49
rect 26 47 27 49
rect 23 42 27 47
rect 43 49 47 55
rect 63 54 67 55
rect 63 52 64 54
rect 66 52 67 54
rect 43 47 44 49
rect 46 47 47 49
rect 43 42 47 47
rect 3 40 4 42
rect 6 40 24 42
rect 26 40 44 42
rect 46 40 47 42
rect 3 38 47 40
rect 43 26 47 38
rect 23 24 47 26
rect 23 22 24 24
rect 26 22 44 24
rect 46 22 47 24
rect 13 20 17 22
rect 13 18 14 20
rect 16 18 17 20
rect 13 12 17 18
rect 23 17 27 22
rect 23 15 24 17
rect 26 15 27 17
rect 23 13 27 15
rect 43 17 47 22
rect 63 47 67 52
rect 63 45 64 47
rect 66 45 67 47
rect 63 43 67 45
rect 93 51 97 55
rect 150 51 154 55
rect 157 58 161 64
rect 157 56 158 58
rect 160 56 161 58
rect 157 54 161 56
rect 177 58 181 64
rect 177 56 178 58
rect 180 56 181 58
rect 177 54 181 56
rect 196 58 202 64
rect 196 56 198 58
rect 200 56 202 58
rect 196 55 202 56
rect 217 52 221 64
rect 84 47 97 51
rect 102 50 147 51
rect 102 48 104 50
rect 106 48 124 50
rect 126 49 147 50
rect 126 48 144 49
rect 102 47 144 48
rect 146 47 147 49
rect 150 49 211 51
rect 150 47 208 49
rect 210 47 211 49
rect 84 33 88 47
rect 142 43 147 47
rect 142 42 192 43
rect 142 40 144 42
rect 146 40 168 42
rect 170 40 188 42
rect 190 40 192 42
rect 142 39 192 40
rect 207 42 211 47
rect 207 40 208 42
rect 210 40 211 42
rect 217 50 218 52
rect 220 50 221 52
rect 217 44 221 50
rect 217 42 218 44
rect 220 42 221 44
rect 217 40 221 42
rect 84 31 85 33
rect 87 31 88 33
rect 84 29 88 31
rect 173 26 177 39
rect 153 24 177 26
rect 153 22 154 24
rect 156 22 174 24
rect 176 22 177 24
rect 153 18 158 22
rect 43 15 44 17
rect 46 16 68 17
rect 46 15 64 16
rect 43 14 64 15
rect 66 14 68 16
rect 13 10 14 12
rect 16 10 17 12
rect 13 8 17 10
rect 33 12 37 14
rect 43 13 68 14
rect 82 17 158 18
rect 82 15 84 17
rect 86 15 104 17
rect 106 15 154 17
rect 156 15 158 17
rect 82 14 158 15
rect 163 16 167 18
rect 163 14 164 16
rect 166 14 167 16
rect 33 10 34 12
rect 36 10 37 12
rect 33 8 37 10
rect 163 8 167 14
rect 173 17 177 22
rect 173 15 174 17
rect 176 15 177 17
rect 173 13 177 15
rect 183 24 187 26
rect 183 22 184 24
rect 186 22 187 24
rect 183 16 187 22
rect 207 24 211 40
rect 207 22 208 24
rect 210 22 211 24
rect 183 14 184 16
rect 186 14 187 16
rect 183 8 187 14
rect 197 19 201 21
rect 207 20 211 22
rect 197 17 198 19
rect 200 17 201 19
rect 197 8 201 17
rect 217 19 221 21
rect 217 17 218 19
rect 220 17 221 19
rect 217 8 221 17
<< labels >>
rlabel alu0 25 19 25 19 6 a1n
rlabel alu0 5 44 5 44 6 a1n
rlabel alu0 25 44 25 44 6 a1n
rlabel alu0 45 36 45 36 6 a1n
rlabel alu0 55 15 55 15 6 a1n
rlabel alu0 86 40 86 40 6 sn
rlabel alu0 65 51 65 51 6 a1n
rlabel alu0 120 16 120 16 6 a0n
rlabel alu0 155 20 155 20 6 a0n
rlabel alu0 124 49 124 49 6 a0n
rlabel alu0 144 45 144 45 6 a0n
rlabel alu0 175 28 175 28 6 a0n
rlabel alu0 209 35 209 35 6 sn
rlabel alu0 167 41 167 41 6 a0n
rlabel alu1 4 24 4 24 6 a1
rlabel polyct1 20 32 20 32 6 a1
rlabel polyct1 12 32 12 32 6 a1
rlabel alu1 100 32 100 32 6 z
rlabel alu1 108 24 108 24 6 z
rlabel alu1 92 24 92 24 6 z
rlabel alu1 76 32 76 32 6 z
rlabel alu1 60 24 60 24 6 z
rlabel alu1 68 24 68 24 6 z
rlabel alu1 84 24 84 24 6 z
rlabel alu1 108 40 108 40 6 z
rlabel alu1 112 4 112 4 6 vss
rlabel alu1 116 24 116 24 6 z
rlabel alu1 148 28 148 28 6 a0
rlabel alu1 156 32 156 32 6 a0
rlabel alu1 164 32 164 32 6 a0
rlabel alu1 132 28 132 28 6 s
rlabel alu1 124 32 124 32 6 s
rlabel alu1 132 40 132 40 6 z
rlabel alu1 124 40 124 40 6 z
rlabel alu1 116 40 116 40 6 z
rlabel alu1 112 68 112 68 6 vdd
<< end >>
