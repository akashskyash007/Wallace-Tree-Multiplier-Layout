magic
tech scmos
timestamp 1199201813
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 9 60 11 65
rect 21 60 23 65
rect 61 62 63 67
rect 39 54 41 59
rect 49 54 51 59
rect 9 45 11 48
rect 9 43 15 45
rect 9 41 11 43
rect 13 41 15 43
rect 9 39 15 41
rect 9 18 11 39
rect 21 35 23 48
rect 61 43 63 46
rect 60 41 66 43
rect 60 39 62 41
rect 64 39 66 41
rect 39 35 41 38
rect 17 33 23 35
rect 17 31 19 33
rect 21 31 23 33
rect 17 29 23 31
rect 33 33 41 35
rect 33 31 35 33
rect 37 31 41 33
rect 49 35 51 38
rect 60 37 66 39
rect 49 33 55 35
rect 49 31 51 33
rect 53 31 55 33
rect 33 29 45 31
rect 49 29 55 31
rect 21 26 23 29
rect 43 26 45 29
rect 53 26 55 29
rect 60 26 62 37
rect 21 15 23 20
rect 9 7 11 12
rect 43 15 45 20
rect 53 14 55 19
rect 60 14 62 19
<< ndif >>
rect 13 20 21 26
rect 23 24 30 26
rect 23 22 26 24
rect 28 22 30 24
rect 23 20 30 22
rect 34 20 43 26
rect 45 24 53 26
rect 45 22 48 24
rect 50 22 53 24
rect 45 20 53 22
rect 13 18 19 20
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 12 19 18
rect 13 7 19 12
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
rect 34 7 41 20
rect 48 19 53 20
rect 55 19 60 26
rect 62 23 69 26
rect 62 21 65 23
rect 67 21 69 23
rect 62 19 69 21
rect 34 5 37 7
rect 39 5 41 7
rect 34 3 41 5
<< pdif >>
rect 13 67 19 69
rect 13 65 15 67
rect 17 65 19 67
rect 13 60 19 65
rect 53 60 61 62
rect 4 54 9 60
rect 2 52 9 54
rect 2 50 4 52
rect 6 50 9 52
rect 2 48 9 50
rect 11 48 21 60
rect 23 54 28 60
rect 53 58 55 60
rect 57 58 61 60
rect 53 54 61 58
rect 23 52 30 54
rect 23 50 26 52
rect 28 50 30 52
rect 23 48 30 50
rect 34 44 39 54
rect 32 42 39 44
rect 32 40 34 42
rect 36 40 39 42
rect 32 38 39 40
rect 41 50 49 54
rect 41 48 44 50
rect 46 48 49 50
rect 41 38 49 48
rect 51 46 61 54
rect 63 59 68 62
rect 63 57 70 59
rect 63 55 66 57
rect 68 55 70 57
rect 63 50 70 55
rect 63 48 66 50
rect 68 48 70 50
rect 63 46 70 48
rect 51 38 58 46
<< alu1 >>
rect -2 67 74 72
rect -2 65 15 67
rect 17 65 37 67
rect 39 65 45 67
rect 47 65 74 67
rect -2 64 74 65
rect 10 53 22 59
rect 10 43 14 53
rect 10 41 11 43
rect 13 41 14 43
rect 10 39 14 41
rect 18 35 22 43
rect 10 33 22 35
rect 10 31 19 33
rect 21 31 22 33
rect 10 29 22 31
rect 33 43 38 51
rect 33 42 46 43
rect 33 40 34 42
rect 36 40 46 42
rect 33 37 46 40
rect 57 41 70 43
rect 57 39 62 41
rect 64 39 70 41
rect 57 38 70 39
rect 10 21 14 29
rect 42 25 46 37
rect 42 24 52 25
rect 42 22 48 24
rect 50 22 52 24
rect 42 21 52 22
rect 66 29 70 38
rect -2 7 74 8
rect -2 5 15 7
rect 17 5 26 7
rect 28 5 37 7
rect 39 5 57 7
rect 59 5 65 7
rect 67 5 74 7
rect -2 0 74 5
<< ptie >>
rect 24 7 30 9
rect 24 5 26 7
rect 28 5 30 7
rect 24 3 30 5
rect 55 7 69 9
rect 55 5 57 7
rect 59 5 65 7
rect 67 5 69 7
rect 55 3 69 5
<< ntie >>
rect 35 67 49 69
rect 35 65 37 67
rect 39 65 45 67
rect 47 65 49 67
rect 35 63 49 65
<< nmos >>
rect 21 20 23 26
rect 43 20 45 26
rect 9 12 11 18
rect 53 19 55 26
rect 60 19 62 26
<< pmos >>
rect 9 48 11 60
rect 21 48 23 60
rect 39 38 41 54
rect 49 38 51 54
rect 61 46 63 62
<< polyct0 >>
rect 35 31 37 33
rect 51 31 53 33
<< polyct1 >>
rect 11 41 13 43
rect 62 39 64 41
rect 19 31 21 33
<< ndifct0 >>
rect 26 22 28 24
rect 4 14 6 16
rect 65 21 67 23
<< ndifct1 >>
rect 48 22 50 24
rect 15 5 17 7
rect 37 5 39 7
<< ntiect1 >>
rect 37 65 39 67
rect 45 65 47 67
<< ptiect1 >>
rect 26 5 28 7
rect 57 5 59 7
rect 65 5 67 7
<< pdifct0 >>
rect 4 50 6 52
rect 55 58 57 60
rect 26 50 28 52
rect 44 48 46 50
rect 66 55 68 57
rect 66 48 68 50
<< pdifct1 >>
rect 15 65 17 67
rect 34 40 36 42
<< alu0 >>
rect 54 60 58 64
rect 2 52 7 54
rect 2 50 4 52
rect 6 50 7 52
rect 2 48 7 50
rect 54 58 55 60
rect 57 58 58 60
rect 54 56 58 58
rect 64 57 70 58
rect 64 55 66 57
rect 68 55 70 57
rect 2 17 6 48
rect 25 52 29 54
rect 25 50 26 52
rect 28 50 29 52
rect 64 51 70 55
rect 25 34 29 50
rect 42 50 70 51
rect 42 48 44 50
rect 46 48 66 50
rect 68 48 70 50
rect 42 47 70 48
rect 25 33 39 34
rect 25 31 35 33
rect 37 31 39 33
rect 25 30 39 31
rect 25 24 29 30
rect 25 22 26 24
rect 28 22 29 24
rect 25 20 29 22
rect 49 33 60 34
rect 49 31 51 33
rect 53 31 60 33
rect 49 30 60 31
rect 56 17 60 30
rect 2 16 60 17
rect 2 14 4 16
rect 6 14 60 16
rect 2 13 60 14
rect 64 23 68 25
rect 64 21 65 23
rect 67 21 68 23
rect 64 8 68 21
<< labels >>
rlabel alu0 4 33 4 33 6 a2n
rlabel alu0 27 37 27 37 6 bn
rlabel alu0 32 32 32 32 6 bn
rlabel alu0 31 15 31 15 6 a2n
rlabel alu0 54 32 54 32 6 a2n
rlabel alu0 56 49 56 49 6 n1
rlabel alu0 67 52 67 52 6 n1
rlabel alu1 12 28 12 28 6 b
rlabel alu1 12 52 12 52 6 a2
rlabel alu1 20 36 20 36 6 b
rlabel alu1 20 56 20 56 6 a2
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 44 32 44 32 6 z
rlabel alu1 36 40 36 40 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 40 60 40 6 a1
rlabel alu1 68 36 68 36 6 a1
<< end >>
