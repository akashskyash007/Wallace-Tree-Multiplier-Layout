magic
tech scmos
timestamp 1199203594
<< ab >>
rect 0 0 136 80
<< nwell >>
rect -5 36 141 88
<< pwell >>
rect -5 -8 141 36
<< poly >>
rect 20 70 22 74
rect 30 70 32 74
rect 45 70 47 74
rect 55 70 57 74
rect 85 70 87 74
rect 95 70 97 74
rect 105 70 107 74
rect 115 70 117 74
rect 125 70 127 74
rect 71 62 77 64
rect 71 60 73 62
rect 75 60 77 62
rect 65 55 67 60
rect 71 58 77 60
rect 75 55 77 58
rect 20 39 22 42
rect 30 39 32 42
rect 45 39 47 42
rect 55 39 57 42
rect 9 37 51 39
rect 9 35 11 37
rect 13 35 21 37
rect 9 33 21 35
rect 9 30 11 33
rect 19 30 21 33
rect 39 30 41 37
rect 49 30 51 37
rect 55 37 61 39
rect 55 35 57 37
rect 59 35 61 37
rect 65 37 67 42
rect 75 37 77 42
rect 85 39 87 42
rect 95 39 97 42
rect 105 39 107 42
rect 85 37 97 39
rect 101 37 107 39
rect 65 35 80 37
rect 55 33 61 35
rect 59 30 61 33
rect 66 30 68 35
rect 78 30 80 35
rect 85 35 87 37
rect 89 35 91 37
rect 85 33 91 35
rect 101 35 103 37
rect 105 35 107 37
rect 101 33 107 35
rect 115 39 117 42
rect 125 39 127 42
rect 115 37 127 39
rect 115 35 123 37
rect 125 35 127 37
rect 115 33 127 35
rect 85 30 87 33
rect 115 30 117 33
rect 125 30 127 33
rect 9 15 11 19
rect 19 8 21 13
rect 39 11 41 16
rect 49 11 51 16
rect 115 12 117 16
rect 125 12 127 16
rect 59 6 61 11
rect 66 6 68 11
rect 78 6 80 11
rect 85 6 87 11
<< ndif >>
rect 2 23 9 30
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 19 19 26
rect 14 13 19 19
rect 21 17 28 30
rect 21 15 24 17
rect 26 15 28 17
rect 32 28 39 30
rect 32 26 34 28
rect 36 26 39 28
rect 32 21 39 26
rect 32 19 34 21
rect 36 19 39 21
rect 32 16 39 19
rect 41 28 49 30
rect 41 26 44 28
rect 46 26 49 28
rect 41 16 49 26
rect 51 28 59 30
rect 51 26 54 28
rect 56 26 59 28
rect 51 21 59 26
rect 51 19 54 21
rect 56 19 59 21
rect 51 16 59 19
rect 21 13 28 15
rect 54 11 59 16
rect 61 11 66 30
rect 68 11 78 30
rect 80 11 85 30
rect 87 23 92 30
rect 87 21 94 23
rect 87 19 90 21
rect 92 19 94 21
rect 87 17 94 19
rect 108 20 115 30
rect 108 18 110 20
rect 112 18 115 20
rect 87 11 92 17
rect 108 16 115 18
rect 117 28 125 30
rect 117 26 120 28
rect 122 26 125 28
rect 117 21 125 26
rect 117 19 120 21
rect 122 19 125 21
rect 117 16 125 19
rect 127 20 134 30
rect 127 18 130 20
rect 132 18 134 20
rect 127 16 134 18
rect 70 9 72 11
rect 74 9 76 11
rect 70 7 76 9
<< pdif >>
rect 13 68 20 70
rect 13 66 15 68
rect 17 66 20 68
rect 13 61 20 66
rect 13 59 15 61
rect 17 59 20 61
rect 13 42 20 59
rect 22 53 30 70
rect 22 51 25 53
rect 27 51 30 53
rect 22 46 30 51
rect 22 44 25 46
rect 27 44 30 46
rect 22 42 30 44
rect 32 68 45 70
rect 32 66 37 68
rect 39 66 45 68
rect 32 61 45 66
rect 32 59 37 61
rect 39 59 45 61
rect 32 42 45 59
rect 47 61 55 70
rect 47 59 50 61
rect 52 59 55 61
rect 47 54 55 59
rect 47 52 50 54
rect 52 52 55 54
rect 47 42 55 52
rect 57 55 62 70
rect 80 55 85 70
rect 57 53 65 55
rect 57 51 60 53
rect 62 51 65 53
rect 57 46 65 51
rect 57 44 60 46
rect 62 44 65 46
rect 57 42 65 44
rect 67 46 75 55
rect 67 44 70 46
rect 72 44 75 46
rect 67 42 75 44
rect 77 53 85 55
rect 77 51 80 53
rect 82 51 85 53
rect 77 42 85 51
rect 87 62 95 70
rect 87 60 90 62
rect 92 60 95 62
rect 87 46 95 60
rect 87 44 90 46
rect 92 44 95 46
rect 87 42 95 44
rect 97 61 105 70
rect 97 59 100 61
rect 102 59 105 61
rect 97 54 105 59
rect 97 52 100 54
rect 102 52 105 54
rect 97 42 105 52
rect 107 53 115 70
rect 107 51 110 53
rect 112 51 115 53
rect 107 46 115 51
rect 107 44 110 46
rect 112 44 115 46
rect 107 42 115 44
rect 117 68 125 70
rect 117 66 120 68
rect 122 66 125 68
rect 117 61 125 66
rect 117 59 120 61
rect 122 59 125 61
rect 117 42 125 59
rect 127 55 132 70
rect 127 53 134 55
rect 127 51 130 53
rect 132 51 134 53
rect 127 46 134 51
rect 127 44 130 46
rect 132 44 134 46
rect 127 42 134 44
<< alu1 >>
rect -2 81 138 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 138 81
rect -2 68 138 79
rect 98 61 103 63
rect 98 59 100 61
rect 102 59 103 61
rect 98 54 103 59
rect 58 53 100 54
rect 58 51 60 53
rect 62 51 80 53
rect 82 52 100 53
rect 102 52 103 54
rect 82 51 103 52
rect 58 50 103 51
rect 2 39 6 47
rect 58 46 63 50
rect 34 44 60 46
rect 62 44 63 46
rect 34 42 63 44
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 34 29 38 42
rect 32 28 38 29
rect 32 26 34 28
rect 36 26 38 28
rect 32 22 38 26
rect 121 37 134 39
rect 121 35 123 37
rect 125 35 134 37
rect 121 34 134 35
rect 53 28 57 30
rect 53 26 54 28
rect 56 26 57 28
rect 53 22 57 26
rect 32 21 95 22
rect 32 19 34 21
rect 36 19 54 21
rect 56 19 90 21
rect 92 19 95 21
rect 32 18 95 19
rect 130 25 134 34
rect -2 11 138 12
rect -2 9 72 11
rect 74 9 138 11
rect -2 1 138 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 138 1
rect -2 -2 138 -1
<< ptie >>
rect 0 1 136 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 136 1
rect 0 -3 136 -1
<< ntie >>
rect 0 81 136 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 136 81
rect 0 77 136 79
<< nmos >>
rect 9 19 11 30
rect 19 13 21 30
rect 39 16 41 30
rect 49 16 51 30
rect 59 11 61 30
rect 66 11 68 30
rect 78 11 80 30
rect 85 11 87 30
rect 115 16 117 30
rect 125 16 127 30
<< pmos >>
rect 20 42 22 70
rect 30 42 32 70
rect 45 42 47 70
rect 55 42 57 70
rect 65 42 67 55
rect 75 42 77 55
rect 85 42 87 70
rect 95 42 97 70
rect 105 42 107 70
rect 115 42 117 70
rect 125 42 127 70
<< polyct0 >>
rect 73 60 75 62
rect 57 35 59 37
rect 87 35 89 37
rect 103 35 105 37
<< polyct1 >>
rect 11 35 13 37
rect 123 35 125 37
<< ndifct0 >>
rect 4 21 6 23
rect 14 26 16 28
rect 24 15 26 17
rect 44 26 46 28
rect 110 18 112 20
rect 120 26 122 28
rect 120 19 122 21
rect 130 18 132 20
<< ndifct1 >>
rect 34 26 36 28
rect 34 19 36 21
rect 54 26 56 28
rect 54 19 56 21
rect 90 19 92 21
rect 72 9 74 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
<< pdifct0 >>
rect 15 66 17 68
rect 15 59 17 61
rect 25 51 27 53
rect 25 44 27 46
rect 37 66 39 68
rect 37 59 39 61
rect 50 59 52 61
rect 50 52 52 54
rect 70 44 72 46
rect 90 60 92 62
rect 90 44 92 46
rect 110 51 112 53
rect 110 44 112 46
rect 120 66 122 68
rect 120 59 122 61
rect 130 51 132 53
rect 130 44 132 46
<< pdifct1 >>
rect 60 51 62 53
rect 60 44 62 46
rect 80 51 82 53
rect 100 59 102 61
rect 100 52 102 54
<< alu0 >>
rect 14 66 15 68
rect 17 66 18 68
rect 14 61 18 66
rect 14 59 15 61
rect 17 59 18 61
rect 14 57 18 59
rect 35 66 37 68
rect 39 66 41 68
rect 35 61 41 66
rect 119 66 120 68
rect 122 66 123 68
rect 35 59 37 61
rect 39 59 41 61
rect 35 58 41 59
rect 49 62 94 63
rect 49 61 73 62
rect 49 59 50 61
rect 52 60 73 61
rect 75 60 90 62
rect 92 60 94 62
rect 52 59 94 60
rect 49 54 53 59
rect 119 61 123 66
rect 119 59 120 61
rect 122 59 123 61
rect 119 57 123 59
rect 23 53 50 54
rect 23 51 25 53
rect 27 52 50 53
rect 52 52 53 54
rect 27 51 53 52
rect 23 50 53 51
rect 108 53 113 55
rect 108 51 110 53
rect 112 51 113 53
rect 23 46 28 50
rect 108 47 113 51
rect 129 53 134 55
rect 129 51 130 53
rect 132 51 134 53
rect 129 47 134 51
rect 23 44 25 46
rect 27 44 28 46
rect 23 42 28 44
rect 68 46 74 47
rect 68 44 70 46
rect 72 44 74 46
rect 23 29 27 42
rect 68 38 74 44
rect 88 46 94 47
rect 108 46 134 47
rect 88 44 90 46
rect 92 44 103 46
rect 88 42 103 44
rect 108 44 110 46
rect 112 44 130 46
rect 132 44 134 46
rect 108 43 134 44
rect 99 38 103 42
rect 12 28 27 29
rect 12 26 14 28
rect 16 26 27 28
rect 12 25 27 26
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 12 7 21
rect 42 37 93 38
rect 42 35 57 37
rect 59 35 87 37
rect 89 35 93 37
rect 42 34 93 35
rect 99 37 107 38
rect 99 35 103 37
rect 105 35 107 37
rect 99 34 107 35
rect 42 28 48 34
rect 89 30 93 34
rect 112 30 116 43
rect 42 26 44 28
rect 46 26 48 28
rect 42 25 48 26
rect 89 28 123 30
rect 89 26 120 28
rect 122 26 123 28
rect 23 17 27 19
rect 109 20 113 22
rect 109 18 110 20
rect 112 18 113 20
rect 23 15 24 17
rect 26 15 27 17
rect 23 12 27 15
rect 109 12 113 18
rect 119 21 123 26
rect 119 19 120 21
rect 122 19 123 21
rect 119 17 123 19
rect 128 20 134 21
rect 128 18 130 20
rect 132 18 134 20
rect 128 12 134 18
<< labels >>
rlabel alu0 19 27 19 27 6 bn
rlabel alu0 45 31 45 31 6 an
rlabel alu0 51 56 51 56 6 bn
rlabel alu0 38 52 38 52 6 bn
rlabel alu0 25 48 25 48 6 bn
rlabel alu0 71 40 71 40 6 an
rlabel alu0 67 36 67 36 6 an
rlabel alu0 95 44 95 44 6 bn
rlabel alu0 71 61 71 61 6 bn
rlabel alu0 121 23 121 23 6 an
rlabel alu0 121 45 121 45 6 an
rlabel alu0 103 36 103 36 6 bn
rlabel alu0 131 49 131 49 6 an
rlabel alu0 110 49 110 49 6 an
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 40 4 40 6 b
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 36 28 36 28 6 z
rlabel alu1 44 44 44 44 6 z
rlabel alu1 52 44 52 44 6 z
rlabel alu1 60 44 60 44 6 z
rlabel alu1 68 6 68 6 6 vss
rlabel alu1 76 20 76 20 6 z
rlabel alu1 84 20 84 20 6 z
rlabel alu1 92 20 92 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 92 52 92 52 6 z
rlabel alu1 100 56 100 56 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 68 74 68 74 6 vdd
rlabel polyct1 124 36 124 36 6 a
rlabel alu1 132 32 132 32 6 a
<< end >>
