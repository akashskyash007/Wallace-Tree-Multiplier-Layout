magic
tech scmos
timestamp 1199203343
<< ab >>
rect 0 0 16 80
<< nwell >>
rect -5 36 21 88
<< pwell >>
rect -5 -8 21 36
<< alu1 >>
rect -2 81 18 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 18 81
rect -2 68 18 79
rect -2 1 18 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 18 1
rect -2 -2 18 -1
<< ptie >>
rect 0 1 16 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 16 1
rect 0 -3 16 -1
<< ntie >>
rect 0 81 16 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 16 81
rect 0 77 16 79
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
<< labels >>
rlabel alu1 8 6 8 6 6 vss
rlabel alu1 8 74 8 74 6 vdd
<< end >>
