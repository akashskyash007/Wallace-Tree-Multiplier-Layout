magic
tech scmos
timestamp 1199203251
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 24 65 26 70
rect 31 65 33 70
rect 38 65 40 70
rect 13 57 15 63
rect 13 42 15 45
rect 9 40 15 42
rect 9 38 11 40
rect 13 38 15 40
rect 9 36 15 38
rect 9 18 11 36
rect 24 35 26 40
rect 19 33 26 35
rect 19 31 21 33
rect 23 32 26 33
rect 23 31 25 32
rect 19 29 25 31
rect 19 18 21 29
rect 31 27 33 40
rect 38 37 40 40
rect 38 35 47 37
rect 41 33 43 35
rect 45 33 47 35
rect 41 31 47 33
rect 29 25 36 27
rect 29 23 32 25
rect 34 23 36 25
rect 29 21 36 23
rect 29 18 31 21
rect 41 18 43 31
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 41 7 43 12
<< ndif >>
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 16 19 18
rect 11 14 14 16
rect 16 14 19 16
rect 11 12 19 14
rect 21 16 29 18
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 31 12 41 18
rect 43 16 50 18
rect 43 14 46 16
rect 48 14 50 16
rect 43 12 50 14
rect 33 7 39 12
rect 33 5 35 7
rect 37 5 39 7
rect 33 3 39 5
<< pdif >>
rect 17 63 24 65
rect 17 61 19 63
rect 21 61 24 63
rect 17 57 24 61
rect 6 55 13 57
rect 6 53 8 55
rect 10 53 13 55
rect 6 51 13 53
rect 8 45 13 51
rect 15 45 24 57
rect 17 40 24 45
rect 26 40 31 65
rect 33 40 38 65
rect 40 60 45 65
rect 40 58 47 60
rect 40 56 43 58
rect 45 56 47 58
rect 40 54 47 56
rect 40 40 45 54
<< alu1 >>
rect -2 67 58 72
rect -2 65 5 67
rect 7 65 58 67
rect -2 64 58 65
rect 2 55 15 58
rect 2 53 8 55
rect 10 53 15 55
rect 2 52 15 53
rect 2 17 6 52
rect 34 45 46 51
rect 26 35 30 43
rect 42 35 46 45
rect 17 33 30 35
rect 17 31 21 33
rect 23 31 30 33
rect 17 30 30 31
rect 34 26 38 35
rect 42 33 43 35
rect 45 33 46 35
rect 42 31 46 33
rect 30 25 47 26
rect 30 23 32 25
rect 34 23 47 25
rect 30 22 47 23
rect 2 16 8 17
rect 2 14 4 16
rect 6 14 8 16
rect 2 13 8 14
rect -2 7 58 8
rect -2 5 35 7
rect 37 5 58 7
rect -2 0 58 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 12 11 18
rect 19 12 21 18
rect 29 12 31 18
rect 41 12 43 18
<< pmos >>
rect 13 45 15 57
rect 24 40 26 65
rect 31 40 33 65
rect 38 40 40 65
<< polyct0 >>
rect 11 38 13 40
<< polyct1 >>
rect 21 31 23 33
rect 43 33 45 35
rect 32 23 34 25
<< ndifct0 >>
rect 14 14 16 16
rect 24 14 26 16
rect 46 14 48 16
<< ndifct1 >>
rect 4 14 6 16
rect 35 5 37 7
<< ntiect1 >>
rect 5 65 7 67
<< pdifct0 >>
rect 19 61 21 63
rect 43 56 45 58
<< pdifct1 >>
rect 8 53 10 55
<< alu0 >>
rect 18 63 22 64
rect 18 61 19 63
rect 21 61 22 63
rect 18 59 22 61
rect 26 58 47 59
rect 26 56 43 58
rect 45 56 47 58
rect 26 55 47 56
rect 26 51 30 55
rect 18 47 30 51
rect 18 44 22 47
rect 10 40 22 44
rect 10 38 11 40
rect 13 38 14 40
rect 10 25 14 38
rect 10 21 26 25
rect 22 17 26 21
rect 12 16 18 17
rect 12 14 14 16
rect 16 14 18 16
rect 12 8 18 14
rect 22 16 50 17
rect 22 14 24 16
rect 26 14 46 16
rect 48 14 50 16
rect 22 13 50 14
<< labels >>
rlabel alu0 12 32 12 32 6 zn
rlabel alu0 36 15 36 15 6 zn
rlabel alu0 36 57 36 57 6 zn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 32 20 32 6 a
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 28 36 28 6 b
rlabel alu1 28 40 28 40 6 a
rlabel alu1 36 48 36 48 6 c
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 24 44 24 6 b
rlabel alu1 44 44 44 44 6 c
<< end >>
