magic
tech scmos
timestamp 1199543931
<< ab >>
rect 0 0 240 100
<< nwell >>
rect -5 48 245 105
<< pwell >>
rect -5 -5 245 48
<< poly >>
rect 119 94 121 98
rect 155 94 157 98
rect 167 94 169 98
rect 179 94 181 98
rect 191 94 193 98
rect 203 94 205 98
rect 215 94 217 98
rect 227 94 229 98
rect 11 85 13 89
rect 23 85 25 89
rect 31 85 33 89
rect 49 85 51 89
rect 57 85 59 89
rect 83 86 85 90
rect 95 85 97 89
rect 11 51 13 65
rect 23 63 25 66
rect 17 61 25 63
rect 17 59 19 61
rect 21 59 25 61
rect 17 57 25 59
rect 31 53 33 66
rect 49 63 51 66
rect 57 63 59 66
rect 83 63 85 66
rect 131 86 133 90
rect 119 73 121 76
rect 115 71 121 73
rect 115 69 117 71
rect 119 69 121 71
rect 115 67 121 69
rect 143 85 145 89
rect 47 61 53 63
rect 47 59 49 61
rect 51 59 53 61
rect 47 57 53 59
rect 57 61 63 63
rect 57 59 59 61
rect 61 59 63 61
rect 57 57 63 59
rect 83 61 91 63
rect 83 59 87 61
rect 89 59 91 61
rect 83 57 91 59
rect 27 51 33 53
rect 77 51 83 53
rect 95 51 97 65
rect 131 63 133 66
rect 155 73 157 76
rect 155 71 163 73
rect 155 69 159 71
rect 161 69 163 71
rect 155 67 163 69
rect 127 61 133 63
rect 127 59 129 61
rect 131 59 133 61
rect 127 57 133 59
rect 127 51 133 53
rect 143 51 145 65
rect 167 63 169 75
rect 161 61 169 63
rect 161 59 163 61
rect 165 59 169 61
rect 161 57 169 59
rect 179 51 181 75
rect 191 73 193 76
rect 185 71 193 73
rect 185 69 187 71
rect 189 69 193 71
rect 185 67 193 69
rect 203 53 205 75
rect 203 51 211 53
rect 11 49 29 51
rect 31 49 51 51
rect 11 25 13 49
rect 27 47 33 49
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 17 31 25 33
rect 17 29 19 31
rect 21 29 25 31
rect 17 27 25 29
rect 23 24 25 27
rect 31 24 33 37
rect 49 24 51 49
rect 77 49 79 51
rect 81 49 129 51
rect 131 49 193 51
rect 77 47 83 49
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 57 27 63 29
rect 83 31 91 33
rect 83 29 87 31
rect 89 29 91 31
rect 83 27 91 29
rect 57 24 59 27
rect 83 24 85 27
rect 95 25 97 49
rect 127 47 133 49
rect 101 41 107 43
rect 137 41 145 43
rect 179 41 187 43
rect 101 39 103 41
rect 105 39 139 41
rect 141 39 183 41
rect 185 39 187 41
rect 101 37 107 39
rect 137 37 145 39
rect 117 31 123 33
rect 117 29 119 31
rect 121 29 123 31
rect 117 27 123 29
rect 127 31 133 33
rect 127 29 129 31
rect 131 29 133 31
rect 127 27 133 29
rect 11 11 13 15
rect 23 11 25 15
rect 31 11 33 15
rect 49 11 51 15
rect 57 11 59 15
rect 119 24 121 27
rect 131 24 133 27
rect 143 25 145 37
rect 179 37 187 39
rect 161 31 169 33
rect 161 29 163 31
rect 165 29 169 31
rect 161 27 169 29
rect 83 10 85 14
rect 95 11 97 15
rect 119 11 121 15
rect 131 11 133 15
rect 143 11 145 15
rect 155 21 163 23
rect 155 19 159 21
rect 161 19 163 21
rect 155 17 163 19
rect 155 14 157 17
rect 167 15 169 27
rect 179 25 181 37
rect 191 25 193 49
rect 203 49 207 51
rect 209 49 211 51
rect 203 47 211 49
rect 215 43 217 55
rect 227 43 229 55
rect 205 41 229 43
rect 205 39 207 41
rect 209 39 229 41
rect 205 37 229 39
rect 203 31 211 33
rect 203 29 207 31
rect 209 29 211 31
rect 203 27 211 29
rect 203 24 205 27
rect 215 25 217 37
rect 227 25 229 37
rect 179 11 181 15
rect 191 11 193 15
rect 203 11 205 15
rect 155 2 157 6
rect 167 2 169 6
rect 215 2 217 6
rect 227 2 229 6
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 24 18 25
rect 37 31 47 33
rect 37 29 39 31
rect 41 29 47 31
rect 37 24 47 29
rect 90 24 95 25
rect 13 15 23 24
rect 25 15 31 24
rect 33 15 49 24
rect 51 15 57 24
rect 59 15 67 24
rect 15 11 21 15
rect 61 11 67 15
rect 75 21 83 24
rect 75 19 77 21
rect 79 19 83 21
rect 75 14 83 19
rect 85 15 95 24
rect 97 21 105 25
rect 138 24 143 25
rect 97 19 101 21
rect 103 19 105 21
rect 97 15 105 19
rect 111 15 119 24
rect 121 15 131 24
rect 133 21 143 24
rect 133 19 137 21
rect 139 19 143 21
rect 133 15 143 19
rect 145 15 153 25
rect 85 14 93 15
rect 15 9 17 11
rect 19 9 21 11
rect 61 9 63 11
rect 65 9 67 11
rect 87 11 93 14
rect 111 11 117 15
rect 147 14 153 15
rect 171 21 179 25
rect 171 19 173 21
rect 175 19 179 21
rect 171 15 179 19
rect 181 21 191 25
rect 181 19 185 21
rect 187 19 191 21
rect 181 15 191 19
rect 193 24 198 25
rect 210 24 215 25
rect 193 15 203 24
rect 205 21 215 24
rect 205 19 209 21
rect 211 19 215 21
rect 205 15 215 19
rect 162 14 167 15
rect 15 7 21 9
rect 61 7 67 9
rect 87 9 89 11
rect 91 9 93 11
rect 87 7 93 9
rect 111 9 113 11
rect 115 9 117 11
rect 111 7 117 9
rect 147 6 155 14
rect 157 11 167 14
rect 157 9 161 11
rect 163 9 167 11
rect 157 6 167 9
rect 169 6 177 15
rect 207 11 215 15
rect 207 9 209 11
rect 211 9 215 11
rect 207 6 215 9
rect 217 21 227 25
rect 217 19 221 21
rect 223 19 227 21
rect 217 6 227 19
rect 229 21 237 25
rect 229 19 233 21
rect 235 19 237 21
rect 229 11 237 19
rect 229 9 233 11
rect 235 9 237 11
rect 229 6 237 9
<< pdif >>
rect 15 91 21 93
rect 61 91 67 93
rect 15 89 17 91
rect 19 89 21 91
rect 61 89 63 91
rect 65 89 67 91
rect 87 91 93 93
rect 15 85 21 89
rect 61 85 67 89
rect 87 89 89 91
rect 91 89 93 91
rect 111 91 119 94
rect 111 89 113 91
rect 115 89 119 91
rect 87 86 93 89
rect 3 71 11 85
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 66 23 85
rect 25 66 31 85
rect 33 71 49 85
rect 33 69 39 71
rect 41 69 49 71
rect 33 66 49 69
rect 51 66 57 85
rect 59 66 67 85
rect 75 71 83 86
rect 75 69 77 71
rect 79 69 83 71
rect 75 66 83 69
rect 85 85 93 86
rect 85 66 95 85
rect 13 65 18 66
rect 90 65 95 66
rect 97 71 105 85
rect 111 76 119 89
rect 121 86 129 94
rect 121 76 131 86
rect 97 69 101 71
rect 103 69 105 71
rect 97 65 105 69
rect 123 66 131 76
rect 133 85 141 86
rect 147 85 155 94
rect 133 71 143 85
rect 133 69 137 71
rect 139 69 143 71
rect 133 66 143 69
rect 138 65 143 66
rect 145 76 155 85
rect 157 91 167 94
rect 157 89 161 91
rect 163 89 167 91
rect 157 76 167 89
rect 145 65 153 76
rect 162 75 167 76
rect 169 81 179 94
rect 169 79 173 81
rect 175 79 179 81
rect 169 75 179 79
rect 181 81 191 94
rect 181 79 185 81
rect 187 79 191 81
rect 181 76 191 79
rect 193 76 203 94
rect 181 75 186 76
rect 198 75 203 76
rect 205 91 215 94
rect 205 89 209 91
rect 211 89 215 91
rect 205 81 215 89
rect 205 79 209 81
rect 211 79 215 81
rect 205 75 215 79
rect 207 71 215 75
rect 207 69 209 71
rect 211 69 215 71
rect 207 61 215 69
rect 207 59 209 61
rect 211 59 215 61
rect 207 55 215 59
rect 217 81 227 94
rect 217 79 221 81
rect 223 79 227 81
rect 217 71 227 79
rect 217 69 221 71
rect 223 69 227 71
rect 217 61 227 69
rect 217 59 221 61
rect 223 59 227 61
rect 217 55 227 59
rect 229 91 237 94
rect 229 89 233 91
rect 235 89 237 91
rect 229 81 237 89
rect 229 79 233 81
rect 235 79 237 81
rect 229 71 237 79
rect 229 69 233 71
rect 235 69 237 71
rect 229 61 237 69
rect 229 59 233 61
rect 235 59 237 61
rect 229 55 237 59
<< alu1 >>
rect -2 95 242 100
rect -2 93 29 95
rect 31 93 49 95
rect 51 93 242 95
rect -2 91 242 93
rect -2 89 17 91
rect 19 89 63 91
rect 65 89 89 91
rect 91 89 113 91
rect 115 89 161 91
rect 163 89 209 91
rect 211 89 233 91
rect 235 89 242 91
rect -2 88 242 89
rect 4 71 8 73
rect 4 69 5 71
rect 7 69 8 71
rect 4 22 8 69
rect 18 61 22 83
rect 18 59 19 61
rect 21 59 22 61
rect 18 31 22 59
rect 28 51 32 83
rect 28 49 29 51
rect 31 49 32 51
rect 28 47 32 49
rect 38 78 122 82
rect 38 71 42 78
rect 38 69 39 71
rect 41 69 42 71
rect 18 29 19 31
rect 21 29 22 31
rect 18 27 22 29
rect 28 41 32 43
rect 28 39 29 41
rect 31 39 32 41
rect 28 22 32 39
rect 38 31 42 69
rect 38 29 39 31
rect 41 29 42 31
rect 38 27 42 29
rect 48 61 52 63
rect 48 59 49 61
rect 51 59 52 61
rect 48 22 52 59
rect 4 21 52 22
rect 4 19 5 21
rect 7 19 52 21
rect 4 18 52 19
rect 58 61 62 73
rect 58 59 59 61
rect 61 59 62 61
rect 58 31 62 59
rect 58 29 59 31
rect 61 29 62 31
rect 4 17 8 18
rect 58 17 62 29
rect 76 71 80 73
rect 76 69 77 71
rect 79 69 80 71
rect 76 52 80 69
rect 88 62 92 73
rect 85 61 92 62
rect 85 59 87 61
rect 89 59 92 61
rect 85 58 92 59
rect 76 51 83 52
rect 76 49 79 51
rect 81 49 83 51
rect 76 48 83 49
rect 76 21 80 48
rect 88 32 92 58
rect 85 31 92 32
rect 85 29 87 31
rect 89 29 92 31
rect 85 28 92 29
rect 76 19 77 21
rect 79 19 80 21
rect 76 17 80 19
rect 88 17 92 28
rect 100 71 104 73
rect 118 72 122 78
rect 172 81 176 83
rect 172 79 173 81
rect 175 79 176 81
rect 172 72 176 79
rect 183 81 200 82
rect 183 79 185 81
rect 187 79 200 81
rect 183 78 200 79
rect 100 69 101 71
rect 103 69 104 71
rect 100 42 104 69
rect 115 71 122 72
rect 115 69 117 71
rect 119 69 122 71
rect 115 68 122 69
rect 135 71 152 72
rect 135 69 137 71
rect 139 69 152 71
rect 135 68 152 69
rect 157 71 176 72
rect 157 69 159 71
rect 161 69 176 71
rect 157 68 176 69
rect 100 41 107 42
rect 100 39 103 41
rect 105 39 107 41
rect 100 38 107 39
rect 100 21 104 38
rect 118 31 122 68
rect 148 62 152 68
rect 127 61 142 62
rect 127 59 129 61
rect 131 59 142 61
rect 127 58 142 59
rect 118 29 119 31
rect 121 29 122 31
rect 118 27 122 29
rect 128 51 132 53
rect 128 49 129 51
rect 131 49 132 51
rect 128 31 132 49
rect 138 41 142 58
rect 138 39 139 41
rect 141 39 142 41
rect 138 37 142 39
rect 148 61 167 62
rect 148 59 163 61
rect 165 59 167 61
rect 148 58 167 59
rect 128 29 129 31
rect 131 29 132 31
rect 128 27 132 29
rect 148 32 152 58
rect 148 31 167 32
rect 148 29 163 31
rect 165 29 167 31
rect 148 28 167 29
rect 148 22 152 28
rect 172 22 176 68
rect 184 71 191 72
rect 184 69 187 71
rect 189 69 191 71
rect 184 68 191 69
rect 184 42 188 68
rect 181 41 188 42
rect 181 39 183 41
rect 185 39 188 41
rect 181 38 188 39
rect 196 42 200 78
rect 208 81 212 88
rect 208 79 209 81
rect 211 79 212 81
rect 208 71 212 79
rect 208 69 209 71
rect 211 69 212 71
rect 208 61 212 69
rect 208 59 209 61
rect 211 59 212 61
rect 208 57 212 59
rect 218 82 222 83
rect 218 81 225 82
rect 218 79 221 81
rect 223 79 225 81
rect 218 78 225 79
rect 232 81 236 88
rect 232 79 233 81
rect 235 79 236 81
rect 218 72 222 78
rect 218 71 225 72
rect 218 69 221 71
rect 223 69 225 71
rect 218 68 225 69
rect 232 71 236 79
rect 232 69 233 71
rect 235 69 236 71
rect 218 62 222 68
rect 218 61 225 62
rect 218 59 221 61
rect 223 59 225 61
rect 218 58 225 59
rect 232 61 236 69
rect 232 59 233 61
rect 235 59 236 61
rect 218 52 222 58
rect 232 57 236 59
rect 205 51 224 52
rect 205 49 207 51
rect 209 49 224 51
rect 205 48 224 49
rect 196 41 211 42
rect 196 39 207 41
rect 209 39 211 41
rect 196 38 211 39
rect 196 22 200 38
rect 218 32 222 48
rect 205 31 224 32
rect 205 29 207 31
rect 209 29 224 31
rect 205 28 224 29
rect 100 19 101 21
rect 103 19 104 21
rect 100 17 104 19
rect 135 21 152 22
rect 135 19 137 21
rect 139 19 152 21
rect 135 18 152 19
rect 157 21 176 22
rect 157 19 159 21
rect 161 19 173 21
rect 175 19 176 21
rect 157 18 176 19
rect 183 21 200 22
rect 183 19 185 21
rect 187 19 200 21
rect 183 18 200 19
rect 208 21 212 23
rect 208 19 209 21
rect 211 19 212 21
rect 172 17 176 18
rect 208 12 212 19
rect 218 22 222 28
rect 218 21 225 22
rect 218 19 221 21
rect 223 19 225 21
rect 218 18 225 19
rect 232 21 236 23
rect 232 19 233 21
rect 235 19 236 21
rect 218 17 222 18
rect 232 12 236 19
rect -2 11 242 12
rect -2 9 17 11
rect 19 9 63 11
rect 65 9 89 11
rect 91 9 113 11
rect 115 9 161 11
rect 163 9 209 11
rect 211 9 233 11
rect 235 9 242 11
rect -2 7 242 9
rect -2 5 29 7
rect 31 5 49 7
rect 51 5 125 7
rect 127 5 137 7
rect 139 5 185 7
rect 187 5 197 7
rect 199 5 242 7
rect -2 0 242 5
<< ptie >>
rect 27 7 53 9
rect 123 7 141 9
rect 27 5 29 7
rect 31 5 49 7
rect 51 5 53 7
rect 27 3 53 5
rect 123 5 125 7
rect 127 5 137 7
rect 139 5 141 7
rect 183 7 201 9
rect 123 3 141 5
rect 183 5 185 7
rect 187 5 197 7
rect 199 5 201 7
rect 183 3 201 5
<< ntie >>
rect 27 95 53 97
rect 27 93 29 95
rect 31 93 49 95
rect 51 93 53 95
rect 27 91 53 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 24
rect 31 15 33 24
rect 49 15 51 24
rect 57 15 59 24
rect 83 14 85 24
rect 95 15 97 25
rect 119 15 121 24
rect 131 15 133 24
rect 143 15 145 25
rect 179 15 181 25
rect 191 15 193 25
rect 203 15 205 24
rect 155 6 157 14
rect 167 6 169 15
rect 215 6 217 25
rect 227 6 229 25
<< pmos >>
rect 11 65 13 85
rect 23 66 25 85
rect 31 66 33 85
rect 49 66 51 85
rect 57 66 59 85
rect 83 66 85 86
rect 95 65 97 85
rect 119 76 121 94
rect 131 66 133 86
rect 143 65 145 85
rect 155 76 157 94
rect 167 75 169 94
rect 179 75 181 94
rect 191 76 193 94
rect 203 75 205 94
rect 215 55 217 94
rect 227 55 229 94
<< polyct1 >>
rect 19 59 21 61
rect 117 69 119 71
rect 49 59 51 61
rect 59 59 61 61
rect 87 59 89 61
rect 159 69 161 71
rect 129 59 131 61
rect 163 59 165 61
rect 187 69 189 71
rect 29 49 31 51
rect 29 39 31 41
rect 19 29 21 31
rect 79 49 81 51
rect 129 49 131 51
rect 59 29 61 31
rect 87 29 89 31
rect 103 39 105 41
rect 139 39 141 41
rect 183 39 185 41
rect 119 29 121 31
rect 129 29 131 31
rect 163 29 165 31
rect 159 19 161 21
rect 207 49 209 51
rect 207 39 209 41
rect 207 29 209 31
<< ndifct1 >>
rect 5 19 7 21
rect 39 29 41 31
rect 77 19 79 21
rect 101 19 103 21
rect 137 19 139 21
rect 17 9 19 11
rect 63 9 65 11
rect 173 19 175 21
rect 185 19 187 21
rect 209 19 211 21
rect 89 9 91 11
rect 113 9 115 11
rect 161 9 163 11
rect 209 9 211 11
rect 221 19 223 21
rect 233 19 235 21
rect 233 9 235 11
<< ntiect1 >>
rect 29 93 31 95
rect 49 93 51 95
<< ptiect1 >>
rect 29 5 31 7
rect 49 5 51 7
rect 125 5 127 7
rect 137 5 139 7
rect 185 5 187 7
rect 197 5 199 7
<< pdifct1 >>
rect 17 89 19 91
rect 63 89 65 91
rect 89 89 91 91
rect 113 89 115 91
rect 5 69 7 71
rect 39 69 41 71
rect 77 69 79 71
rect 101 69 103 71
rect 137 69 139 71
rect 161 89 163 91
rect 173 79 175 81
rect 185 79 187 81
rect 209 89 211 91
rect 209 79 211 81
rect 209 69 211 71
rect 209 59 211 61
rect 221 79 223 81
rect 221 69 223 71
rect 221 59 223 61
rect 233 89 235 91
rect 233 79 235 81
rect 233 69 235 71
rect 233 59 235 61
<< labels >>
rlabel alu1 20 55 20 55 6 i0
rlabel alu1 30 65 30 65 6 cmd
rlabel alu1 90 45 90 45 6 ck
rlabel alu1 60 45 60 45 6 i1
rlabel alu1 120 6 120 6 6 vss
rlabel alu1 120 94 120 94 6 vdd
rlabel alu1 210 30 210 30 6 q
rlabel alu1 220 50 220 50 6 q
rlabel alu1 210 50 210 50 6 q
<< end >>
