magic
tech scmos
timestamp 1199472707
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -2 48 62 104
<< pwell >>
rect -2 -4 62 48
<< alu1 >>
rect -2 95 62 100
rect -2 93 5 95
rect 7 93 14 95
rect 16 93 24 95
rect 26 93 34 95
rect 36 93 44 95
rect 46 93 53 95
rect 55 93 62 95
rect -2 88 62 93
rect -2 7 62 12
rect -2 5 5 7
rect 7 5 14 7
rect 16 5 24 7
rect 26 5 34 7
rect 36 5 44 7
rect 46 5 53 7
rect 55 5 62 7
rect -2 0 62 5
<< ptie >>
rect 3 7 57 39
rect 3 5 5 7
rect 7 5 14 7
rect 16 5 24 7
rect 26 5 34 7
rect 36 5 44 7
rect 46 5 53 7
rect 55 5 57 7
rect 3 3 57 5
<< ntie >>
rect 3 95 57 97
rect 3 93 5 95
rect 7 93 14 95
rect 16 93 24 95
rect 26 93 34 95
rect 36 93 44 95
rect 46 93 53 95
rect 55 93 57 95
rect 3 55 57 93
<< ntiect1 >>
rect 5 93 7 95
rect 14 93 16 95
rect 24 93 26 95
rect 34 93 36 95
rect 44 93 46 95
rect 53 93 55 95
<< ptiect1 >>
rect 5 5 7 7
rect 14 5 16 7
rect 24 5 26 7
rect 34 5 36 7
rect 44 5 46 7
rect 53 5 55 7
<< labels >>
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 30 94 30 94 6 vdd
<< end >>
