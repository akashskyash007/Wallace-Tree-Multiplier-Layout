magic
tech scmos
timestamp 1199201872
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 81 70 83 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 24 37
rect 26 35 31 37
rect 19 33 31 35
rect 12 25 14 33
rect 19 25 21 33
rect 29 30 31 33
rect 36 37 42 39
rect 36 35 38 37
rect 40 35 42 37
rect 36 33 42 35
rect 49 37 55 39
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 59 37 71 39
rect 59 35 66 37
rect 68 35 71 37
rect 81 39 83 42
rect 81 37 87 39
rect 81 35 83 37
rect 85 35 87 37
rect 59 33 71 35
rect 36 30 38 33
rect 52 30 54 33
rect 59 30 61 33
rect 69 30 71 33
rect 76 33 87 35
rect 76 30 78 33
rect 69 15 71 20
rect 76 15 78 20
rect 12 10 14 15
rect 19 10 21 15
rect 29 10 31 15
rect 36 10 38 15
rect 52 10 54 15
rect 59 10 61 15
<< ndif >>
rect 24 25 29 30
rect 4 15 12 25
rect 14 15 19 25
rect 21 20 29 25
rect 21 18 24 20
rect 26 18 29 20
rect 21 15 29 18
rect 31 15 36 30
rect 38 19 52 30
rect 38 17 44 19
rect 46 17 52 19
rect 38 15 52 17
rect 54 15 59 30
rect 61 26 69 30
rect 61 24 64 26
rect 66 24 69 26
rect 61 20 69 24
rect 71 20 76 30
rect 78 24 88 30
rect 78 22 83 24
rect 85 22 88 24
rect 78 20 88 22
rect 61 15 66 20
rect 4 11 10 15
rect 4 9 6 11
rect 8 9 10 11
rect 4 7 10 9
<< pdif >>
rect 73 70 79 72
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 42 9 58
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 62 29 70
rect 21 60 24 62
rect 26 60 29 62
rect 21 42 29 60
rect 31 53 39 70
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 61 49 70
rect 41 59 44 61
rect 46 59 49 61
rect 41 54 49 59
rect 41 52 44 54
rect 46 52 49 54
rect 41 42 49 52
rect 51 68 59 70
rect 51 66 54 68
rect 56 66 59 68
rect 51 61 59 66
rect 51 59 54 61
rect 56 59 59 61
rect 51 42 59 59
rect 61 61 69 70
rect 61 59 64 61
rect 66 59 69 61
rect 61 54 69 59
rect 61 52 64 54
rect 66 52 69 54
rect 61 42 69 52
rect 71 68 75 70
rect 77 68 81 70
rect 71 42 81 68
rect 83 63 88 70
rect 83 61 90 63
rect 83 59 86 61
rect 88 59 90 61
rect 83 54 90 59
rect 83 52 86 54
rect 88 52 90 54
rect 83 50 90 52
rect 83 42 88 50
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 70 98 79
rect -2 68 75 70
rect 77 68 98 70
rect 2 53 39 55
rect 2 51 14 53
rect 16 51 34 53
rect 36 51 39 53
rect 2 50 39 51
rect 2 21 6 50
rect 74 46 78 55
rect 10 42 42 46
rect 10 37 14 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 25 14 35
rect 18 37 31 38
rect 18 35 24 37
rect 26 35 31 37
rect 18 34 31 35
rect 36 37 42 42
rect 36 35 38 37
rect 40 35 42 37
rect 36 34 42 35
rect 49 42 86 46
rect 49 37 55 42
rect 49 35 51 37
rect 53 35 55 37
rect 49 34 55 35
rect 64 37 78 38
rect 64 35 66 37
rect 68 35 78 37
rect 64 34 78 35
rect 18 25 22 34
rect 33 26 67 30
rect 33 21 39 26
rect 63 24 64 26
rect 66 24 67 26
rect 63 22 67 24
rect 2 20 39 21
rect 2 18 24 20
rect 26 18 39 20
rect 2 17 39 18
rect 74 17 78 34
rect 82 37 86 42
rect 82 35 83 37
rect 85 35 86 37
rect 82 33 86 35
rect -2 11 98 12
rect -2 9 6 11
rect 8 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 12 15 14 25
rect 19 15 21 25
rect 29 15 31 30
rect 36 15 38 30
rect 52 15 54 30
rect 59 15 61 30
rect 69 20 71 30
rect 76 20 78 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 81 42 83 70
<< polyct1 >>
rect 11 35 13 37
rect 24 35 26 37
rect 38 35 40 37
rect 51 35 53 37
rect 66 35 68 37
rect 83 35 85 37
<< ndifct0 >>
rect 44 17 46 19
rect 83 22 85 24
<< ndifct1 >>
rect 24 18 26 20
rect 64 24 66 26
rect 6 9 8 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 60 6 62
rect 24 60 26 62
rect 44 59 46 61
rect 44 52 46 54
rect 54 66 56 68
rect 54 59 56 61
rect 64 59 66 61
rect 64 52 66 54
rect 86 59 88 61
rect 86 52 88 54
<< pdifct1 >>
rect 14 51 16 53
rect 34 51 36 53
rect 75 68 77 70
<< alu0 >>
rect 52 66 54 68
rect 56 66 58 68
rect 73 67 79 68
rect 2 62 47 63
rect 2 60 4 62
rect 6 60 24 62
rect 26 61 47 62
rect 26 60 44 61
rect 2 59 44 60
rect 46 59 47 61
rect 43 54 47 59
rect 52 61 58 66
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
rect 63 61 89 63
rect 63 59 64 61
rect 66 59 86 61
rect 88 59 89 61
rect 63 54 67 59
rect 43 52 44 54
rect 46 52 64 54
rect 66 52 67 54
rect 43 50 67 52
rect 85 54 89 59
rect 85 52 86 54
rect 88 52 89 54
rect 85 50 89 52
rect 43 19 47 21
rect 43 17 44 19
rect 46 17 47 19
rect 82 24 86 26
rect 82 22 83 24
rect 85 22 86 24
rect 43 12 47 17
rect 82 12 86 22
<< labels >>
rlabel alu0 45 56 45 56 6 n3
rlabel alu0 24 61 24 61 6 n3
rlabel alu0 65 56 65 56 6 n3
rlabel alu0 87 56 87 56 6 n3
rlabel alu1 12 32 12 32 6 b1
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 28 20 28 6 b2
rlabel alu1 20 44 20 44 6 b1
rlabel alu1 28 36 28 36 6 b2
rlabel alu1 28 44 28 44 6 b1
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 36 24 36 24 6 z
rlabel alu1 44 28 44 28 6 z
rlabel alu1 52 28 52 28 6 z
rlabel alu1 36 44 36 44 6 b1
rlabel alu1 52 40 52 40 6 a1
rlabel alu1 36 52 36 52 6 z
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 60 28 60 28 6 z
rlabel alu1 76 24 76 24 6 a2
rlabel alu1 60 44 60 44 6 a1
rlabel alu1 68 36 68 36 6 a2
rlabel alu1 68 44 68 44 6 a1
rlabel alu1 76 48 76 48 6 a1
rlabel polyct1 84 36 84 36 6 a1
<< end >>
