magic
tech scmos
timestamp 1199202924
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 37 28 39
rect 33 39 35 42
rect 43 39 45 42
rect 33 37 45 39
rect 50 39 52 42
rect 60 39 62 42
rect 50 37 62 39
rect 22 35 24 37
rect 26 35 28 37
rect 22 33 28 35
rect 35 35 41 37
rect 35 33 37 35
rect 39 33 41 35
rect 50 35 52 37
rect 54 35 56 37
rect 50 33 56 35
rect 9 31 18 33
rect 12 29 14 31
rect 16 29 18 31
rect 12 27 18 29
rect 13 24 15 27
rect 23 24 25 33
rect 35 31 41 33
rect 45 31 56 33
rect 67 31 69 42
rect 35 28 37 31
rect 45 28 47 31
rect 63 29 69 31
rect 63 27 65 29
rect 67 27 69 29
rect 63 25 69 27
rect 13 6 15 11
rect 23 6 25 11
rect 35 6 37 11
rect 45 6 47 11
<< ndif >>
rect 27 24 35 28
rect 4 11 13 24
rect 15 21 23 24
rect 15 19 18 21
rect 20 19 23 21
rect 15 11 23 19
rect 25 11 35 24
rect 37 21 45 28
rect 37 19 40 21
rect 42 19 45 21
rect 37 11 45 19
rect 47 22 55 28
rect 47 20 50 22
rect 52 20 55 22
rect 47 15 55 20
rect 47 13 50 15
rect 52 13 55 15
rect 47 11 55 13
rect 4 9 7 11
rect 9 9 11 11
rect 4 7 11 9
rect 27 9 29 11
rect 31 9 33 11
rect 27 7 33 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 42 16 70
rect 18 53 26 70
rect 18 51 21 53
rect 23 51 26 53
rect 18 46 26 51
rect 18 44 21 46
rect 23 44 26 46
rect 18 42 26 44
rect 28 42 33 70
rect 35 68 43 70
rect 35 66 38 68
rect 40 66 43 68
rect 35 61 43 66
rect 35 59 38 61
rect 40 59 43 61
rect 35 42 43 59
rect 45 42 50 70
rect 52 53 60 70
rect 52 51 55 53
rect 57 51 60 53
rect 52 46 60 51
rect 52 44 55 46
rect 57 44 60 46
rect 52 42 60 44
rect 62 42 67 70
rect 69 68 77 70
rect 69 66 72 68
rect 74 66 77 68
rect 69 61 77 66
rect 69 59 72 61
rect 74 59 77 61
rect 69 42 77 59
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 19 53 59 54
rect 19 51 21 53
rect 23 51 55 53
rect 57 51 59 53
rect 19 50 59 51
rect 19 47 24 50
rect 2 46 24 47
rect 54 46 59 50
rect 2 44 21 46
rect 23 44 24 46
rect 2 42 24 44
rect 28 42 50 46
rect 54 44 55 46
rect 57 44 63 46
rect 54 42 63 44
rect 2 22 6 42
rect 28 38 32 42
rect 22 37 32 38
rect 46 38 50 42
rect 46 37 63 38
rect 22 35 24 37
rect 26 35 32 37
rect 22 34 32 35
rect 36 35 40 37
rect 36 33 37 35
rect 39 33 40 35
rect 46 35 52 37
rect 54 35 63 37
rect 46 34 63 35
rect 13 31 17 33
rect 13 29 14 31
rect 16 30 17 31
rect 36 30 40 33
rect 16 29 70 30
rect 13 27 65 29
rect 67 27 70 29
rect 13 26 70 27
rect 2 21 44 22
rect 2 19 18 21
rect 20 19 40 21
rect 42 19 44 21
rect 2 18 44 19
rect 66 17 70 26
rect -2 11 82 12
rect -2 9 7 11
rect 9 9 29 11
rect 31 9 82 11
rect -2 1 82 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 13 11 15 24
rect 23 11 25 24
rect 35 11 37 28
rect 45 11 47 28
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
<< polyct1 >>
rect 24 35 26 37
rect 37 33 39 35
rect 52 35 54 37
rect 14 29 16 31
rect 65 27 67 29
<< ndifct0 >>
rect 50 20 52 22
rect 50 13 52 15
<< ndifct1 >>
rect 18 19 20 21
rect 40 19 42 21
rect 7 9 9 11
rect 29 9 31 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 38 66 40 68
rect 38 59 40 61
rect 72 66 74 68
rect 72 59 74 61
<< pdifct1 >>
rect 21 51 23 53
rect 21 44 23 46
rect 55 51 57 53
rect 55 44 57 46
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 36 66 38 68
rect 40 66 42 68
rect 36 61 42 66
rect 36 59 38 61
rect 40 59 42 61
rect 36 58 42 59
rect 70 66 72 68
rect 74 66 76 68
rect 70 61 76 66
rect 70 59 72 61
rect 74 59 76 61
rect 70 58 76 59
rect 48 22 54 23
rect 48 20 50 22
rect 52 20 54 22
rect 48 15 54 20
rect 48 13 50 15
rect 52 13 54 15
rect 48 12 54 13
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 28 36 28 36 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 28 44 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 52 28 52 28 6 a
rlabel alu1 60 28 60 28 6 a
rlabel alu1 52 36 52 36 6 b
rlabel alu1 60 36 60 36 6 b
rlabel alu1 60 44 60 44 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 68 20 68 20 6 a
<< end >>
