magic
tech scmos
timestamp 1199201799
<< ab >>
rect 0 0 168 72
<< nwell >>
rect -5 32 173 77
<< pwell >>
rect -5 -5 173 32
<< poly >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 50 66 52 70
rect 60 66 62 70
rect 67 66 69 70
rect 77 66 79 70
rect 107 66 109 70
rect 117 66 119 70
rect 127 66 129 70
rect 137 66 139 70
rect 147 66 149 70
rect 157 66 159 70
rect 87 52 89 57
rect 97 52 99 57
rect 9 25 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 16 33 28 35
rect 16 31 19 33
rect 21 31 23 33
rect 33 31 35 38
rect 43 31 45 38
rect 50 35 52 38
rect 60 35 62 38
rect 50 33 62 35
rect 50 31 52 33
rect 54 31 56 33
rect 16 29 23 31
rect 32 29 46 31
rect 50 29 56 31
rect 32 27 34 29
rect 28 25 34 27
rect 44 26 46 29
rect 54 26 56 29
rect 67 28 69 38
rect 77 35 79 38
rect 87 35 89 38
rect 97 35 99 38
rect 107 35 109 38
rect 117 35 119 38
rect 77 33 119 35
rect 127 35 129 38
rect 137 35 139 38
rect 147 35 149 38
rect 157 35 159 38
rect 127 33 159 35
rect 81 31 83 33
rect 85 31 87 33
rect 81 29 87 31
rect 113 31 115 33
rect 117 31 119 33
rect 113 29 119 31
rect 130 31 132 33
rect 134 31 136 33
rect 130 29 136 31
rect 66 26 72 28
rect 9 23 30 25
rect 32 23 34 25
rect 28 21 34 23
rect 66 24 68 26
rect 70 24 72 26
rect 91 27 109 29
rect 113 27 126 29
rect 91 25 97 27
rect 66 22 72 24
rect 44 2 46 6
rect 54 2 56 6
rect 91 23 93 25
rect 95 23 97 25
rect 107 24 109 27
rect 114 24 116 27
rect 124 24 126 27
rect 131 24 133 29
rect 91 21 97 23
rect 107 2 109 7
rect 114 2 116 7
rect 124 2 126 7
rect 131 2 133 7
<< ndif >>
rect 36 7 44 26
rect 36 5 38 7
rect 40 6 44 7
rect 46 17 54 26
rect 46 15 49 17
rect 51 15 54 17
rect 46 6 54 15
rect 56 7 64 26
rect 56 6 60 7
rect 40 5 42 6
rect 36 3 42 5
rect 58 5 60 6
rect 62 5 64 7
rect 58 3 64 5
rect 99 7 107 24
rect 109 7 114 24
rect 116 17 124 24
rect 116 15 119 17
rect 121 15 124 17
rect 116 7 124 15
rect 126 7 131 24
rect 133 18 146 24
rect 133 16 141 18
rect 143 16 146 18
rect 133 11 146 16
rect 133 9 141 11
rect 143 9 146 11
rect 133 7 146 9
rect 99 5 101 7
rect 103 5 105 7
rect 99 3 105 5
<< pdif >>
rect 4 60 9 66
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 54 9 56
rect 4 38 9 54
rect 11 38 16 66
rect 18 49 26 66
rect 18 47 21 49
rect 23 47 26 49
rect 18 38 26 47
rect 28 38 33 66
rect 35 58 43 66
rect 35 56 38 58
rect 40 56 43 58
rect 35 38 43 56
rect 45 38 50 66
rect 52 49 60 66
rect 52 47 55 49
rect 57 47 60 49
rect 52 42 60 47
rect 52 40 55 42
rect 57 40 60 42
rect 52 38 60 40
rect 62 38 67 66
rect 69 57 77 66
rect 69 55 72 57
rect 74 55 77 57
rect 69 50 77 55
rect 69 48 72 50
rect 74 48 77 50
rect 69 43 77 48
rect 69 41 72 43
rect 74 41 77 43
rect 69 38 77 41
rect 79 64 86 66
rect 79 62 82 64
rect 84 62 86 64
rect 79 60 86 62
rect 79 52 85 60
rect 100 64 107 66
rect 100 62 102 64
rect 104 62 107 64
rect 100 60 107 62
rect 101 52 107 60
rect 79 50 87 52
rect 79 48 82 50
rect 84 48 87 50
rect 79 38 87 48
rect 89 49 97 52
rect 89 47 92 49
rect 94 47 97 49
rect 89 42 97 47
rect 89 40 92 42
rect 94 40 97 42
rect 89 38 97 40
rect 99 50 107 52
rect 99 48 102 50
rect 104 48 107 50
rect 99 38 107 48
rect 109 57 117 66
rect 109 55 112 57
rect 114 55 117 57
rect 109 50 117 55
rect 109 48 112 50
rect 114 48 117 50
rect 109 43 117 48
rect 109 41 112 43
rect 114 41 117 43
rect 109 38 117 41
rect 119 64 127 66
rect 119 62 122 64
rect 124 62 127 64
rect 119 57 127 62
rect 119 55 122 57
rect 124 55 127 57
rect 119 38 127 55
rect 129 56 137 66
rect 129 54 132 56
rect 134 54 137 56
rect 129 49 137 54
rect 129 47 132 49
rect 134 47 137 49
rect 129 38 137 47
rect 139 64 147 66
rect 139 62 142 64
rect 144 62 147 64
rect 139 57 147 62
rect 139 55 142 57
rect 144 55 147 57
rect 139 38 147 55
rect 149 57 157 66
rect 149 55 152 57
rect 154 55 157 57
rect 149 50 157 55
rect 149 48 152 50
rect 154 48 157 50
rect 149 43 157 48
rect 149 41 152 43
rect 154 41 157 43
rect 149 38 157 41
rect 159 64 166 66
rect 159 62 162 64
rect 164 62 166 64
rect 159 57 166 62
rect 159 55 162 57
rect 164 55 166 57
rect 159 38 166 55
<< alu1 >>
rect -2 67 170 72
rect -2 65 92 67
rect 94 65 170 67
rect -2 64 170 65
rect 2 49 59 50
rect 2 47 21 49
rect 23 47 55 49
rect 57 47 59 49
rect 2 46 59 47
rect 2 18 6 46
rect 53 42 59 46
rect 17 34 23 42
rect 53 40 55 42
rect 57 40 59 42
rect 53 39 59 40
rect 17 33 56 34
rect 17 31 19 33
rect 21 31 52 33
rect 54 31 56 33
rect 17 30 56 31
rect 17 22 23 30
rect 66 26 71 35
rect 28 25 68 26
rect 28 23 30 25
rect 32 24 68 25
rect 70 24 71 26
rect 32 23 71 24
rect 28 22 71 23
rect 81 33 119 34
rect 81 31 83 33
rect 85 31 115 33
rect 117 31 119 33
rect 81 30 119 31
rect 130 33 134 43
rect 130 31 132 33
rect 81 22 87 30
rect 130 26 134 31
rect 91 25 134 26
rect 91 23 93 25
rect 95 23 134 25
rect 91 22 134 23
rect 2 17 123 18
rect 2 15 49 17
rect 51 15 119 17
rect 121 15 123 17
rect 2 14 123 15
rect 130 13 134 22
rect -2 7 170 8
rect -2 5 5 7
rect 7 5 13 7
rect 15 5 38 7
rect 40 5 60 7
rect 62 5 80 7
rect 82 5 101 7
rect 103 5 153 7
rect 155 5 161 7
rect 163 5 170 7
rect -2 0 170 5
<< ptie >>
rect 3 7 17 20
rect 3 5 5 7
rect 7 5 13 7
rect 15 5 17 7
rect 3 3 17 5
rect 75 7 87 24
rect 75 5 80 7
rect 82 5 87 7
rect 75 3 87 5
rect 151 7 165 24
rect 151 5 153 7
rect 155 5 161 7
rect 163 5 165 7
rect 151 3 165 5
<< ntie >>
rect 90 67 96 69
rect 90 65 92 67
rect 94 65 96 67
rect 90 59 96 65
<< nmos >>
rect 44 6 46 26
rect 54 6 56 26
rect 107 7 109 24
rect 114 7 116 24
rect 124 7 126 24
rect 131 7 133 24
<< pmos >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 38 45 66
rect 50 38 52 66
rect 60 38 62 66
rect 67 38 69 66
rect 77 38 79 66
rect 87 38 89 52
rect 97 38 99 52
rect 107 38 109 66
rect 117 38 119 66
rect 127 38 129 66
rect 137 38 139 66
rect 147 38 149 66
rect 157 38 159 66
<< polyct1 >>
rect 19 31 21 33
rect 52 31 54 33
rect 83 31 85 33
rect 115 31 117 33
rect 132 31 134 33
rect 30 23 32 25
rect 68 24 70 26
rect 93 23 95 25
<< ndifct0 >>
rect 141 16 143 18
rect 141 9 143 11
<< ndifct1 >>
rect 38 5 40 7
rect 49 15 51 17
rect 60 5 62 7
rect 119 15 121 17
rect 101 5 103 7
<< ntiect1 >>
rect 92 65 94 67
<< ptiect1 >>
rect 5 5 7 7
rect 13 5 15 7
rect 80 5 82 7
rect 153 5 155 7
rect 161 5 163 7
<< pdifct0 >>
rect 4 56 6 58
rect 38 56 40 58
rect 72 55 74 57
rect 72 48 74 50
rect 72 41 74 43
rect 82 62 84 64
rect 102 62 104 64
rect 82 48 84 50
rect 92 47 94 49
rect 92 40 94 42
rect 102 48 104 50
rect 112 55 114 57
rect 112 48 114 50
rect 112 41 114 43
rect 122 62 124 64
rect 122 55 124 57
rect 132 54 134 56
rect 132 47 134 49
rect 142 62 144 64
rect 142 55 144 57
rect 152 55 154 57
rect 152 48 154 50
rect 152 41 154 43
rect 162 62 164 64
rect 162 55 164 57
<< pdifct1 >>
rect 21 47 23 49
rect 55 47 57 49
rect 55 40 57 42
<< alu0 >>
rect 80 62 82 64
rect 84 62 86 64
rect 2 58 75 59
rect 2 56 4 58
rect 6 56 38 58
rect 40 57 75 58
rect 40 56 72 57
rect 2 55 72 56
rect 74 55 75 57
rect 71 50 75 55
rect 71 48 72 50
rect 74 48 75 50
rect 71 43 75 48
rect 80 50 86 62
rect 100 62 102 64
rect 104 62 106 64
rect 80 48 82 50
rect 84 48 86 50
rect 80 47 86 48
rect 91 49 95 51
rect 91 47 92 49
rect 94 47 95 49
rect 100 50 106 62
rect 120 62 122 64
rect 124 62 126 64
rect 100 48 102 50
rect 104 48 106 50
rect 100 47 106 48
rect 111 57 115 59
rect 111 55 112 57
rect 114 55 115 57
rect 111 50 115 55
rect 120 57 126 62
rect 140 62 142 64
rect 144 62 146 64
rect 120 55 122 57
rect 124 55 126 57
rect 120 54 126 55
rect 131 56 135 58
rect 131 54 132 56
rect 134 54 135 56
rect 140 57 146 62
rect 161 62 162 64
rect 164 62 165 64
rect 140 55 142 57
rect 144 55 146 57
rect 140 54 146 55
rect 151 57 155 59
rect 151 55 152 57
rect 154 55 155 57
rect 131 50 135 54
rect 151 50 155 55
rect 161 57 165 62
rect 161 55 162 57
rect 164 55 165 57
rect 161 53 165 55
rect 111 48 112 50
rect 114 49 152 50
rect 114 48 132 49
rect 111 47 132 48
rect 134 48 152 49
rect 154 48 155 50
rect 134 47 155 48
rect 91 43 95 47
rect 111 46 155 47
rect 111 43 115 46
rect 151 43 155 46
rect 71 41 72 43
rect 74 42 112 43
rect 74 41 92 42
rect 71 40 92 41
rect 94 41 112 42
rect 114 41 115 43
rect 94 40 115 41
rect 71 39 115 40
rect 151 41 152 43
rect 154 41 155 43
rect 151 39 155 41
rect 134 29 135 35
rect 139 18 145 19
rect 139 16 141 18
rect 143 16 145 18
rect 139 11 145 16
rect 139 9 141 11
rect 143 9 145 11
rect 139 8 145 9
<< labels >>
rlabel pdifct0 73 49 73 49 6 n1
rlabel alu0 38 57 38 57 6 n1
rlabel alu0 93 45 93 45 6 n1
rlabel pdifct0 133 48 133 48 6 n1
rlabel pdifct0 153 49 153 49 6 n1
rlabel alu0 133 52 133 52 6 n1
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 28 32 28 32 6 c
rlabel polyct1 20 32 20 32 6 c
rlabel alu1 28 48 28 48 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 60 16 60 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 60 24 60 24 6 b
rlabel alu1 52 24 52 24 6 b
rlabel alu1 44 24 44 24 6 b
rlabel alu1 36 24 36 24 6 b
rlabel alu1 52 32 52 32 6 c
rlabel alu1 44 32 44 32 6 c
rlabel alu1 36 32 36 32 6 c
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 84 4 84 4 6 vss
rlabel alu1 92 16 92 16 6 z
rlabel alu1 84 16 84 16 6 z
rlabel alu1 76 16 76 16 6 z
rlabel alu1 68 16 68 16 6 z
rlabel alu1 92 32 92 32 6 a2
rlabel alu1 84 28 84 28 6 a2
rlabel alu1 68 28 68 28 6 b
rlabel alu1 84 68 84 68 6 vdd
rlabel alu1 116 16 116 16 6 z
rlabel alu1 108 16 108 16 6 z
rlabel alu1 100 16 100 16 6 z
rlabel alu1 100 24 100 24 6 a1
rlabel alu1 124 24 124 24 6 a1
rlabel alu1 116 24 116 24 6 a1
rlabel alu1 108 24 108 24 6 a1
rlabel polyct1 116 32 116 32 6 a2
rlabel alu1 108 32 108 32 6 a2
rlabel alu1 132 28 132 28 6 a1
rlabel alu1 100 32 100 32 6 a2
<< end >>
