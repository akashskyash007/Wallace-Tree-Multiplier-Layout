magic
tech scmos
timestamp 1199201841
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 29 66 31 71
rect 9 58 11 63
rect 19 58 21 63
rect 29 47 31 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 9 39 11 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 35 21 42
rect 29 41 35 43
rect 19 33 25 35
rect 12 25 14 33
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 22 26 24 29
rect 29 26 31 41
rect 12 15 14 19
rect 22 15 24 19
rect 29 15 31 19
<< ndif >>
rect 17 25 22 26
rect 3 19 12 25
rect 14 23 22 25
rect 14 21 17 23
rect 19 21 22 23
rect 14 19 22 21
rect 24 19 29 26
rect 31 19 38 26
rect 3 11 10 19
rect 33 13 38 19
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
rect 32 11 38 13
rect 32 9 34 11
rect 36 9 38 11
rect 32 7 38 9
<< pdif >>
rect 21 71 27 73
rect 21 69 23 71
rect 25 69 27 71
rect 21 66 27 69
rect 21 65 29 66
rect 23 58 29 65
rect 4 55 9 58
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 56 19 58
rect 11 54 14 56
rect 16 54 19 56
rect 11 42 19 54
rect 21 50 29 58
rect 31 63 36 66
rect 31 61 38 63
rect 31 59 34 61
rect 36 59 38 61
rect 31 54 38 59
rect 31 52 34 54
rect 36 52 38 54
rect 31 50 38 52
rect 21 42 27 50
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 71 42 79
rect -2 69 23 71
rect 25 69 42 71
rect -2 68 42 69
rect 2 53 6 55
rect 2 51 4 53
rect 2 46 6 51
rect 2 44 4 46
rect 2 23 6 44
rect 26 47 30 55
rect 10 41 22 47
rect 26 45 38 47
rect 26 43 31 45
rect 33 43 38 45
rect 26 41 38 43
rect 10 37 14 41
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 19 33 25 34
rect 19 31 21 33
rect 23 31 30 33
rect 19 29 30 31
rect 26 23 30 29
rect 2 21 17 23
rect 19 21 22 23
rect 2 17 22 21
rect 26 17 38 23
rect -2 11 42 12
rect -2 9 6 11
rect 8 9 34 11
rect 36 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 12 19 14 25
rect 22 19 24 26
rect 29 19 31 26
<< pmos >>
rect 9 42 11 58
rect 19 42 21 58
rect 29 50 31 66
<< polyct1 >>
rect 31 43 33 45
rect 11 35 13 37
rect 21 31 23 33
<< ndifct1 >>
rect 17 21 19 23
rect 6 9 8 11
rect 34 9 36 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 54 16 56
rect 34 59 36 61
rect 34 52 36 54
<< pdifct1 >>
rect 23 69 25 71
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 13 61 37 63
rect 13 59 34 61
rect 36 59 37 61
rect 13 56 17 59
rect 6 42 7 55
rect 13 54 14 56
rect 16 54 17 56
rect 13 52 17 54
rect 33 54 37 59
rect 33 52 34 54
rect 36 52 37 54
rect 33 50 37 52
rect 16 23 20 25
<< labels >>
rlabel alu0 15 57 15 57 6 n1
rlabel alu0 35 56 35 56 6 n1
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 24 28 24 6 a2
rlabel alu1 20 44 20 44 6 b
rlabel alu1 28 48 28 48 6 a1
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 20 36 20 6 a2
rlabel alu1 36 44 36 44 6 a1
<< end >>
