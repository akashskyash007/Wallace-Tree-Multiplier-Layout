magic
tech scmos
timestamp 1554086911
<< ab >>
rect 11 9 91 297
rect 93 9 311 297
rect 319 9 359 297
rect 361 9 579 297
rect 587 9 627 297
rect 628 9 846 297
<< nwell >>
rect 6 185 851 265
rect 6 41 851 121
<< pwell >>
rect 6 265 851 302
rect 6 121 851 185
rect 6 4 851 41
<< poly >>
rect 20 284 22 289
rect 27 284 29 289
rect 40 282 42 286
rect 60 284 62 289
rect 67 284 69 289
rect 102 291 104 295
rect 80 282 82 286
rect 112 288 114 293
rect 152 291 154 295
rect 159 291 161 295
rect 170 291 172 295
rect 191 291 193 295
rect 122 285 124 290
rect 132 285 134 290
rect 102 275 104 278
rect 102 273 108 275
rect 20 260 22 273
rect 27 268 29 273
rect 40 268 42 273
rect 26 266 32 268
rect 26 264 28 266
rect 30 264 32 266
rect 26 262 32 264
rect 36 266 42 268
rect 36 264 38 266
rect 40 264 42 266
rect 36 262 42 264
rect 16 258 22 260
rect 16 256 18 258
rect 20 256 22 258
rect 16 254 22 256
rect 20 251 22 254
rect 30 251 32 262
rect 40 258 42 262
rect 60 260 62 273
rect 67 268 69 273
rect 80 268 82 273
rect 66 266 72 268
rect 66 264 68 266
rect 70 264 72 266
rect 66 262 72 264
rect 76 266 82 268
rect 76 264 78 266
rect 80 264 82 266
rect 76 262 82 264
rect 56 258 62 260
rect 56 256 58 258
rect 60 256 62 258
rect 56 254 62 256
rect 60 251 62 254
rect 70 251 72 262
rect 80 258 82 262
rect 102 271 104 273
rect 106 271 108 273
rect 102 269 108 271
rect 20 233 22 238
rect 30 233 32 238
rect 40 236 42 240
rect 102 256 104 269
rect 112 265 114 278
rect 201 288 203 293
rect 241 291 243 295
rect 248 291 250 295
rect 259 291 261 295
rect 211 285 213 290
rect 221 285 223 290
rect 108 263 114 265
rect 108 261 110 263
rect 112 261 114 263
rect 122 268 124 271
rect 132 268 134 271
rect 152 268 154 271
rect 159 268 161 271
rect 170 268 172 277
rect 191 275 193 278
rect 191 273 197 275
rect 191 271 193 273
rect 195 271 197 273
rect 191 269 197 271
rect 122 266 128 268
rect 122 264 124 266
rect 126 264 128 266
rect 122 262 128 264
rect 132 266 154 268
rect 132 264 143 266
rect 145 264 150 266
rect 152 264 154 266
rect 132 262 154 264
rect 158 266 164 268
rect 158 264 160 266
rect 162 264 164 266
rect 158 262 164 264
rect 168 266 174 268
rect 168 264 170 266
rect 172 264 174 266
rect 168 262 174 264
rect 108 259 117 261
rect 125 259 127 262
rect 132 259 134 262
rect 150 259 152 262
rect 160 259 162 262
rect 170 259 172 262
rect 115 256 117 259
rect 60 233 62 238
rect 70 233 72 238
rect 80 236 82 240
rect 115 238 117 243
rect 102 227 104 231
rect 125 229 127 234
rect 132 229 134 234
rect 191 256 193 269
rect 201 265 203 278
rect 280 285 282 290
rect 197 263 203 265
rect 197 261 199 263
rect 201 261 203 263
rect 211 268 213 271
rect 221 268 223 271
rect 241 268 243 271
rect 248 268 250 271
rect 259 268 261 277
rect 290 284 292 289
rect 300 282 302 286
rect 328 284 330 289
rect 335 284 337 289
rect 370 291 372 295
rect 280 268 282 271
rect 290 268 292 276
rect 300 268 302 274
rect 348 282 350 286
rect 380 288 382 293
rect 420 291 422 295
rect 427 291 429 295
rect 438 291 440 295
rect 459 291 461 295
rect 390 285 392 290
rect 400 285 402 290
rect 370 275 372 278
rect 370 273 376 275
rect 211 266 217 268
rect 211 264 213 266
rect 215 264 217 266
rect 211 262 217 264
rect 221 266 243 268
rect 221 264 232 266
rect 234 264 239 266
rect 241 264 243 266
rect 221 262 243 264
rect 247 266 253 268
rect 247 264 249 266
rect 251 264 253 266
rect 247 262 253 264
rect 257 266 263 268
rect 257 264 259 266
rect 261 264 263 266
rect 257 262 263 264
rect 280 266 286 268
rect 280 264 282 266
rect 284 264 286 266
rect 280 262 286 264
rect 290 266 296 268
rect 290 264 292 266
rect 294 264 296 266
rect 290 262 296 264
rect 300 266 309 268
rect 300 264 305 266
rect 307 264 309 266
rect 300 262 309 264
rect 197 259 206 261
rect 214 259 216 262
rect 221 259 223 262
rect 239 259 241 262
rect 249 259 251 262
rect 259 259 261 262
rect 280 259 282 262
rect 293 259 295 262
rect 300 259 302 262
rect 328 260 330 273
rect 335 268 337 273
rect 348 268 350 273
rect 334 266 340 268
rect 334 264 336 266
rect 338 264 340 266
rect 334 262 340 264
rect 344 266 350 268
rect 344 264 346 266
rect 348 264 350 266
rect 344 262 350 264
rect 204 256 206 259
rect 204 238 206 243
rect 150 227 152 231
rect 160 227 162 231
rect 170 227 172 231
rect 191 227 193 231
rect 214 229 216 234
rect 221 229 223 234
rect 239 227 241 231
rect 249 227 251 231
rect 259 227 261 231
rect 280 227 282 231
rect 324 258 330 260
rect 324 256 326 258
rect 328 256 330 258
rect 324 254 330 256
rect 328 251 330 254
rect 338 251 340 262
rect 348 258 350 262
rect 370 271 372 273
rect 374 271 376 273
rect 370 269 376 271
rect 370 256 372 269
rect 380 265 382 278
rect 469 288 471 293
rect 509 291 511 295
rect 516 291 518 295
rect 527 291 529 295
rect 479 285 481 290
rect 489 285 491 290
rect 376 263 382 265
rect 376 261 378 263
rect 380 261 382 263
rect 390 268 392 271
rect 400 268 402 271
rect 420 268 422 271
rect 427 268 429 271
rect 438 268 440 277
rect 459 275 461 278
rect 459 273 465 275
rect 459 271 461 273
rect 463 271 465 273
rect 459 269 465 271
rect 390 266 396 268
rect 390 264 392 266
rect 394 264 396 266
rect 390 262 396 264
rect 400 266 422 268
rect 400 264 411 266
rect 413 264 418 266
rect 420 264 422 266
rect 400 262 422 264
rect 426 266 432 268
rect 426 264 428 266
rect 430 264 432 266
rect 426 262 432 264
rect 436 266 442 268
rect 436 264 438 266
rect 440 264 442 266
rect 436 262 442 264
rect 376 259 385 261
rect 393 259 395 262
rect 400 259 402 262
rect 418 259 420 262
rect 428 259 430 262
rect 438 259 440 262
rect 383 256 385 259
rect 328 233 330 238
rect 338 233 340 238
rect 348 236 350 240
rect 293 227 295 231
rect 300 227 302 231
rect 383 238 385 243
rect 370 227 372 231
rect 393 229 395 234
rect 400 229 402 234
rect 459 256 461 269
rect 469 265 471 278
rect 548 285 550 290
rect 465 263 471 265
rect 465 261 467 263
rect 469 261 471 263
rect 479 268 481 271
rect 489 268 491 271
rect 509 268 511 271
rect 516 268 518 271
rect 527 268 529 277
rect 558 284 560 289
rect 568 282 570 286
rect 596 284 598 289
rect 603 284 605 289
rect 637 291 639 295
rect 548 268 550 271
rect 558 268 560 276
rect 568 268 570 274
rect 616 282 618 286
rect 647 288 649 293
rect 687 291 689 295
rect 694 291 696 295
rect 705 291 707 295
rect 726 291 728 295
rect 657 285 659 290
rect 667 285 669 290
rect 637 275 639 278
rect 637 273 643 275
rect 479 266 485 268
rect 479 264 481 266
rect 483 264 485 266
rect 479 262 485 264
rect 489 266 511 268
rect 489 264 500 266
rect 502 264 507 266
rect 509 264 511 266
rect 489 262 511 264
rect 515 266 521 268
rect 515 264 517 266
rect 519 264 521 266
rect 515 262 521 264
rect 525 266 531 268
rect 525 264 527 266
rect 529 264 531 266
rect 525 262 531 264
rect 548 266 554 268
rect 548 264 550 266
rect 552 264 554 266
rect 548 262 554 264
rect 558 266 564 268
rect 558 264 560 266
rect 562 264 564 266
rect 558 262 564 264
rect 568 266 577 268
rect 568 264 573 266
rect 575 264 577 266
rect 568 262 577 264
rect 465 259 474 261
rect 482 259 484 262
rect 489 259 491 262
rect 507 259 509 262
rect 517 259 519 262
rect 527 259 529 262
rect 548 259 550 262
rect 561 259 563 262
rect 568 259 570 262
rect 596 260 598 273
rect 603 268 605 273
rect 616 268 618 273
rect 602 266 608 268
rect 602 264 604 266
rect 606 264 608 266
rect 602 262 608 264
rect 612 266 618 268
rect 612 264 614 266
rect 616 264 618 266
rect 612 262 618 264
rect 472 256 474 259
rect 472 238 474 243
rect 418 227 420 231
rect 428 227 430 231
rect 438 227 440 231
rect 459 227 461 231
rect 482 229 484 234
rect 489 229 491 234
rect 507 227 509 231
rect 517 227 519 231
rect 527 227 529 231
rect 548 227 550 231
rect 592 258 598 260
rect 592 256 594 258
rect 596 256 598 258
rect 592 254 598 256
rect 596 251 598 254
rect 606 251 608 262
rect 616 258 618 262
rect 637 271 639 273
rect 641 271 643 273
rect 637 269 643 271
rect 637 256 639 269
rect 647 265 649 278
rect 736 288 738 293
rect 776 291 778 295
rect 783 291 785 295
rect 794 291 796 295
rect 746 285 748 290
rect 756 285 758 290
rect 643 263 649 265
rect 643 261 645 263
rect 647 261 649 263
rect 657 268 659 271
rect 667 268 669 271
rect 687 268 689 271
rect 694 268 696 271
rect 705 268 707 277
rect 726 275 728 278
rect 726 273 732 275
rect 726 271 728 273
rect 730 271 732 273
rect 726 269 732 271
rect 657 266 663 268
rect 657 264 659 266
rect 661 264 663 266
rect 657 262 663 264
rect 667 266 689 268
rect 667 264 678 266
rect 680 264 685 266
rect 687 264 689 266
rect 667 262 689 264
rect 693 266 699 268
rect 693 264 695 266
rect 697 264 699 266
rect 693 262 699 264
rect 703 266 709 268
rect 703 264 705 266
rect 707 264 709 266
rect 703 262 709 264
rect 643 259 652 261
rect 660 259 662 262
rect 667 259 669 262
rect 685 259 687 262
rect 695 259 697 262
rect 705 259 707 262
rect 650 256 652 259
rect 596 233 598 238
rect 606 233 608 238
rect 616 236 618 240
rect 561 227 563 231
rect 568 227 570 231
rect 650 238 652 243
rect 637 227 639 231
rect 660 229 662 234
rect 667 229 669 234
rect 726 256 728 269
rect 736 265 738 278
rect 815 285 817 290
rect 732 263 738 265
rect 732 261 734 263
rect 736 261 738 263
rect 746 268 748 271
rect 756 268 758 271
rect 776 268 778 271
rect 783 268 785 271
rect 794 268 796 277
rect 825 284 827 289
rect 835 282 837 286
rect 815 268 817 271
rect 825 268 827 276
rect 835 268 837 274
rect 746 266 752 268
rect 746 264 748 266
rect 750 264 752 266
rect 746 262 752 264
rect 756 266 778 268
rect 756 264 767 266
rect 769 264 774 266
rect 776 264 778 266
rect 756 262 778 264
rect 782 266 788 268
rect 782 264 784 266
rect 786 264 788 266
rect 782 262 788 264
rect 792 266 798 268
rect 792 264 794 266
rect 796 264 798 266
rect 792 262 798 264
rect 815 266 821 268
rect 815 264 817 266
rect 819 264 821 266
rect 815 262 821 264
rect 825 266 831 268
rect 825 264 827 266
rect 829 264 831 266
rect 825 262 831 264
rect 835 266 844 268
rect 835 264 840 266
rect 842 264 844 266
rect 835 262 844 264
rect 732 259 741 261
rect 749 259 751 262
rect 756 259 758 262
rect 774 259 776 262
rect 784 259 786 262
rect 794 259 796 262
rect 815 259 817 262
rect 828 259 830 262
rect 835 259 837 262
rect 739 256 741 259
rect 739 238 741 243
rect 685 227 687 231
rect 695 227 697 231
rect 705 227 707 231
rect 726 227 728 231
rect 749 229 751 234
rect 756 229 758 234
rect 774 227 776 231
rect 784 227 786 231
rect 794 227 796 231
rect 815 227 817 231
rect 828 227 830 231
rect 835 227 837 231
rect 20 212 22 217
rect 30 212 32 217
rect 102 219 104 223
rect 40 210 42 214
rect 60 212 62 217
rect 70 212 72 217
rect 20 196 22 199
rect 16 194 22 196
rect 16 192 18 194
rect 20 192 22 194
rect 16 190 22 192
rect 20 177 22 190
rect 30 188 32 199
rect 80 210 82 214
rect 60 196 62 199
rect 56 194 62 196
rect 56 192 58 194
rect 60 192 62 194
rect 40 188 42 192
rect 56 190 62 192
rect 26 186 32 188
rect 26 184 28 186
rect 30 184 32 186
rect 26 182 32 184
rect 36 186 42 188
rect 36 184 38 186
rect 40 184 42 186
rect 36 182 42 184
rect 27 177 29 182
rect 40 177 42 182
rect 60 177 62 190
rect 70 188 72 199
rect 125 216 127 221
rect 132 216 134 221
rect 150 219 152 223
rect 160 219 162 223
rect 170 219 172 223
rect 191 219 193 223
rect 115 207 117 212
rect 80 188 82 192
rect 66 186 72 188
rect 66 184 68 186
rect 70 184 72 186
rect 66 182 72 184
rect 76 186 82 188
rect 76 184 78 186
rect 80 184 82 186
rect 76 182 82 184
rect 67 177 69 182
rect 80 177 82 182
rect 102 181 104 194
rect 115 191 117 194
rect 214 216 216 221
rect 221 216 223 221
rect 239 219 241 223
rect 249 219 251 223
rect 259 219 261 223
rect 280 219 282 223
rect 204 207 206 212
rect 108 189 117 191
rect 108 187 110 189
rect 112 187 114 189
rect 125 188 127 191
rect 132 188 134 191
rect 150 188 152 191
rect 160 188 162 191
rect 170 188 172 191
rect 108 185 114 187
rect 102 179 108 181
rect 102 177 104 179
rect 106 177 108 179
rect 20 161 22 166
rect 27 161 29 166
rect 40 164 42 168
rect 102 175 108 177
rect 102 172 104 175
rect 112 172 114 185
rect 122 186 128 188
rect 122 184 124 186
rect 126 184 128 186
rect 122 182 128 184
rect 132 186 154 188
rect 132 184 143 186
rect 145 184 150 186
rect 152 184 154 186
rect 132 182 154 184
rect 158 186 164 188
rect 158 184 160 186
rect 162 184 164 186
rect 158 182 164 184
rect 168 186 174 188
rect 168 184 170 186
rect 172 184 174 186
rect 168 182 174 184
rect 122 179 124 182
rect 132 179 134 182
rect 152 179 154 182
rect 159 179 161 182
rect 60 161 62 166
rect 67 161 69 166
rect 80 164 82 168
rect 102 155 104 159
rect 112 157 114 162
rect 122 160 124 165
rect 132 160 134 165
rect 170 173 172 182
rect 191 181 193 194
rect 204 191 206 194
rect 293 219 295 223
rect 300 219 302 223
rect 370 219 372 223
rect 328 212 330 217
rect 338 212 340 217
rect 348 210 350 214
rect 328 196 330 199
rect 324 194 330 196
rect 324 192 326 194
rect 328 192 330 194
rect 197 189 206 191
rect 197 187 199 189
rect 201 187 203 189
rect 214 188 216 191
rect 221 188 223 191
rect 239 188 241 191
rect 249 188 251 191
rect 259 188 261 191
rect 280 188 282 191
rect 293 188 295 191
rect 300 188 302 191
rect 324 190 330 192
rect 197 185 203 187
rect 191 179 197 181
rect 191 177 193 179
rect 195 177 197 179
rect 191 175 197 177
rect 191 172 193 175
rect 201 172 203 185
rect 211 186 217 188
rect 211 184 213 186
rect 215 184 217 186
rect 211 182 217 184
rect 221 186 243 188
rect 221 184 232 186
rect 234 184 239 186
rect 241 184 243 186
rect 221 182 243 184
rect 247 186 253 188
rect 247 184 249 186
rect 251 184 253 186
rect 247 182 253 184
rect 257 186 263 188
rect 257 184 259 186
rect 261 184 263 186
rect 257 182 263 184
rect 280 186 286 188
rect 280 184 282 186
rect 284 184 286 186
rect 280 182 286 184
rect 290 186 296 188
rect 290 184 292 186
rect 294 184 296 186
rect 290 182 296 184
rect 300 186 309 188
rect 300 184 305 186
rect 307 184 309 186
rect 300 182 309 184
rect 211 179 213 182
rect 221 179 223 182
rect 241 179 243 182
rect 248 179 250 182
rect 152 155 154 159
rect 159 155 161 159
rect 170 155 172 159
rect 191 155 193 159
rect 201 157 203 162
rect 211 160 213 165
rect 221 160 223 165
rect 259 173 261 182
rect 280 179 282 182
rect 290 174 292 182
rect 300 176 302 182
rect 328 177 330 190
rect 338 188 340 199
rect 393 216 395 221
rect 400 216 402 221
rect 418 219 420 223
rect 428 219 430 223
rect 438 219 440 223
rect 459 219 461 223
rect 383 207 385 212
rect 348 188 350 192
rect 334 186 340 188
rect 334 184 336 186
rect 338 184 340 186
rect 334 182 340 184
rect 344 186 350 188
rect 344 184 346 186
rect 348 184 350 186
rect 344 182 350 184
rect 335 177 337 182
rect 348 177 350 182
rect 370 181 372 194
rect 383 191 385 194
rect 482 216 484 221
rect 489 216 491 221
rect 507 219 509 223
rect 517 219 519 223
rect 527 219 529 223
rect 548 219 550 223
rect 472 207 474 212
rect 376 189 385 191
rect 376 187 378 189
rect 380 187 382 189
rect 393 188 395 191
rect 400 188 402 191
rect 418 188 420 191
rect 428 188 430 191
rect 438 188 440 191
rect 376 185 382 187
rect 370 179 376 181
rect 370 177 372 179
rect 374 177 376 179
rect 280 160 282 165
rect 290 161 292 166
rect 300 164 302 168
rect 370 175 376 177
rect 370 172 372 175
rect 380 172 382 185
rect 390 186 396 188
rect 390 184 392 186
rect 394 184 396 186
rect 390 182 396 184
rect 400 186 422 188
rect 400 184 411 186
rect 413 184 418 186
rect 420 184 422 186
rect 400 182 422 184
rect 426 186 432 188
rect 426 184 428 186
rect 430 184 432 186
rect 426 182 432 184
rect 436 186 442 188
rect 436 184 438 186
rect 440 184 442 186
rect 436 182 442 184
rect 390 179 392 182
rect 400 179 402 182
rect 420 179 422 182
rect 427 179 429 182
rect 328 161 330 166
rect 335 161 337 166
rect 241 155 243 159
rect 248 155 250 159
rect 259 155 261 159
rect 348 164 350 168
rect 370 155 372 159
rect 380 157 382 162
rect 390 160 392 165
rect 400 160 402 165
rect 438 173 440 182
rect 459 181 461 194
rect 472 191 474 194
rect 561 219 563 223
rect 568 219 570 223
rect 637 219 639 223
rect 596 212 598 217
rect 606 212 608 217
rect 616 210 618 214
rect 596 196 598 199
rect 592 194 598 196
rect 592 192 594 194
rect 596 192 598 194
rect 465 189 474 191
rect 465 187 467 189
rect 469 187 471 189
rect 482 188 484 191
rect 489 188 491 191
rect 507 188 509 191
rect 517 188 519 191
rect 527 188 529 191
rect 548 188 550 191
rect 561 188 563 191
rect 568 188 570 191
rect 592 190 598 192
rect 465 185 471 187
rect 459 179 465 181
rect 459 177 461 179
rect 463 177 465 179
rect 459 175 465 177
rect 459 172 461 175
rect 469 172 471 185
rect 479 186 485 188
rect 479 184 481 186
rect 483 184 485 186
rect 479 182 485 184
rect 489 186 511 188
rect 489 184 500 186
rect 502 184 507 186
rect 509 184 511 186
rect 489 182 511 184
rect 515 186 521 188
rect 515 184 517 186
rect 519 184 521 186
rect 515 182 521 184
rect 525 186 531 188
rect 525 184 527 186
rect 529 184 531 186
rect 525 182 531 184
rect 548 186 554 188
rect 548 184 550 186
rect 552 184 554 186
rect 548 182 554 184
rect 558 186 564 188
rect 558 184 560 186
rect 562 184 564 186
rect 558 182 564 184
rect 568 186 577 188
rect 568 184 573 186
rect 575 184 577 186
rect 568 182 577 184
rect 479 179 481 182
rect 489 179 491 182
rect 509 179 511 182
rect 516 179 518 182
rect 420 155 422 159
rect 427 155 429 159
rect 438 155 440 159
rect 459 155 461 159
rect 469 157 471 162
rect 479 160 481 165
rect 489 160 491 165
rect 527 173 529 182
rect 548 179 550 182
rect 558 174 560 182
rect 568 176 570 182
rect 596 177 598 190
rect 606 188 608 199
rect 660 216 662 221
rect 667 216 669 221
rect 685 219 687 223
rect 695 219 697 223
rect 705 219 707 223
rect 726 219 728 223
rect 650 207 652 212
rect 616 188 618 192
rect 602 186 608 188
rect 602 184 604 186
rect 606 184 608 186
rect 602 182 608 184
rect 612 186 618 188
rect 612 184 614 186
rect 616 184 618 186
rect 612 182 618 184
rect 603 177 605 182
rect 616 177 618 182
rect 637 181 639 194
rect 650 191 652 194
rect 749 216 751 221
rect 756 216 758 221
rect 774 219 776 223
rect 784 219 786 223
rect 794 219 796 223
rect 815 219 817 223
rect 739 207 741 212
rect 643 189 652 191
rect 643 187 645 189
rect 647 187 649 189
rect 660 188 662 191
rect 667 188 669 191
rect 685 188 687 191
rect 695 188 697 191
rect 705 188 707 191
rect 643 185 649 187
rect 637 179 643 181
rect 637 177 639 179
rect 641 177 643 179
rect 548 160 550 165
rect 558 161 560 166
rect 568 164 570 168
rect 637 175 643 177
rect 637 172 639 175
rect 647 172 649 185
rect 657 186 663 188
rect 657 184 659 186
rect 661 184 663 186
rect 657 182 663 184
rect 667 186 689 188
rect 667 184 678 186
rect 680 184 685 186
rect 687 184 689 186
rect 667 182 689 184
rect 693 186 699 188
rect 693 184 695 186
rect 697 184 699 186
rect 693 182 699 184
rect 703 186 709 188
rect 703 184 705 186
rect 707 184 709 186
rect 703 182 709 184
rect 657 179 659 182
rect 667 179 669 182
rect 687 179 689 182
rect 694 179 696 182
rect 596 161 598 166
rect 603 161 605 166
rect 509 155 511 159
rect 516 155 518 159
rect 527 155 529 159
rect 616 164 618 168
rect 637 155 639 159
rect 647 157 649 162
rect 657 160 659 165
rect 667 160 669 165
rect 705 173 707 182
rect 726 181 728 194
rect 739 191 741 194
rect 828 219 830 223
rect 835 219 837 223
rect 732 189 741 191
rect 732 187 734 189
rect 736 187 738 189
rect 749 188 751 191
rect 756 188 758 191
rect 774 188 776 191
rect 784 188 786 191
rect 794 188 796 191
rect 815 188 817 191
rect 828 188 830 191
rect 835 188 837 191
rect 732 185 738 187
rect 726 179 732 181
rect 726 177 728 179
rect 730 177 732 179
rect 726 175 732 177
rect 726 172 728 175
rect 736 172 738 185
rect 746 186 752 188
rect 746 184 748 186
rect 750 184 752 186
rect 746 182 752 184
rect 756 186 778 188
rect 756 184 767 186
rect 769 184 774 186
rect 776 184 778 186
rect 756 182 778 184
rect 782 186 788 188
rect 782 184 784 186
rect 786 184 788 186
rect 782 182 788 184
rect 792 186 798 188
rect 792 184 794 186
rect 796 184 798 186
rect 792 182 798 184
rect 815 186 821 188
rect 815 184 817 186
rect 819 184 821 186
rect 815 182 821 184
rect 825 186 831 188
rect 825 184 827 186
rect 829 184 831 186
rect 825 182 831 184
rect 835 186 844 188
rect 835 184 840 186
rect 842 184 844 186
rect 835 182 844 184
rect 746 179 748 182
rect 756 179 758 182
rect 776 179 778 182
rect 783 179 785 182
rect 687 155 689 159
rect 694 155 696 159
rect 705 155 707 159
rect 726 155 728 159
rect 736 157 738 162
rect 746 160 748 165
rect 756 160 758 165
rect 794 173 796 182
rect 815 179 817 182
rect 825 174 827 182
rect 835 176 837 182
rect 815 160 817 165
rect 825 161 827 166
rect 835 164 837 168
rect 776 155 778 159
rect 783 155 785 159
rect 794 155 796 159
rect 20 140 22 145
rect 27 140 29 145
rect 40 138 42 142
rect 60 140 62 145
rect 67 140 69 145
rect 102 147 104 151
rect 80 138 82 142
rect 112 144 114 149
rect 152 147 154 151
rect 159 147 161 151
rect 170 147 172 151
rect 191 147 193 151
rect 122 141 124 146
rect 132 141 134 146
rect 102 131 104 134
rect 102 129 108 131
rect 20 116 22 129
rect 27 124 29 129
rect 40 124 42 129
rect 26 122 32 124
rect 26 120 28 122
rect 30 120 32 122
rect 26 118 32 120
rect 36 122 42 124
rect 36 120 38 122
rect 40 120 42 122
rect 36 118 42 120
rect 16 114 22 116
rect 16 112 18 114
rect 20 112 22 114
rect 16 110 22 112
rect 20 107 22 110
rect 30 107 32 118
rect 40 114 42 118
rect 60 116 62 129
rect 67 124 69 129
rect 80 124 82 129
rect 66 122 72 124
rect 66 120 68 122
rect 70 120 72 122
rect 66 118 72 120
rect 76 122 82 124
rect 76 120 78 122
rect 80 120 82 122
rect 76 118 82 120
rect 56 114 62 116
rect 56 112 58 114
rect 60 112 62 114
rect 56 110 62 112
rect 60 107 62 110
rect 70 107 72 118
rect 80 114 82 118
rect 102 127 104 129
rect 106 127 108 129
rect 102 125 108 127
rect 20 89 22 94
rect 30 89 32 94
rect 40 92 42 96
rect 102 112 104 125
rect 112 121 114 134
rect 201 144 203 149
rect 241 147 243 151
rect 248 147 250 151
rect 259 147 261 151
rect 211 141 213 146
rect 221 141 223 146
rect 108 119 114 121
rect 108 117 110 119
rect 112 117 114 119
rect 122 124 124 127
rect 132 124 134 127
rect 152 124 154 127
rect 159 124 161 127
rect 170 124 172 133
rect 191 131 193 134
rect 191 129 197 131
rect 191 127 193 129
rect 195 127 197 129
rect 191 125 197 127
rect 122 122 128 124
rect 122 120 124 122
rect 126 120 128 122
rect 122 118 128 120
rect 132 122 154 124
rect 132 120 143 122
rect 145 120 150 122
rect 152 120 154 122
rect 132 118 154 120
rect 158 122 164 124
rect 158 120 160 122
rect 162 120 164 122
rect 158 118 164 120
rect 168 122 174 124
rect 168 120 170 122
rect 172 120 174 122
rect 168 118 174 120
rect 108 115 117 117
rect 125 115 127 118
rect 132 115 134 118
rect 150 115 152 118
rect 160 115 162 118
rect 170 115 172 118
rect 115 112 117 115
rect 60 89 62 94
rect 70 89 72 94
rect 80 92 82 96
rect 115 94 117 99
rect 102 83 104 87
rect 125 85 127 90
rect 132 85 134 90
rect 191 112 193 125
rect 201 121 203 134
rect 280 141 282 146
rect 197 119 203 121
rect 197 117 199 119
rect 201 117 203 119
rect 211 124 213 127
rect 221 124 223 127
rect 241 124 243 127
rect 248 124 250 127
rect 259 124 261 133
rect 290 140 292 145
rect 300 138 302 142
rect 328 140 330 145
rect 335 140 337 145
rect 370 147 372 151
rect 280 124 282 127
rect 290 124 292 132
rect 300 124 302 130
rect 348 138 350 142
rect 380 144 382 149
rect 420 147 422 151
rect 427 147 429 151
rect 438 147 440 151
rect 459 147 461 151
rect 390 141 392 146
rect 400 141 402 146
rect 370 131 372 134
rect 370 129 376 131
rect 211 122 217 124
rect 211 120 213 122
rect 215 120 217 122
rect 211 118 217 120
rect 221 122 243 124
rect 221 120 232 122
rect 234 120 239 122
rect 241 120 243 122
rect 221 118 243 120
rect 247 122 253 124
rect 247 120 249 122
rect 251 120 253 122
rect 247 118 253 120
rect 257 122 263 124
rect 257 120 259 122
rect 261 120 263 122
rect 257 118 263 120
rect 280 122 286 124
rect 280 120 282 122
rect 284 120 286 122
rect 280 118 286 120
rect 290 122 296 124
rect 290 120 292 122
rect 294 120 296 122
rect 290 118 296 120
rect 300 122 309 124
rect 300 120 305 122
rect 307 120 309 122
rect 300 118 309 120
rect 197 115 206 117
rect 214 115 216 118
rect 221 115 223 118
rect 239 115 241 118
rect 249 115 251 118
rect 259 115 261 118
rect 280 115 282 118
rect 293 115 295 118
rect 300 115 302 118
rect 328 116 330 129
rect 335 124 337 129
rect 348 124 350 129
rect 334 122 340 124
rect 334 120 336 122
rect 338 120 340 122
rect 334 118 340 120
rect 344 122 350 124
rect 344 120 346 122
rect 348 120 350 122
rect 344 118 350 120
rect 204 112 206 115
rect 204 94 206 99
rect 150 83 152 87
rect 160 83 162 87
rect 170 83 172 87
rect 191 83 193 87
rect 214 85 216 90
rect 221 85 223 90
rect 239 83 241 87
rect 249 83 251 87
rect 259 83 261 87
rect 280 83 282 87
rect 324 114 330 116
rect 324 112 326 114
rect 328 112 330 114
rect 324 110 330 112
rect 328 107 330 110
rect 338 107 340 118
rect 348 114 350 118
rect 370 127 372 129
rect 374 127 376 129
rect 370 125 376 127
rect 370 112 372 125
rect 380 121 382 134
rect 469 144 471 149
rect 509 147 511 151
rect 516 147 518 151
rect 527 147 529 151
rect 479 141 481 146
rect 489 141 491 146
rect 376 119 382 121
rect 376 117 378 119
rect 380 117 382 119
rect 390 124 392 127
rect 400 124 402 127
rect 420 124 422 127
rect 427 124 429 127
rect 438 124 440 133
rect 459 131 461 134
rect 459 129 465 131
rect 459 127 461 129
rect 463 127 465 129
rect 459 125 465 127
rect 390 122 396 124
rect 390 120 392 122
rect 394 120 396 122
rect 390 118 396 120
rect 400 122 422 124
rect 400 120 411 122
rect 413 120 418 122
rect 420 120 422 122
rect 400 118 422 120
rect 426 122 432 124
rect 426 120 428 122
rect 430 120 432 122
rect 426 118 432 120
rect 436 122 442 124
rect 436 120 438 122
rect 440 120 442 122
rect 436 118 442 120
rect 376 115 385 117
rect 393 115 395 118
rect 400 115 402 118
rect 418 115 420 118
rect 428 115 430 118
rect 438 115 440 118
rect 383 112 385 115
rect 328 89 330 94
rect 338 89 340 94
rect 348 92 350 96
rect 293 83 295 87
rect 300 83 302 87
rect 383 94 385 99
rect 370 83 372 87
rect 393 85 395 90
rect 400 85 402 90
rect 459 112 461 125
rect 469 121 471 134
rect 548 141 550 146
rect 465 119 471 121
rect 465 117 467 119
rect 469 117 471 119
rect 479 124 481 127
rect 489 124 491 127
rect 509 124 511 127
rect 516 124 518 127
rect 527 124 529 133
rect 558 140 560 145
rect 568 138 570 142
rect 596 140 598 145
rect 603 140 605 145
rect 637 147 639 151
rect 548 124 550 127
rect 558 124 560 132
rect 568 124 570 130
rect 616 138 618 142
rect 647 144 649 149
rect 687 147 689 151
rect 694 147 696 151
rect 705 147 707 151
rect 726 147 728 151
rect 657 141 659 146
rect 667 141 669 146
rect 637 131 639 134
rect 637 129 643 131
rect 479 122 485 124
rect 479 120 481 122
rect 483 120 485 122
rect 479 118 485 120
rect 489 122 511 124
rect 489 120 500 122
rect 502 120 507 122
rect 509 120 511 122
rect 489 118 511 120
rect 515 122 521 124
rect 515 120 517 122
rect 519 120 521 122
rect 515 118 521 120
rect 525 122 531 124
rect 525 120 527 122
rect 529 120 531 122
rect 525 118 531 120
rect 548 122 554 124
rect 548 120 550 122
rect 552 120 554 122
rect 548 118 554 120
rect 558 122 564 124
rect 558 120 560 122
rect 562 120 564 122
rect 558 118 564 120
rect 568 122 577 124
rect 568 120 573 122
rect 575 120 577 122
rect 568 118 577 120
rect 465 115 474 117
rect 482 115 484 118
rect 489 115 491 118
rect 507 115 509 118
rect 517 115 519 118
rect 527 115 529 118
rect 548 115 550 118
rect 561 115 563 118
rect 568 115 570 118
rect 596 116 598 129
rect 603 124 605 129
rect 616 124 618 129
rect 602 122 608 124
rect 602 120 604 122
rect 606 120 608 122
rect 602 118 608 120
rect 612 122 618 124
rect 612 120 614 122
rect 616 120 618 122
rect 612 118 618 120
rect 472 112 474 115
rect 472 94 474 99
rect 418 83 420 87
rect 428 83 430 87
rect 438 83 440 87
rect 459 83 461 87
rect 482 85 484 90
rect 489 85 491 90
rect 507 83 509 87
rect 517 83 519 87
rect 527 83 529 87
rect 548 83 550 87
rect 592 114 598 116
rect 592 112 594 114
rect 596 112 598 114
rect 592 110 598 112
rect 596 107 598 110
rect 606 107 608 118
rect 616 114 618 118
rect 637 127 639 129
rect 641 127 643 129
rect 637 125 643 127
rect 637 112 639 125
rect 647 121 649 134
rect 736 144 738 149
rect 776 147 778 151
rect 783 147 785 151
rect 794 147 796 151
rect 746 141 748 146
rect 756 141 758 146
rect 643 119 649 121
rect 643 117 645 119
rect 647 117 649 119
rect 657 124 659 127
rect 667 124 669 127
rect 687 124 689 127
rect 694 124 696 127
rect 705 124 707 133
rect 726 131 728 134
rect 726 129 732 131
rect 726 127 728 129
rect 730 127 732 129
rect 726 125 732 127
rect 657 122 663 124
rect 657 120 659 122
rect 661 120 663 122
rect 657 118 663 120
rect 667 122 689 124
rect 667 120 678 122
rect 680 120 685 122
rect 687 120 689 122
rect 667 118 689 120
rect 693 122 699 124
rect 693 120 695 122
rect 697 120 699 122
rect 693 118 699 120
rect 703 122 709 124
rect 703 120 705 122
rect 707 120 709 122
rect 703 118 709 120
rect 643 115 652 117
rect 660 115 662 118
rect 667 115 669 118
rect 685 115 687 118
rect 695 115 697 118
rect 705 115 707 118
rect 650 112 652 115
rect 596 89 598 94
rect 606 89 608 94
rect 616 92 618 96
rect 561 83 563 87
rect 568 83 570 87
rect 650 94 652 99
rect 637 83 639 87
rect 660 85 662 90
rect 667 85 669 90
rect 726 112 728 125
rect 736 121 738 134
rect 815 141 817 146
rect 732 119 738 121
rect 732 117 734 119
rect 736 117 738 119
rect 746 124 748 127
rect 756 124 758 127
rect 776 124 778 127
rect 783 124 785 127
rect 794 124 796 133
rect 825 140 827 145
rect 835 138 837 142
rect 815 124 817 127
rect 825 124 827 132
rect 835 124 837 130
rect 746 122 752 124
rect 746 120 748 122
rect 750 120 752 122
rect 746 118 752 120
rect 756 122 778 124
rect 756 120 767 122
rect 769 120 774 122
rect 776 120 778 122
rect 756 118 778 120
rect 782 122 788 124
rect 782 120 784 122
rect 786 120 788 122
rect 782 118 788 120
rect 792 122 798 124
rect 792 120 794 122
rect 796 120 798 122
rect 792 118 798 120
rect 815 122 821 124
rect 815 120 817 122
rect 819 120 821 122
rect 815 118 821 120
rect 825 122 831 124
rect 825 120 827 122
rect 829 120 831 122
rect 825 118 831 120
rect 835 122 844 124
rect 835 120 840 122
rect 842 120 844 122
rect 835 118 844 120
rect 732 115 741 117
rect 749 115 751 118
rect 756 115 758 118
rect 774 115 776 118
rect 784 115 786 118
rect 794 115 796 118
rect 815 115 817 118
rect 828 115 830 118
rect 835 115 837 118
rect 739 112 741 115
rect 739 94 741 99
rect 685 83 687 87
rect 695 83 697 87
rect 705 83 707 87
rect 726 83 728 87
rect 749 85 751 90
rect 756 85 758 90
rect 774 83 776 87
rect 784 83 786 87
rect 794 83 796 87
rect 815 83 817 87
rect 828 83 830 87
rect 835 83 837 87
rect 20 68 22 73
rect 30 68 32 73
rect 102 75 104 79
rect 40 66 42 70
rect 60 68 62 73
rect 70 68 72 73
rect 20 52 22 55
rect 16 50 22 52
rect 16 48 18 50
rect 20 48 22 50
rect 16 46 22 48
rect 20 33 22 46
rect 30 44 32 55
rect 80 66 82 70
rect 60 52 62 55
rect 56 50 62 52
rect 56 48 58 50
rect 60 48 62 50
rect 40 44 42 48
rect 56 46 62 48
rect 26 42 32 44
rect 26 40 28 42
rect 30 40 32 42
rect 26 38 32 40
rect 36 42 42 44
rect 36 40 38 42
rect 40 40 42 42
rect 36 38 42 40
rect 27 33 29 38
rect 40 33 42 38
rect 60 33 62 46
rect 70 44 72 55
rect 125 72 127 77
rect 132 72 134 77
rect 150 75 152 79
rect 160 75 162 79
rect 170 75 172 79
rect 191 75 193 79
rect 115 63 117 68
rect 80 44 82 48
rect 66 42 72 44
rect 66 40 68 42
rect 70 40 72 42
rect 66 38 72 40
rect 76 42 82 44
rect 76 40 78 42
rect 80 40 82 42
rect 76 38 82 40
rect 67 33 69 38
rect 80 33 82 38
rect 102 37 104 50
rect 115 47 117 50
rect 214 72 216 77
rect 221 72 223 77
rect 239 75 241 79
rect 249 75 251 79
rect 259 75 261 79
rect 280 75 282 79
rect 204 63 206 68
rect 108 45 117 47
rect 108 43 110 45
rect 112 43 114 45
rect 125 44 127 47
rect 132 44 134 47
rect 150 44 152 47
rect 160 44 162 47
rect 170 44 172 47
rect 108 41 114 43
rect 102 35 108 37
rect 102 33 104 35
rect 106 33 108 35
rect 20 17 22 22
rect 27 17 29 22
rect 40 20 42 24
rect 102 31 108 33
rect 102 28 104 31
rect 112 28 114 41
rect 122 42 128 44
rect 122 40 124 42
rect 126 40 128 42
rect 122 38 128 40
rect 132 42 154 44
rect 132 40 143 42
rect 145 40 150 42
rect 152 40 154 42
rect 132 38 154 40
rect 158 42 164 44
rect 158 40 160 42
rect 162 40 164 42
rect 158 38 164 40
rect 168 42 174 44
rect 168 40 170 42
rect 172 40 174 42
rect 168 38 174 40
rect 122 35 124 38
rect 132 35 134 38
rect 152 35 154 38
rect 159 35 161 38
rect 60 17 62 22
rect 67 17 69 22
rect 80 20 82 24
rect 102 11 104 15
rect 112 13 114 18
rect 122 16 124 21
rect 132 16 134 21
rect 170 29 172 38
rect 191 37 193 50
rect 204 47 206 50
rect 293 75 295 79
rect 300 75 302 79
rect 370 75 372 79
rect 328 68 330 73
rect 338 68 340 73
rect 348 66 350 70
rect 328 52 330 55
rect 324 50 330 52
rect 324 48 326 50
rect 328 48 330 50
rect 197 45 206 47
rect 197 43 199 45
rect 201 43 203 45
rect 214 44 216 47
rect 221 44 223 47
rect 239 44 241 47
rect 249 44 251 47
rect 259 44 261 47
rect 280 44 282 47
rect 293 44 295 47
rect 300 44 302 47
rect 324 46 330 48
rect 197 41 203 43
rect 191 35 197 37
rect 191 33 193 35
rect 195 33 197 35
rect 191 31 197 33
rect 191 28 193 31
rect 201 28 203 41
rect 211 42 217 44
rect 211 40 213 42
rect 215 40 217 42
rect 211 38 217 40
rect 221 42 243 44
rect 221 40 232 42
rect 234 40 239 42
rect 241 40 243 42
rect 221 38 243 40
rect 247 42 253 44
rect 247 40 249 42
rect 251 40 253 42
rect 247 38 253 40
rect 257 42 263 44
rect 257 40 259 42
rect 261 40 263 42
rect 257 38 263 40
rect 280 42 286 44
rect 280 40 282 42
rect 284 40 286 42
rect 280 38 286 40
rect 290 42 296 44
rect 290 40 292 42
rect 294 40 296 42
rect 290 38 296 40
rect 300 42 309 44
rect 300 40 305 42
rect 307 40 309 42
rect 300 38 309 40
rect 211 35 213 38
rect 221 35 223 38
rect 241 35 243 38
rect 248 35 250 38
rect 152 11 154 15
rect 159 11 161 15
rect 170 11 172 15
rect 191 11 193 15
rect 201 13 203 18
rect 211 16 213 21
rect 221 16 223 21
rect 259 29 261 38
rect 280 35 282 38
rect 290 30 292 38
rect 300 32 302 38
rect 328 33 330 46
rect 338 44 340 55
rect 393 72 395 77
rect 400 72 402 77
rect 418 75 420 79
rect 428 75 430 79
rect 438 75 440 79
rect 459 75 461 79
rect 383 63 385 68
rect 348 44 350 48
rect 334 42 340 44
rect 334 40 336 42
rect 338 40 340 42
rect 334 38 340 40
rect 344 42 350 44
rect 344 40 346 42
rect 348 40 350 42
rect 344 38 350 40
rect 335 33 337 38
rect 348 33 350 38
rect 370 37 372 50
rect 383 47 385 50
rect 482 72 484 77
rect 489 72 491 77
rect 507 75 509 79
rect 517 75 519 79
rect 527 75 529 79
rect 548 75 550 79
rect 472 63 474 68
rect 376 45 385 47
rect 376 43 378 45
rect 380 43 382 45
rect 393 44 395 47
rect 400 44 402 47
rect 418 44 420 47
rect 428 44 430 47
rect 438 44 440 47
rect 376 41 382 43
rect 370 35 376 37
rect 370 33 372 35
rect 374 33 376 35
rect 280 16 282 21
rect 290 17 292 22
rect 300 20 302 24
rect 370 31 376 33
rect 370 28 372 31
rect 380 28 382 41
rect 390 42 396 44
rect 390 40 392 42
rect 394 40 396 42
rect 390 38 396 40
rect 400 42 422 44
rect 400 40 411 42
rect 413 40 418 42
rect 420 40 422 42
rect 400 38 422 40
rect 426 42 432 44
rect 426 40 428 42
rect 430 40 432 42
rect 426 38 432 40
rect 436 42 442 44
rect 436 40 438 42
rect 440 40 442 42
rect 436 38 442 40
rect 390 35 392 38
rect 400 35 402 38
rect 420 35 422 38
rect 427 35 429 38
rect 328 17 330 22
rect 335 17 337 22
rect 241 11 243 15
rect 248 11 250 15
rect 259 11 261 15
rect 348 20 350 24
rect 370 11 372 15
rect 380 13 382 18
rect 390 16 392 21
rect 400 16 402 21
rect 438 29 440 38
rect 459 37 461 50
rect 472 47 474 50
rect 561 75 563 79
rect 568 75 570 79
rect 637 75 639 79
rect 596 68 598 73
rect 606 68 608 73
rect 616 66 618 70
rect 596 52 598 55
rect 592 50 598 52
rect 592 48 594 50
rect 596 48 598 50
rect 465 45 474 47
rect 465 43 467 45
rect 469 43 471 45
rect 482 44 484 47
rect 489 44 491 47
rect 507 44 509 47
rect 517 44 519 47
rect 527 44 529 47
rect 548 44 550 47
rect 561 44 563 47
rect 568 44 570 47
rect 592 46 598 48
rect 465 41 471 43
rect 459 35 465 37
rect 459 33 461 35
rect 463 33 465 35
rect 459 31 465 33
rect 459 28 461 31
rect 469 28 471 41
rect 479 42 485 44
rect 479 40 481 42
rect 483 40 485 42
rect 479 38 485 40
rect 489 42 511 44
rect 489 40 500 42
rect 502 40 507 42
rect 509 40 511 42
rect 489 38 511 40
rect 515 42 521 44
rect 515 40 517 42
rect 519 40 521 42
rect 515 38 521 40
rect 525 42 531 44
rect 525 40 527 42
rect 529 40 531 42
rect 525 38 531 40
rect 548 42 554 44
rect 548 40 550 42
rect 552 40 554 42
rect 548 38 554 40
rect 558 42 564 44
rect 558 40 560 42
rect 562 40 564 42
rect 558 38 564 40
rect 568 42 577 44
rect 568 40 573 42
rect 575 40 577 42
rect 568 38 577 40
rect 479 35 481 38
rect 489 35 491 38
rect 509 35 511 38
rect 516 35 518 38
rect 420 11 422 15
rect 427 11 429 15
rect 438 11 440 15
rect 459 11 461 15
rect 469 13 471 18
rect 479 16 481 21
rect 489 16 491 21
rect 527 29 529 38
rect 548 35 550 38
rect 558 30 560 38
rect 568 32 570 38
rect 596 33 598 46
rect 606 44 608 55
rect 660 72 662 77
rect 667 72 669 77
rect 685 75 687 79
rect 695 75 697 79
rect 705 75 707 79
rect 726 75 728 79
rect 650 63 652 68
rect 616 44 618 48
rect 602 42 608 44
rect 602 40 604 42
rect 606 40 608 42
rect 602 38 608 40
rect 612 42 618 44
rect 612 40 614 42
rect 616 40 618 42
rect 612 38 618 40
rect 603 33 605 38
rect 616 33 618 38
rect 637 37 639 50
rect 650 47 652 50
rect 749 72 751 77
rect 756 72 758 77
rect 774 75 776 79
rect 784 75 786 79
rect 794 75 796 79
rect 815 75 817 79
rect 739 63 741 68
rect 643 45 652 47
rect 643 43 645 45
rect 647 43 649 45
rect 660 44 662 47
rect 667 44 669 47
rect 685 44 687 47
rect 695 44 697 47
rect 705 44 707 47
rect 643 41 649 43
rect 637 35 643 37
rect 637 33 639 35
rect 641 33 643 35
rect 548 16 550 21
rect 558 17 560 22
rect 568 20 570 24
rect 637 31 643 33
rect 637 28 639 31
rect 647 28 649 41
rect 657 42 663 44
rect 657 40 659 42
rect 661 40 663 42
rect 657 38 663 40
rect 667 42 689 44
rect 667 40 678 42
rect 680 40 685 42
rect 687 40 689 42
rect 667 38 689 40
rect 693 42 699 44
rect 693 40 695 42
rect 697 40 699 42
rect 693 38 699 40
rect 703 42 709 44
rect 703 40 705 42
rect 707 40 709 42
rect 703 38 709 40
rect 657 35 659 38
rect 667 35 669 38
rect 687 35 689 38
rect 694 35 696 38
rect 596 17 598 22
rect 603 17 605 22
rect 509 11 511 15
rect 516 11 518 15
rect 527 11 529 15
rect 616 20 618 24
rect 637 11 639 15
rect 647 13 649 18
rect 657 16 659 21
rect 667 16 669 21
rect 705 29 707 38
rect 726 37 728 50
rect 739 47 741 50
rect 828 75 830 79
rect 835 75 837 79
rect 732 45 741 47
rect 732 43 734 45
rect 736 43 738 45
rect 749 44 751 47
rect 756 44 758 47
rect 774 44 776 47
rect 784 44 786 47
rect 794 44 796 47
rect 815 44 817 47
rect 828 44 830 47
rect 835 44 837 47
rect 732 41 738 43
rect 726 35 732 37
rect 726 33 728 35
rect 730 33 732 35
rect 726 31 732 33
rect 726 28 728 31
rect 736 28 738 41
rect 746 42 752 44
rect 746 40 748 42
rect 750 40 752 42
rect 746 38 752 40
rect 756 42 778 44
rect 756 40 767 42
rect 769 40 774 42
rect 776 40 778 42
rect 756 38 778 40
rect 782 42 788 44
rect 782 40 784 42
rect 786 40 788 42
rect 782 38 788 40
rect 792 42 798 44
rect 792 40 794 42
rect 796 40 798 42
rect 792 38 798 40
rect 815 42 821 44
rect 815 40 817 42
rect 819 40 821 42
rect 815 38 821 40
rect 825 42 831 44
rect 825 40 827 42
rect 829 40 831 42
rect 825 38 831 40
rect 835 42 844 44
rect 835 40 840 42
rect 842 40 844 42
rect 835 38 844 40
rect 746 35 748 38
rect 756 35 758 38
rect 776 35 778 38
rect 783 35 785 38
rect 687 11 689 15
rect 694 11 696 15
rect 705 11 707 15
rect 726 11 728 15
rect 736 13 738 18
rect 746 16 748 21
rect 756 16 758 21
rect 794 29 796 38
rect 815 35 817 38
rect 825 30 827 38
rect 835 32 837 38
rect 815 16 817 21
rect 825 17 827 22
rect 835 20 837 24
rect 776 11 778 15
rect 783 11 785 15
rect 794 11 796 15
<< ndif >>
rect 31 292 38 294
rect 31 290 34 292
rect 36 290 38 292
rect 31 284 38 290
rect 71 292 78 294
rect 71 290 74 292
rect 76 290 78 292
rect 13 282 20 284
rect 13 280 15 282
rect 17 280 20 282
rect 13 278 20 280
rect 15 273 20 278
rect 22 273 27 284
rect 29 282 38 284
rect 71 284 78 290
rect 53 282 60 284
rect 29 273 40 282
rect 42 280 49 282
rect 42 278 45 280
rect 47 278 49 280
rect 53 280 55 282
rect 57 280 60 282
rect 53 278 60 280
rect 42 276 49 278
rect 42 273 47 276
rect 55 273 60 278
rect 62 273 67 284
rect 69 282 78 284
rect 97 284 102 291
rect 95 282 102 284
rect 69 273 80 282
rect 82 280 89 282
rect 82 278 85 280
rect 87 278 89 280
rect 95 280 97 282
rect 99 280 102 282
rect 95 278 102 280
rect 104 288 109 291
rect 104 286 112 288
rect 104 284 107 286
rect 109 284 112 286
rect 104 278 112 284
rect 114 285 119 288
rect 114 283 122 285
rect 114 281 117 283
rect 119 281 122 283
rect 114 278 122 281
rect 82 276 89 278
rect 82 273 87 276
rect 117 271 122 278
rect 124 275 132 285
rect 124 273 127 275
rect 129 273 132 275
rect 124 271 132 273
rect 134 282 141 285
rect 147 284 152 291
rect 134 280 137 282
rect 139 280 141 282
rect 134 275 141 280
rect 145 282 152 284
rect 145 280 147 282
rect 149 280 152 282
rect 145 278 152 280
rect 134 273 137 275
rect 139 273 141 275
rect 134 271 141 273
rect 147 271 152 278
rect 154 271 159 291
rect 161 289 170 291
rect 161 287 164 289
rect 166 287 170 289
rect 161 277 170 287
rect 172 284 177 291
rect 186 284 191 291
rect 172 282 179 284
rect 172 280 175 282
rect 177 280 179 282
rect 172 277 179 280
rect 184 282 191 284
rect 184 280 186 282
rect 188 280 191 282
rect 184 278 191 280
rect 193 288 198 291
rect 193 286 201 288
rect 193 284 196 286
rect 198 284 201 286
rect 193 278 201 284
rect 203 285 208 288
rect 203 283 211 285
rect 203 281 206 283
rect 208 281 211 283
rect 203 278 211 281
rect 161 271 168 277
rect 206 271 211 278
rect 213 275 221 285
rect 213 273 216 275
rect 218 273 221 275
rect 213 271 221 273
rect 223 282 230 285
rect 236 284 241 291
rect 223 280 226 282
rect 228 280 230 282
rect 223 275 230 280
rect 234 282 241 284
rect 234 280 236 282
rect 238 280 241 282
rect 234 278 241 280
rect 223 273 226 275
rect 228 273 230 275
rect 223 271 230 273
rect 236 271 241 278
rect 243 271 248 291
rect 250 289 259 291
rect 250 287 253 289
rect 255 287 259 289
rect 250 277 259 287
rect 261 284 266 291
rect 261 282 268 284
rect 261 280 264 282
rect 266 280 268 282
rect 261 277 268 280
rect 273 282 280 285
rect 273 280 275 282
rect 277 280 280 282
rect 250 271 257 277
rect 273 275 280 280
rect 273 273 275 275
rect 277 273 280 275
rect 273 271 280 273
rect 282 284 287 285
rect 339 292 346 294
rect 339 290 342 292
rect 344 290 346 292
rect 282 282 290 284
rect 282 280 285 282
rect 287 280 290 282
rect 282 276 290 280
rect 292 282 297 284
rect 339 284 346 290
rect 321 282 328 284
rect 292 280 300 282
rect 292 278 295 280
rect 297 278 300 280
rect 292 276 300 278
rect 282 271 287 276
rect 295 274 300 276
rect 302 280 309 282
rect 302 278 305 280
rect 307 278 309 280
rect 321 280 323 282
rect 325 280 328 282
rect 321 278 328 280
rect 302 274 309 278
rect 323 273 328 278
rect 330 273 335 284
rect 337 282 346 284
rect 365 284 370 291
rect 363 282 370 284
rect 337 273 348 282
rect 350 280 357 282
rect 350 278 353 280
rect 355 278 357 280
rect 363 280 365 282
rect 367 280 370 282
rect 363 278 370 280
rect 372 288 377 291
rect 372 286 380 288
rect 372 284 375 286
rect 377 284 380 286
rect 372 278 380 284
rect 382 285 387 288
rect 382 283 390 285
rect 382 281 385 283
rect 387 281 390 283
rect 382 278 390 281
rect 350 276 357 278
rect 350 273 355 276
rect 385 271 390 278
rect 392 275 400 285
rect 392 273 395 275
rect 397 273 400 275
rect 392 271 400 273
rect 402 282 409 285
rect 415 284 420 291
rect 402 280 405 282
rect 407 280 409 282
rect 402 275 409 280
rect 413 282 420 284
rect 413 280 415 282
rect 417 280 420 282
rect 413 278 420 280
rect 402 273 405 275
rect 407 273 409 275
rect 402 271 409 273
rect 415 271 420 278
rect 422 271 427 291
rect 429 289 438 291
rect 429 287 432 289
rect 434 287 438 289
rect 429 277 438 287
rect 440 284 445 291
rect 454 284 459 291
rect 440 282 447 284
rect 440 280 443 282
rect 445 280 447 282
rect 440 277 447 280
rect 452 282 459 284
rect 452 280 454 282
rect 456 280 459 282
rect 452 278 459 280
rect 461 288 466 291
rect 461 286 469 288
rect 461 284 464 286
rect 466 284 469 286
rect 461 278 469 284
rect 471 285 476 288
rect 471 283 479 285
rect 471 281 474 283
rect 476 281 479 283
rect 471 278 479 281
rect 429 271 436 277
rect 474 271 479 278
rect 481 275 489 285
rect 481 273 484 275
rect 486 273 489 275
rect 481 271 489 273
rect 491 282 498 285
rect 504 284 509 291
rect 491 280 494 282
rect 496 280 498 282
rect 491 275 498 280
rect 502 282 509 284
rect 502 280 504 282
rect 506 280 509 282
rect 502 278 509 280
rect 491 273 494 275
rect 496 273 498 275
rect 491 271 498 273
rect 504 271 509 278
rect 511 271 516 291
rect 518 289 527 291
rect 518 287 521 289
rect 523 287 527 289
rect 518 277 527 287
rect 529 284 534 291
rect 529 282 536 284
rect 529 280 532 282
rect 534 280 536 282
rect 529 277 536 280
rect 541 282 548 285
rect 541 280 543 282
rect 545 280 548 282
rect 518 271 525 277
rect 541 275 548 280
rect 541 273 543 275
rect 545 273 548 275
rect 541 271 548 273
rect 550 284 555 285
rect 607 292 614 294
rect 607 290 610 292
rect 612 290 614 292
rect 550 282 558 284
rect 550 280 553 282
rect 555 280 558 282
rect 550 276 558 280
rect 560 282 565 284
rect 607 284 614 290
rect 589 282 596 284
rect 560 280 568 282
rect 560 278 563 280
rect 565 278 568 280
rect 560 276 568 278
rect 550 271 555 276
rect 563 274 568 276
rect 570 280 577 282
rect 570 278 573 280
rect 575 278 577 280
rect 589 280 591 282
rect 593 280 596 282
rect 589 278 596 280
rect 570 274 577 278
rect 591 273 596 278
rect 598 273 603 284
rect 605 282 614 284
rect 632 284 637 291
rect 630 282 637 284
rect 605 273 616 282
rect 618 280 625 282
rect 618 278 621 280
rect 623 278 625 280
rect 630 280 632 282
rect 634 280 637 282
rect 630 278 637 280
rect 639 288 644 291
rect 639 286 647 288
rect 639 284 642 286
rect 644 284 647 286
rect 639 278 647 284
rect 649 285 654 288
rect 649 283 657 285
rect 649 281 652 283
rect 654 281 657 283
rect 649 278 657 281
rect 618 276 625 278
rect 618 273 623 276
rect 652 271 657 278
rect 659 275 667 285
rect 659 273 662 275
rect 664 273 667 275
rect 659 271 667 273
rect 669 282 676 285
rect 682 284 687 291
rect 669 280 672 282
rect 674 280 676 282
rect 669 275 676 280
rect 680 282 687 284
rect 680 280 682 282
rect 684 280 687 282
rect 680 278 687 280
rect 669 273 672 275
rect 674 273 676 275
rect 669 271 676 273
rect 682 271 687 278
rect 689 271 694 291
rect 696 289 705 291
rect 696 287 699 289
rect 701 287 705 289
rect 696 277 705 287
rect 707 284 712 291
rect 721 284 726 291
rect 707 282 714 284
rect 707 280 710 282
rect 712 280 714 282
rect 707 277 714 280
rect 719 282 726 284
rect 719 280 721 282
rect 723 280 726 282
rect 719 278 726 280
rect 728 288 733 291
rect 728 286 736 288
rect 728 284 731 286
rect 733 284 736 286
rect 728 278 736 284
rect 738 285 743 288
rect 738 283 746 285
rect 738 281 741 283
rect 743 281 746 283
rect 738 278 746 281
rect 696 271 703 277
rect 741 271 746 278
rect 748 275 756 285
rect 748 273 751 275
rect 753 273 756 275
rect 748 271 756 273
rect 758 282 765 285
rect 771 284 776 291
rect 758 280 761 282
rect 763 280 765 282
rect 758 275 765 280
rect 769 282 776 284
rect 769 280 771 282
rect 773 280 776 282
rect 769 278 776 280
rect 758 273 761 275
rect 763 273 765 275
rect 758 271 765 273
rect 771 271 776 278
rect 778 271 783 291
rect 785 289 794 291
rect 785 287 788 289
rect 790 287 794 289
rect 785 277 794 287
rect 796 284 801 291
rect 796 282 803 284
rect 796 280 799 282
rect 801 280 803 282
rect 796 277 803 280
rect 808 282 815 285
rect 808 280 810 282
rect 812 280 815 282
rect 785 271 792 277
rect 808 275 815 280
rect 808 273 810 275
rect 812 273 815 275
rect 808 271 815 273
rect 817 284 822 285
rect 817 282 825 284
rect 817 280 820 282
rect 822 280 825 282
rect 817 276 825 280
rect 827 282 832 284
rect 827 280 835 282
rect 827 278 830 280
rect 832 278 835 280
rect 827 276 835 278
rect 817 271 822 276
rect 830 274 835 276
rect 837 280 844 282
rect 837 278 840 280
rect 842 278 844 280
rect 837 274 844 278
rect 15 172 20 177
rect 13 170 20 172
rect 13 168 15 170
rect 17 168 20 170
rect 13 166 20 168
rect 22 166 27 177
rect 29 168 40 177
rect 42 174 47 177
rect 42 172 49 174
rect 55 172 60 177
rect 42 170 45 172
rect 47 170 49 172
rect 42 168 49 170
rect 53 170 60 172
rect 53 168 55 170
rect 57 168 60 170
rect 29 166 38 168
rect 31 160 38 166
rect 53 166 60 168
rect 62 166 67 177
rect 69 168 80 177
rect 82 174 87 177
rect 82 172 89 174
rect 117 172 122 179
rect 82 170 85 172
rect 87 170 89 172
rect 82 168 89 170
rect 95 170 102 172
rect 95 168 97 170
rect 99 168 102 170
rect 69 166 78 168
rect 31 158 34 160
rect 36 158 38 160
rect 31 156 38 158
rect 71 160 78 166
rect 95 166 102 168
rect 71 158 74 160
rect 76 158 78 160
rect 71 156 78 158
rect 97 159 102 166
rect 104 166 112 172
rect 104 164 107 166
rect 109 164 112 166
rect 104 162 112 164
rect 114 169 122 172
rect 114 167 117 169
rect 119 167 122 169
rect 114 165 122 167
rect 124 177 132 179
rect 124 175 127 177
rect 129 175 132 177
rect 124 165 132 175
rect 134 177 141 179
rect 134 175 137 177
rect 139 175 141 177
rect 134 170 141 175
rect 147 172 152 179
rect 134 168 137 170
rect 139 168 141 170
rect 134 165 141 168
rect 145 170 152 172
rect 145 168 147 170
rect 149 168 152 170
rect 145 166 152 168
rect 114 162 119 165
rect 104 159 109 162
rect 147 159 152 166
rect 154 159 159 179
rect 161 173 168 179
rect 161 163 170 173
rect 161 161 164 163
rect 166 161 170 163
rect 161 159 170 161
rect 172 170 179 173
rect 206 172 211 179
rect 172 168 175 170
rect 177 168 179 170
rect 172 166 179 168
rect 184 170 191 172
rect 184 168 186 170
rect 188 168 191 170
rect 184 166 191 168
rect 172 159 177 166
rect 186 159 191 166
rect 193 166 201 172
rect 193 164 196 166
rect 198 164 201 166
rect 193 162 201 164
rect 203 169 211 172
rect 203 167 206 169
rect 208 167 211 169
rect 203 165 211 167
rect 213 177 221 179
rect 213 175 216 177
rect 218 175 221 177
rect 213 165 221 175
rect 223 177 230 179
rect 223 175 226 177
rect 228 175 230 177
rect 223 170 230 175
rect 236 172 241 179
rect 223 168 226 170
rect 228 168 230 170
rect 223 165 230 168
rect 234 170 241 172
rect 234 168 236 170
rect 238 168 241 170
rect 234 166 241 168
rect 203 162 208 165
rect 193 159 198 162
rect 236 159 241 166
rect 243 159 248 179
rect 250 173 257 179
rect 273 177 280 179
rect 273 175 275 177
rect 277 175 280 177
rect 250 163 259 173
rect 250 161 253 163
rect 255 161 259 163
rect 250 159 259 161
rect 261 170 268 173
rect 261 168 264 170
rect 266 168 268 170
rect 261 166 268 168
rect 273 170 280 175
rect 273 168 275 170
rect 277 168 280 170
rect 261 159 266 166
rect 273 165 280 168
rect 282 174 287 179
rect 295 174 300 176
rect 282 170 290 174
rect 282 168 285 170
rect 287 168 290 170
rect 282 166 290 168
rect 292 172 300 174
rect 292 170 295 172
rect 297 170 300 172
rect 292 168 300 170
rect 302 172 309 176
rect 323 172 328 177
rect 302 170 305 172
rect 307 170 309 172
rect 302 168 309 170
rect 321 170 328 172
rect 321 168 323 170
rect 325 168 328 170
rect 292 166 297 168
rect 282 165 287 166
rect 321 166 328 168
rect 330 166 335 177
rect 337 168 348 177
rect 350 174 355 177
rect 350 172 357 174
rect 385 172 390 179
rect 350 170 353 172
rect 355 170 357 172
rect 350 168 357 170
rect 363 170 370 172
rect 363 168 365 170
rect 367 168 370 170
rect 337 166 346 168
rect 339 160 346 166
rect 363 166 370 168
rect 339 158 342 160
rect 344 158 346 160
rect 339 156 346 158
rect 365 159 370 166
rect 372 166 380 172
rect 372 164 375 166
rect 377 164 380 166
rect 372 162 380 164
rect 382 169 390 172
rect 382 167 385 169
rect 387 167 390 169
rect 382 165 390 167
rect 392 177 400 179
rect 392 175 395 177
rect 397 175 400 177
rect 392 165 400 175
rect 402 177 409 179
rect 402 175 405 177
rect 407 175 409 177
rect 402 170 409 175
rect 415 172 420 179
rect 402 168 405 170
rect 407 168 409 170
rect 402 165 409 168
rect 413 170 420 172
rect 413 168 415 170
rect 417 168 420 170
rect 413 166 420 168
rect 382 162 387 165
rect 372 159 377 162
rect 415 159 420 166
rect 422 159 427 179
rect 429 173 436 179
rect 429 163 438 173
rect 429 161 432 163
rect 434 161 438 163
rect 429 159 438 161
rect 440 170 447 173
rect 474 172 479 179
rect 440 168 443 170
rect 445 168 447 170
rect 440 166 447 168
rect 452 170 459 172
rect 452 168 454 170
rect 456 168 459 170
rect 452 166 459 168
rect 440 159 445 166
rect 454 159 459 166
rect 461 166 469 172
rect 461 164 464 166
rect 466 164 469 166
rect 461 162 469 164
rect 471 169 479 172
rect 471 167 474 169
rect 476 167 479 169
rect 471 165 479 167
rect 481 177 489 179
rect 481 175 484 177
rect 486 175 489 177
rect 481 165 489 175
rect 491 177 498 179
rect 491 175 494 177
rect 496 175 498 177
rect 491 170 498 175
rect 504 172 509 179
rect 491 168 494 170
rect 496 168 498 170
rect 491 165 498 168
rect 502 170 509 172
rect 502 168 504 170
rect 506 168 509 170
rect 502 166 509 168
rect 471 162 476 165
rect 461 159 466 162
rect 504 159 509 166
rect 511 159 516 179
rect 518 173 525 179
rect 541 177 548 179
rect 541 175 543 177
rect 545 175 548 177
rect 518 163 527 173
rect 518 161 521 163
rect 523 161 527 163
rect 518 159 527 161
rect 529 170 536 173
rect 529 168 532 170
rect 534 168 536 170
rect 529 166 536 168
rect 541 170 548 175
rect 541 168 543 170
rect 545 168 548 170
rect 529 159 534 166
rect 541 165 548 168
rect 550 174 555 179
rect 563 174 568 176
rect 550 170 558 174
rect 550 168 553 170
rect 555 168 558 170
rect 550 166 558 168
rect 560 172 568 174
rect 560 170 563 172
rect 565 170 568 172
rect 560 168 568 170
rect 570 172 577 176
rect 591 172 596 177
rect 570 170 573 172
rect 575 170 577 172
rect 570 168 577 170
rect 589 170 596 172
rect 589 168 591 170
rect 593 168 596 170
rect 560 166 565 168
rect 550 165 555 166
rect 589 166 596 168
rect 598 166 603 177
rect 605 168 616 177
rect 618 174 623 177
rect 618 172 625 174
rect 652 172 657 179
rect 618 170 621 172
rect 623 170 625 172
rect 618 168 625 170
rect 630 170 637 172
rect 630 168 632 170
rect 634 168 637 170
rect 605 166 614 168
rect 607 160 614 166
rect 630 166 637 168
rect 607 158 610 160
rect 612 158 614 160
rect 607 156 614 158
rect 632 159 637 166
rect 639 166 647 172
rect 639 164 642 166
rect 644 164 647 166
rect 639 162 647 164
rect 649 169 657 172
rect 649 167 652 169
rect 654 167 657 169
rect 649 165 657 167
rect 659 177 667 179
rect 659 175 662 177
rect 664 175 667 177
rect 659 165 667 175
rect 669 177 676 179
rect 669 175 672 177
rect 674 175 676 177
rect 669 170 676 175
rect 682 172 687 179
rect 669 168 672 170
rect 674 168 676 170
rect 669 165 676 168
rect 680 170 687 172
rect 680 168 682 170
rect 684 168 687 170
rect 680 166 687 168
rect 649 162 654 165
rect 639 159 644 162
rect 682 159 687 166
rect 689 159 694 179
rect 696 173 703 179
rect 696 163 705 173
rect 696 161 699 163
rect 701 161 705 163
rect 696 159 705 161
rect 707 170 714 173
rect 741 172 746 179
rect 707 168 710 170
rect 712 168 714 170
rect 707 166 714 168
rect 719 170 726 172
rect 719 168 721 170
rect 723 168 726 170
rect 719 166 726 168
rect 707 159 712 166
rect 721 159 726 166
rect 728 166 736 172
rect 728 164 731 166
rect 733 164 736 166
rect 728 162 736 164
rect 738 169 746 172
rect 738 167 741 169
rect 743 167 746 169
rect 738 165 746 167
rect 748 177 756 179
rect 748 175 751 177
rect 753 175 756 177
rect 748 165 756 175
rect 758 177 765 179
rect 758 175 761 177
rect 763 175 765 177
rect 758 170 765 175
rect 771 172 776 179
rect 758 168 761 170
rect 763 168 765 170
rect 758 165 765 168
rect 769 170 776 172
rect 769 168 771 170
rect 773 168 776 170
rect 769 166 776 168
rect 738 162 743 165
rect 728 159 733 162
rect 771 159 776 166
rect 778 159 783 179
rect 785 173 792 179
rect 808 177 815 179
rect 808 175 810 177
rect 812 175 815 177
rect 785 163 794 173
rect 785 161 788 163
rect 790 161 794 163
rect 785 159 794 161
rect 796 170 803 173
rect 796 168 799 170
rect 801 168 803 170
rect 796 166 803 168
rect 808 170 815 175
rect 808 168 810 170
rect 812 168 815 170
rect 796 159 801 166
rect 808 165 815 168
rect 817 174 822 179
rect 830 174 835 176
rect 817 170 825 174
rect 817 168 820 170
rect 822 168 825 170
rect 817 166 825 168
rect 827 172 835 174
rect 827 170 830 172
rect 832 170 835 172
rect 827 168 835 170
rect 837 172 844 176
rect 837 170 840 172
rect 842 170 844 172
rect 837 168 844 170
rect 827 166 832 168
rect 817 165 822 166
rect 31 148 38 150
rect 31 146 34 148
rect 36 146 38 148
rect 31 140 38 146
rect 71 148 78 150
rect 71 146 74 148
rect 76 146 78 148
rect 13 138 20 140
rect 13 136 15 138
rect 17 136 20 138
rect 13 134 20 136
rect 15 129 20 134
rect 22 129 27 140
rect 29 138 38 140
rect 71 140 78 146
rect 53 138 60 140
rect 29 129 40 138
rect 42 136 49 138
rect 42 134 45 136
rect 47 134 49 136
rect 53 136 55 138
rect 57 136 60 138
rect 53 134 60 136
rect 42 132 49 134
rect 42 129 47 132
rect 55 129 60 134
rect 62 129 67 140
rect 69 138 78 140
rect 97 140 102 147
rect 95 138 102 140
rect 69 129 80 138
rect 82 136 89 138
rect 82 134 85 136
rect 87 134 89 136
rect 95 136 97 138
rect 99 136 102 138
rect 95 134 102 136
rect 104 144 109 147
rect 104 142 112 144
rect 104 140 107 142
rect 109 140 112 142
rect 104 134 112 140
rect 114 141 119 144
rect 114 139 122 141
rect 114 137 117 139
rect 119 137 122 139
rect 114 134 122 137
rect 82 132 89 134
rect 82 129 87 132
rect 117 127 122 134
rect 124 131 132 141
rect 124 129 127 131
rect 129 129 132 131
rect 124 127 132 129
rect 134 138 141 141
rect 147 140 152 147
rect 134 136 137 138
rect 139 136 141 138
rect 134 131 141 136
rect 145 138 152 140
rect 145 136 147 138
rect 149 136 152 138
rect 145 134 152 136
rect 134 129 137 131
rect 139 129 141 131
rect 134 127 141 129
rect 147 127 152 134
rect 154 127 159 147
rect 161 145 170 147
rect 161 143 164 145
rect 166 143 170 145
rect 161 133 170 143
rect 172 140 177 147
rect 186 140 191 147
rect 172 138 179 140
rect 172 136 175 138
rect 177 136 179 138
rect 172 133 179 136
rect 184 138 191 140
rect 184 136 186 138
rect 188 136 191 138
rect 184 134 191 136
rect 193 144 198 147
rect 193 142 201 144
rect 193 140 196 142
rect 198 140 201 142
rect 193 134 201 140
rect 203 141 208 144
rect 203 139 211 141
rect 203 137 206 139
rect 208 137 211 139
rect 203 134 211 137
rect 161 127 168 133
rect 206 127 211 134
rect 213 131 221 141
rect 213 129 216 131
rect 218 129 221 131
rect 213 127 221 129
rect 223 138 230 141
rect 236 140 241 147
rect 223 136 226 138
rect 228 136 230 138
rect 223 131 230 136
rect 234 138 241 140
rect 234 136 236 138
rect 238 136 241 138
rect 234 134 241 136
rect 223 129 226 131
rect 228 129 230 131
rect 223 127 230 129
rect 236 127 241 134
rect 243 127 248 147
rect 250 145 259 147
rect 250 143 253 145
rect 255 143 259 145
rect 250 133 259 143
rect 261 140 266 147
rect 261 138 268 140
rect 261 136 264 138
rect 266 136 268 138
rect 261 133 268 136
rect 273 138 280 141
rect 273 136 275 138
rect 277 136 280 138
rect 250 127 257 133
rect 273 131 280 136
rect 273 129 275 131
rect 277 129 280 131
rect 273 127 280 129
rect 282 140 287 141
rect 339 148 346 150
rect 339 146 342 148
rect 344 146 346 148
rect 282 138 290 140
rect 282 136 285 138
rect 287 136 290 138
rect 282 132 290 136
rect 292 138 297 140
rect 339 140 346 146
rect 321 138 328 140
rect 292 136 300 138
rect 292 134 295 136
rect 297 134 300 136
rect 292 132 300 134
rect 282 127 287 132
rect 295 130 300 132
rect 302 136 309 138
rect 302 134 305 136
rect 307 134 309 136
rect 321 136 323 138
rect 325 136 328 138
rect 321 134 328 136
rect 302 130 309 134
rect 323 129 328 134
rect 330 129 335 140
rect 337 138 346 140
rect 365 140 370 147
rect 363 138 370 140
rect 337 129 348 138
rect 350 136 357 138
rect 350 134 353 136
rect 355 134 357 136
rect 363 136 365 138
rect 367 136 370 138
rect 363 134 370 136
rect 372 144 377 147
rect 372 142 380 144
rect 372 140 375 142
rect 377 140 380 142
rect 372 134 380 140
rect 382 141 387 144
rect 382 139 390 141
rect 382 137 385 139
rect 387 137 390 139
rect 382 134 390 137
rect 350 132 357 134
rect 350 129 355 132
rect 385 127 390 134
rect 392 131 400 141
rect 392 129 395 131
rect 397 129 400 131
rect 392 127 400 129
rect 402 138 409 141
rect 415 140 420 147
rect 402 136 405 138
rect 407 136 409 138
rect 402 131 409 136
rect 413 138 420 140
rect 413 136 415 138
rect 417 136 420 138
rect 413 134 420 136
rect 402 129 405 131
rect 407 129 409 131
rect 402 127 409 129
rect 415 127 420 134
rect 422 127 427 147
rect 429 145 438 147
rect 429 143 432 145
rect 434 143 438 145
rect 429 133 438 143
rect 440 140 445 147
rect 454 140 459 147
rect 440 138 447 140
rect 440 136 443 138
rect 445 136 447 138
rect 440 133 447 136
rect 452 138 459 140
rect 452 136 454 138
rect 456 136 459 138
rect 452 134 459 136
rect 461 144 466 147
rect 461 142 469 144
rect 461 140 464 142
rect 466 140 469 142
rect 461 134 469 140
rect 471 141 476 144
rect 471 139 479 141
rect 471 137 474 139
rect 476 137 479 139
rect 471 134 479 137
rect 429 127 436 133
rect 474 127 479 134
rect 481 131 489 141
rect 481 129 484 131
rect 486 129 489 131
rect 481 127 489 129
rect 491 138 498 141
rect 504 140 509 147
rect 491 136 494 138
rect 496 136 498 138
rect 491 131 498 136
rect 502 138 509 140
rect 502 136 504 138
rect 506 136 509 138
rect 502 134 509 136
rect 491 129 494 131
rect 496 129 498 131
rect 491 127 498 129
rect 504 127 509 134
rect 511 127 516 147
rect 518 145 527 147
rect 518 143 521 145
rect 523 143 527 145
rect 518 133 527 143
rect 529 140 534 147
rect 529 138 536 140
rect 529 136 532 138
rect 534 136 536 138
rect 529 133 536 136
rect 541 138 548 141
rect 541 136 543 138
rect 545 136 548 138
rect 518 127 525 133
rect 541 131 548 136
rect 541 129 543 131
rect 545 129 548 131
rect 541 127 548 129
rect 550 140 555 141
rect 607 148 614 150
rect 607 146 610 148
rect 612 146 614 148
rect 550 138 558 140
rect 550 136 553 138
rect 555 136 558 138
rect 550 132 558 136
rect 560 138 565 140
rect 607 140 614 146
rect 589 138 596 140
rect 560 136 568 138
rect 560 134 563 136
rect 565 134 568 136
rect 560 132 568 134
rect 550 127 555 132
rect 563 130 568 132
rect 570 136 577 138
rect 570 134 573 136
rect 575 134 577 136
rect 589 136 591 138
rect 593 136 596 138
rect 589 134 596 136
rect 570 130 577 134
rect 591 129 596 134
rect 598 129 603 140
rect 605 138 614 140
rect 632 140 637 147
rect 630 138 637 140
rect 605 129 616 138
rect 618 136 625 138
rect 618 134 621 136
rect 623 134 625 136
rect 630 136 632 138
rect 634 136 637 138
rect 630 134 637 136
rect 639 144 644 147
rect 639 142 647 144
rect 639 140 642 142
rect 644 140 647 142
rect 639 134 647 140
rect 649 141 654 144
rect 649 139 657 141
rect 649 137 652 139
rect 654 137 657 139
rect 649 134 657 137
rect 618 132 625 134
rect 618 129 623 132
rect 652 127 657 134
rect 659 131 667 141
rect 659 129 662 131
rect 664 129 667 131
rect 659 127 667 129
rect 669 138 676 141
rect 682 140 687 147
rect 669 136 672 138
rect 674 136 676 138
rect 669 131 676 136
rect 680 138 687 140
rect 680 136 682 138
rect 684 136 687 138
rect 680 134 687 136
rect 669 129 672 131
rect 674 129 676 131
rect 669 127 676 129
rect 682 127 687 134
rect 689 127 694 147
rect 696 145 705 147
rect 696 143 699 145
rect 701 143 705 145
rect 696 133 705 143
rect 707 140 712 147
rect 721 140 726 147
rect 707 138 714 140
rect 707 136 710 138
rect 712 136 714 138
rect 707 133 714 136
rect 719 138 726 140
rect 719 136 721 138
rect 723 136 726 138
rect 719 134 726 136
rect 728 144 733 147
rect 728 142 736 144
rect 728 140 731 142
rect 733 140 736 142
rect 728 134 736 140
rect 738 141 743 144
rect 738 139 746 141
rect 738 137 741 139
rect 743 137 746 139
rect 738 134 746 137
rect 696 127 703 133
rect 741 127 746 134
rect 748 131 756 141
rect 748 129 751 131
rect 753 129 756 131
rect 748 127 756 129
rect 758 138 765 141
rect 771 140 776 147
rect 758 136 761 138
rect 763 136 765 138
rect 758 131 765 136
rect 769 138 776 140
rect 769 136 771 138
rect 773 136 776 138
rect 769 134 776 136
rect 758 129 761 131
rect 763 129 765 131
rect 758 127 765 129
rect 771 127 776 134
rect 778 127 783 147
rect 785 145 794 147
rect 785 143 788 145
rect 790 143 794 145
rect 785 133 794 143
rect 796 140 801 147
rect 796 138 803 140
rect 796 136 799 138
rect 801 136 803 138
rect 796 133 803 136
rect 808 138 815 141
rect 808 136 810 138
rect 812 136 815 138
rect 785 127 792 133
rect 808 131 815 136
rect 808 129 810 131
rect 812 129 815 131
rect 808 127 815 129
rect 817 140 822 141
rect 817 138 825 140
rect 817 136 820 138
rect 822 136 825 138
rect 817 132 825 136
rect 827 138 832 140
rect 827 136 835 138
rect 827 134 830 136
rect 832 134 835 136
rect 827 132 835 134
rect 817 127 822 132
rect 830 130 835 132
rect 837 136 844 138
rect 837 134 840 136
rect 842 134 844 136
rect 837 130 844 134
rect 15 28 20 33
rect 13 26 20 28
rect 13 24 15 26
rect 17 24 20 26
rect 13 22 20 24
rect 22 22 27 33
rect 29 24 40 33
rect 42 30 47 33
rect 42 28 49 30
rect 55 28 60 33
rect 42 26 45 28
rect 47 26 49 28
rect 42 24 49 26
rect 53 26 60 28
rect 53 24 55 26
rect 57 24 60 26
rect 29 22 38 24
rect 31 16 38 22
rect 53 22 60 24
rect 62 22 67 33
rect 69 24 80 33
rect 82 30 87 33
rect 82 28 89 30
rect 117 28 122 35
rect 82 26 85 28
rect 87 26 89 28
rect 82 24 89 26
rect 95 26 102 28
rect 95 24 97 26
rect 99 24 102 26
rect 69 22 78 24
rect 31 14 34 16
rect 36 14 38 16
rect 31 12 38 14
rect 71 16 78 22
rect 95 22 102 24
rect 71 14 74 16
rect 76 14 78 16
rect 71 12 78 14
rect 97 15 102 22
rect 104 22 112 28
rect 104 20 107 22
rect 109 20 112 22
rect 104 18 112 20
rect 114 25 122 28
rect 114 23 117 25
rect 119 23 122 25
rect 114 21 122 23
rect 124 33 132 35
rect 124 31 127 33
rect 129 31 132 33
rect 124 21 132 31
rect 134 33 141 35
rect 134 31 137 33
rect 139 31 141 33
rect 134 26 141 31
rect 147 28 152 35
rect 134 24 137 26
rect 139 24 141 26
rect 134 21 141 24
rect 145 26 152 28
rect 145 24 147 26
rect 149 24 152 26
rect 145 22 152 24
rect 114 18 119 21
rect 104 15 109 18
rect 147 15 152 22
rect 154 15 159 35
rect 161 29 168 35
rect 161 19 170 29
rect 161 17 164 19
rect 166 17 170 19
rect 161 15 170 17
rect 172 26 179 29
rect 206 28 211 35
rect 172 24 175 26
rect 177 24 179 26
rect 172 22 179 24
rect 184 26 191 28
rect 184 24 186 26
rect 188 24 191 26
rect 184 22 191 24
rect 172 15 177 22
rect 186 15 191 22
rect 193 22 201 28
rect 193 20 196 22
rect 198 20 201 22
rect 193 18 201 20
rect 203 25 211 28
rect 203 23 206 25
rect 208 23 211 25
rect 203 21 211 23
rect 213 33 221 35
rect 213 31 216 33
rect 218 31 221 33
rect 213 21 221 31
rect 223 33 230 35
rect 223 31 226 33
rect 228 31 230 33
rect 223 26 230 31
rect 236 28 241 35
rect 223 24 226 26
rect 228 24 230 26
rect 223 21 230 24
rect 234 26 241 28
rect 234 24 236 26
rect 238 24 241 26
rect 234 22 241 24
rect 203 18 208 21
rect 193 15 198 18
rect 236 15 241 22
rect 243 15 248 35
rect 250 29 257 35
rect 273 33 280 35
rect 273 31 275 33
rect 277 31 280 33
rect 250 19 259 29
rect 250 17 253 19
rect 255 17 259 19
rect 250 15 259 17
rect 261 26 268 29
rect 261 24 264 26
rect 266 24 268 26
rect 261 22 268 24
rect 273 26 280 31
rect 273 24 275 26
rect 277 24 280 26
rect 261 15 266 22
rect 273 21 280 24
rect 282 30 287 35
rect 295 30 300 32
rect 282 26 290 30
rect 282 24 285 26
rect 287 24 290 26
rect 282 22 290 24
rect 292 28 300 30
rect 292 26 295 28
rect 297 26 300 28
rect 292 24 300 26
rect 302 28 309 32
rect 323 28 328 33
rect 302 26 305 28
rect 307 26 309 28
rect 302 24 309 26
rect 321 26 328 28
rect 321 24 323 26
rect 325 24 328 26
rect 292 22 297 24
rect 282 21 287 22
rect 321 22 328 24
rect 330 22 335 33
rect 337 24 348 33
rect 350 30 355 33
rect 350 28 357 30
rect 385 28 390 35
rect 350 26 353 28
rect 355 26 357 28
rect 350 24 357 26
rect 363 26 370 28
rect 363 24 365 26
rect 367 24 370 26
rect 337 22 346 24
rect 339 16 346 22
rect 363 22 370 24
rect 339 14 342 16
rect 344 14 346 16
rect 339 12 346 14
rect 365 15 370 22
rect 372 22 380 28
rect 372 20 375 22
rect 377 20 380 22
rect 372 18 380 20
rect 382 25 390 28
rect 382 23 385 25
rect 387 23 390 25
rect 382 21 390 23
rect 392 33 400 35
rect 392 31 395 33
rect 397 31 400 33
rect 392 21 400 31
rect 402 33 409 35
rect 402 31 405 33
rect 407 31 409 33
rect 402 26 409 31
rect 415 28 420 35
rect 402 24 405 26
rect 407 24 409 26
rect 402 21 409 24
rect 413 26 420 28
rect 413 24 415 26
rect 417 24 420 26
rect 413 22 420 24
rect 382 18 387 21
rect 372 15 377 18
rect 415 15 420 22
rect 422 15 427 35
rect 429 29 436 35
rect 429 19 438 29
rect 429 17 432 19
rect 434 17 438 19
rect 429 15 438 17
rect 440 26 447 29
rect 474 28 479 35
rect 440 24 443 26
rect 445 24 447 26
rect 440 22 447 24
rect 452 26 459 28
rect 452 24 454 26
rect 456 24 459 26
rect 452 22 459 24
rect 440 15 445 22
rect 454 15 459 22
rect 461 22 469 28
rect 461 20 464 22
rect 466 20 469 22
rect 461 18 469 20
rect 471 25 479 28
rect 471 23 474 25
rect 476 23 479 25
rect 471 21 479 23
rect 481 33 489 35
rect 481 31 484 33
rect 486 31 489 33
rect 481 21 489 31
rect 491 33 498 35
rect 491 31 494 33
rect 496 31 498 33
rect 491 26 498 31
rect 504 28 509 35
rect 491 24 494 26
rect 496 24 498 26
rect 491 21 498 24
rect 502 26 509 28
rect 502 24 504 26
rect 506 24 509 26
rect 502 22 509 24
rect 471 18 476 21
rect 461 15 466 18
rect 504 15 509 22
rect 511 15 516 35
rect 518 29 525 35
rect 541 33 548 35
rect 541 31 543 33
rect 545 31 548 33
rect 518 19 527 29
rect 518 17 521 19
rect 523 17 527 19
rect 518 15 527 17
rect 529 26 536 29
rect 529 24 532 26
rect 534 24 536 26
rect 529 22 536 24
rect 541 26 548 31
rect 541 24 543 26
rect 545 24 548 26
rect 529 15 534 22
rect 541 21 548 24
rect 550 30 555 35
rect 563 30 568 32
rect 550 26 558 30
rect 550 24 553 26
rect 555 24 558 26
rect 550 22 558 24
rect 560 28 568 30
rect 560 26 563 28
rect 565 26 568 28
rect 560 24 568 26
rect 570 28 577 32
rect 591 28 596 33
rect 570 26 573 28
rect 575 26 577 28
rect 570 24 577 26
rect 589 26 596 28
rect 589 24 591 26
rect 593 24 596 26
rect 560 22 565 24
rect 550 21 555 22
rect 589 22 596 24
rect 598 22 603 33
rect 605 24 616 33
rect 618 30 623 33
rect 618 28 625 30
rect 652 28 657 35
rect 618 26 621 28
rect 623 26 625 28
rect 618 24 625 26
rect 630 26 637 28
rect 630 24 632 26
rect 634 24 637 26
rect 605 22 614 24
rect 607 16 614 22
rect 630 22 637 24
rect 607 14 610 16
rect 612 14 614 16
rect 607 12 614 14
rect 632 15 637 22
rect 639 22 647 28
rect 639 20 642 22
rect 644 20 647 22
rect 639 18 647 20
rect 649 25 657 28
rect 649 23 652 25
rect 654 23 657 25
rect 649 21 657 23
rect 659 33 667 35
rect 659 31 662 33
rect 664 31 667 33
rect 659 21 667 31
rect 669 33 676 35
rect 669 31 672 33
rect 674 31 676 33
rect 669 26 676 31
rect 682 28 687 35
rect 669 24 672 26
rect 674 24 676 26
rect 669 21 676 24
rect 680 26 687 28
rect 680 24 682 26
rect 684 24 687 26
rect 680 22 687 24
rect 649 18 654 21
rect 639 15 644 18
rect 682 15 687 22
rect 689 15 694 35
rect 696 29 703 35
rect 696 19 705 29
rect 696 17 699 19
rect 701 17 705 19
rect 696 15 705 17
rect 707 26 714 29
rect 741 28 746 35
rect 707 24 710 26
rect 712 24 714 26
rect 707 22 714 24
rect 719 26 726 28
rect 719 24 721 26
rect 723 24 726 26
rect 719 22 726 24
rect 707 15 712 22
rect 721 15 726 22
rect 728 22 736 28
rect 728 20 731 22
rect 733 20 736 22
rect 728 18 736 20
rect 738 25 746 28
rect 738 23 741 25
rect 743 23 746 25
rect 738 21 746 23
rect 748 33 756 35
rect 748 31 751 33
rect 753 31 756 33
rect 748 21 756 31
rect 758 33 765 35
rect 758 31 761 33
rect 763 31 765 33
rect 758 26 765 31
rect 771 28 776 35
rect 758 24 761 26
rect 763 24 765 26
rect 758 21 765 24
rect 769 26 776 28
rect 769 24 771 26
rect 773 24 776 26
rect 769 22 776 24
rect 738 18 743 21
rect 728 15 733 18
rect 771 15 776 22
rect 778 15 783 35
rect 785 29 792 35
rect 808 33 815 35
rect 808 31 810 33
rect 812 31 815 33
rect 785 19 794 29
rect 785 17 788 19
rect 790 17 794 19
rect 785 15 794 17
rect 796 26 803 29
rect 796 24 799 26
rect 801 24 803 26
rect 796 22 803 24
rect 808 26 815 31
rect 808 24 810 26
rect 812 24 815 26
rect 796 15 801 22
rect 808 21 815 24
rect 817 30 822 35
rect 830 30 835 32
rect 817 26 825 30
rect 817 24 820 26
rect 822 24 825 26
rect 817 22 825 24
rect 827 28 835 30
rect 827 26 830 28
rect 832 26 835 28
rect 827 24 835 26
rect 837 28 844 32
rect 837 26 840 28
rect 842 26 844 28
rect 837 24 844 26
rect 827 22 832 24
rect 817 21 822 22
<< pdif >>
rect 34 251 40 258
rect 13 242 20 251
rect 13 240 15 242
rect 17 240 20 242
rect 13 238 20 240
rect 22 249 30 251
rect 22 247 25 249
rect 27 247 30 249
rect 22 242 30 247
rect 22 240 25 242
rect 27 240 30 242
rect 22 238 30 240
rect 32 244 40 251
rect 32 242 35 244
rect 37 242 40 244
rect 32 240 40 242
rect 42 256 49 258
rect 42 254 45 256
rect 47 254 49 256
rect 42 249 49 254
rect 74 251 80 258
rect 42 247 45 249
rect 47 247 49 249
rect 42 245 49 247
rect 42 240 47 245
rect 53 242 60 251
rect 53 240 55 242
rect 57 240 60 242
rect 32 238 38 240
rect 53 238 60 240
rect 62 249 70 251
rect 62 247 65 249
rect 67 247 70 249
rect 62 242 70 247
rect 62 240 65 242
rect 67 240 70 242
rect 62 238 70 240
rect 72 244 80 251
rect 72 242 75 244
rect 77 242 80 244
rect 72 240 80 242
rect 82 256 89 258
rect 120 256 125 259
rect 82 254 85 256
rect 87 254 89 256
rect 82 249 89 254
rect 82 247 85 249
rect 87 247 89 249
rect 82 245 89 247
rect 95 254 102 256
rect 95 252 97 254
rect 99 252 102 254
rect 95 247 102 252
rect 95 245 97 247
rect 99 245 102 247
rect 82 240 87 245
rect 95 243 102 245
rect 72 238 78 240
rect 97 231 102 243
rect 104 243 115 256
rect 117 254 125 256
rect 117 252 120 254
rect 122 252 125 254
rect 117 243 125 252
rect 104 235 113 243
rect 104 233 108 235
rect 110 233 113 235
rect 120 234 125 243
rect 127 234 132 259
rect 134 242 150 259
rect 134 240 143 242
rect 145 240 150 242
rect 134 235 150 240
rect 134 234 143 235
rect 104 231 113 233
rect 136 233 143 234
rect 145 233 150 235
rect 136 231 150 233
rect 152 250 160 259
rect 152 248 155 250
rect 157 248 160 250
rect 152 243 160 248
rect 152 241 155 243
rect 157 241 160 243
rect 152 231 160 241
rect 162 242 170 259
rect 162 240 165 242
rect 167 240 170 242
rect 162 235 170 240
rect 162 233 165 235
rect 167 233 170 235
rect 162 231 170 233
rect 172 257 179 259
rect 172 255 175 257
rect 177 255 179 257
rect 209 256 214 259
rect 172 250 179 255
rect 172 248 175 250
rect 177 248 179 250
rect 172 246 179 248
rect 184 254 191 256
rect 184 252 186 254
rect 188 252 191 254
rect 184 247 191 252
rect 172 231 177 246
rect 184 245 186 247
rect 188 245 191 247
rect 184 243 191 245
rect 186 231 191 243
rect 193 243 204 256
rect 206 254 214 256
rect 206 252 209 254
rect 211 252 214 254
rect 206 243 214 252
rect 193 235 202 243
rect 193 233 197 235
rect 199 233 202 235
rect 209 234 214 243
rect 216 234 221 259
rect 223 242 239 259
rect 223 240 232 242
rect 234 240 239 242
rect 223 235 239 240
rect 223 234 232 235
rect 193 231 202 233
rect 225 233 232 234
rect 234 233 239 235
rect 225 231 239 233
rect 241 250 249 259
rect 241 248 244 250
rect 246 248 249 250
rect 241 243 249 248
rect 241 241 244 243
rect 246 241 249 243
rect 241 231 249 241
rect 251 242 259 259
rect 251 240 254 242
rect 256 240 259 242
rect 251 235 259 240
rect 251 233 254 235
rect 256 233 259 235
rect 251 231 259 233
rect 261 257 268 259
rect 261 255 264 257
rect 266 255 268 257
rect 261 250 268 255
rect 275 250 280 259
rect 261 248 264 250
rect 266 248 268 250
rect 261 246 268 248
rect 273 248 280 250
rect 273 246 275 248
rect 277 246 280 248
rect 261 231 266 246
rect 273 241 280 246
rect 273 239 275 241
rect 277 239 280 241
rect 273 237 280 239
rect 275 231 280 237
rect 282 232 293 259
rect 282 231 286 232
rect 284 230 286 231
rect 288 231 293 232
rect 295 231 300 259
rect 302 243 307 259
rect 342 251 348 258
rect 302 241 309 243
rect 302 239 305 241
rect 307 239 309 241
rect 302 237 309 239
rect 321 242 328 251
rect 321 240 323 242
rect 325 240 328 242
rect 321 238 328 240
rect 330 249 338 251
rect 330 247 333 249
rect 335 247 338 249
rect 330 242 338 247
rect 330 240 333 242
rect 335 240 338 242
rect 330 238 338 240
rect 340 244 348 251
rect 340 242 343 244
rect 345 242 348 244
rect 340 240 348 242
rect 350 256 357 258
rect 388 256 393 259
rect 350 254 353 256
rect 355 254 357 256
rect 350 249 357 254
rect 350 247 353 249
rect 355 247 357 249
rect 350 245 357 247
rect 363 254 370 256
rect 363 252 365 254
rect 367 252 370 254
rect 363 247 370 252
rect 363 245 365 247
rect 367 245 370 247
rect 350 240 355 245
rect 363 243 370 245
rect 340 238 346 240
rect 302 231 307 237
rect 288 230 291 231
rect 284 228 291 230
rect 365 231 370 243
rect 372 243 383 256
rect 385 254 393 256
rect 385 252 388 254
rect 390 252 393 254
rect 385 243 393 252
rect 372 235 381 243
rect 372 233 376 235
rect 378 233 381 235
rect 388 234 393 243
rect 395 234 400 259
rect 402 242 418 259
rect 402 240 411 242
rect 413 240 418 242
rect 402 235 418 240
rect 402 234 411 235
rect 372 231 381 233
rect 404 233 411 234
rect 413 233 418 235
rect 404 231 418 233
rect 420 250 428 259
rect 420 248 423 250
rect 425 248 428 250
rect 420 243 428 248
rect 420 241 423 243
rect 425 241 428 243
rect 420 231 428 241
rect 430 242 438 259
rect 430 240 433 242
rect 435 240 438 242
rect 430 235 438 240
rect 430 233 433 235
rect 435 233 438 235
rect 430 231 438 233
rect 440 257 447 259
rect 440 255 443 257
rect 445 255 447 257
rect 477 256 482 259
rect 440 250 447 255
rect 440 248 443 250
rect 445 248 447 250
rect 440 246 447 248
rect 452 254 459 256
rect 452 252 454 254
rect 456 252 459 254
rect 452 247 459 252
rect 440 231 445 246
rect 452 245 454 247
rect 456 245 459 247
rect 452 243 459 245
rect 454 231 459 243
rect 461 243 472 256
rect 474 254 482 256
rect 474 252 477 254
rect 479 252 482 254
rect 474 243 482 252
rect 461 235 470 243
rect 461 233 465 235
rect 467 233 470 235
rect 477 234 482 243
rect 484 234 489 259
rect 491 242 507 259
rect 491 240 500 242
rect 502 240 507 242
rect 491 235 507 240
rect 491 234 500 235
rect 461 231 470 233
rect 493 233 500 234
rect 502 233 507 235
rect 493 231 507 233
rect 509 250 517 259
rect 509 248 512 250
rect 514 248 517 250
rect 509 243 517 248
rect 509 241 512 243
rect 514 241 517 243
rect 509 231 517 241
rect 519 242 527 259
rect 519 240 522 242
rect 524 240 527 242
rect 519 235 527 240
rect 519 233 522 235
rect 524 233 527 235
rect 519 231 527 233
rect 529 257 536 259
rect 529 255 532 257
rect 534 255 536 257
rect 529 250 536 255
rect 543 250 548 259
rect 529 248 532 250
rect 534 248 536 250
rect 529 246 536 248
rect 541 248 548 250
rect 541 246 543 248
rect 545 246 548 248
rect 529 231 534 246
rect 541 241 548 246
rect 541 239 543 241
rect 545 239 548 241
rect 541 237 548 239
rect 543 231 548 237
rect 550 232 561 259
rect 550 231 554 232
rect 552 230 554 231
rect 556 231 561 232
rect 563 231 568 259
rect 570 243 575 259
rect 610 251 616 258
rect 570 241 577 243
rect 570 239 573 241
rect 575 239 577 241
rect 570 237 577 239
rect 589 242 596 251
rect 589 240 591 242
rect 593 240 596 242
rect 589 238 596 240
rect 598 249 606 251
rect 598 247 601 249
rect 603 247 606 249
rect 598 242 606 247
rect 598 240 601 242
rect 603 240 606 242
rect 598 238 606 240
rect 608 244 616 251
rect 608 242 611 244
rect 613 242 616 244
rect 608 240 616 242
rect 618 256 625 258
rect 655 256 660 259
rect 618 254 621 256
rect 623 254 625 256
rect 618 249 625 254
rect 618 247 621 249
rect 623 247 625 249
rect 618 245 625 247
rect 630 254 637 256
rect 630 252 632 254
rect 634 252 637 254
rect 630 247 637 252
rect 630 245 632 247
rect 634 245 637 247
rect 618 240 623 245
rect 630 243 637 245
rect 608 238 614 240
rect 570 231 575 237
rect 556 230 559 231
rect 552 228 559 230
rect 632 231 637 243
rect 639 243 650 256
rect 652 254 660 256
rect 652 252 655 254
rect 657 252 660 254
rect 652 243 660 252
rect 639 235 648 243
rect 639 233 643 235
rect 645 233 648 235
rect 655 234 660 243
rect 662 234 667 259
rect 669 242 685 259
rect 669 240 678 242
rect 680 240 685 242
rect 669 235 685 240
rect 669 234 678 235
rect 639 231 648 233
rect 671 233 678 234
rect 680 233 685 235
rect 671 231 685 233
rect 687 250 695 259
rect 687 248 690 250
rect 692 248 695 250
rect 687 243 695 248
rect 687 241 690 243
rect 692 241 695 243
rect 687 231 695 241
rect 697 242 705 259
rect 697 240 700 242
rect 702 240 705 242
rect 697 235 705 240
rect 697 233 700 235
rect 702 233 705 235
rect 697 231 705 233
rect 707 257 714 259
rect 707 255 710 257
rect 712 255 714 257
rect 744 256 749 259
rect 707 250 714 255
rect 707 248 710 250
rect 712 248 714 250
rect 707 246 714 248
rect 719 254 726 256
rect 719 252 721 254
rect 723 252 726 254
rect 719 247 726 252
rect 707 231 712 246
rect 719 245 721 247
rect 723 245 726 247
rect 719 243 726 245
rect 721 231 726 243
rect 728 243 739 256
rect 741 254 749 256
rect 741 252 744 254
rect 746 252 749 254
rect 741 243 749 252
rect 728 235 737 243
rect 728 233 732 235
rect 734 233 737 235
rect 744 234 749 243
rect 751 234 756 259
rect 758 242 774 259
rect 758 240 767 242
rect 769 240 774 242
rect 758 235 774 240
rect 758 234 767 235
rect 728 231 737 233
rect 760 233 767 234
rect 769 233 774 235
rect 760 231 774 233
rect 776 250 784 259
rect 776 248 779 250
rect 781 248 784 250
rect 776 243 784 248
rect 776 241 779 243
rect 781 241 784 243
rect 776 231 784 241
rect 786 242 794 259
rect 786 240 789 242
rect 791 240 794 242
rect 786 235 794 240
rect 786 233 789 235
rect 791 233 794 235
rect 786 231 794 233
rect 796 257 803 259
rect 796 255 799 257
rect 801 255 803 257
rect 796 250 803 255
rect 810 250 815 259
rect 796 248 799 250
rect 801 248 803 250
rect 796 246 803 248
rect 808 248 815 250
rect 808 246 810 248
rect 812 246 815 248
rect 796 231 801 246
rect 808 241 815 246
rect 808 239 810 241
rect 812 239 815 241
rect 808 237 815 239
rect 810 231 815 237
rect 817 232 828 259
rect 817 231 821 232
rect 819 230 821 231
rect 823 231 828 232
rect 830 231 835 259
rect 837 243 842 259
rect 837 241 844 243
rect 837 239 840 241
rect 842 239 844 241
rect 837 237 844 239
rect 837 231 842 237
rect 823 230 826 231
rect 819 228 826 230
rect 13 210 20 212
rect 13 208 15 210
rect 17 208 20 210
rect 13 199 20 208
rect 22 210 30 212
rect 22 208 25 210
rect 27 208 30 210
rect 22 203 30 208
rect 22 201 25 203
rect 27 201 30 203
rect 22 199 30 201
rect 32 210 38 212
rect 53 210 60 212
rect 32 208 40 210
rect 32 206 35 208
rect 37 206 40 208
rect 32 199 40 206
rect 34 192 40 199
rect 42 205 47 210
rect 53 208 55 210
rect 57 208 60 210
rect 42 203 49 205
rect 42 201 45 203
rect 47 201 49 203
rect 42 196 49 201
rect 53 199 60 208
rect 62 210 70 212
rect 62 208 65 210
rect 67 208 70 210
rect 62 203 70 208
rect 62 201 65 203
rect 67 201 70 203
rect 62 199 70 201
rect 72 210 78 212
rect 72 208 80 210
rect 72 206 75 208
rect 77 206 80 208
rect 72 199 80 206
rect 42 194 45 196
rect 47 194 49 196
rect 42 192 49 194
rect 74 192 80 199
rect 82 205 87 210
rect 97 207 102 219
rect 95 205 102 207
rect 82 203 89 205
rect 82 201 85 203
rect 87 201 89 203
rect 82 196 89 201
rect 82 194 85 196
rect 87 194 89 196
rect 95 203 97 205
rect 99 203 102 205
rect 95 198 102 203
rect 95 196 97 198
rect 99 196 102 198
rect 95 194 102 196
rect 104 217 113 219
rect 104 215 108 217
rect 110 215 113 217
rect 136 217 150 219
rect 136 216 143 217
rect 104 207 113 215
rect 120 207 125 216
rect 104 194 115 207
rect 117 198 125 207
rect 117 196 120 198
rect 122 196 125 198
rect 117 194 125 196
rect 82 192 89 194
rect 120 191 125 194
rect 127 191 132 216
rect 134 215 143 216
rect 145 215 150 217
rect 134 210 150 215
rect 134 208 143 210
rect 145 208 150 210
rect 134 191 150 208
rect 152 209 160 219
rect 152 207 155 209
rect 157 207 160 209
rect 152 202 160 207
rect 152 200 155 202
rect 157 200 160 202
rect 152 191 160 200
rect 162 217 170 219
rect 162 215 165 217
rect 167 215 170 217
rect 162 210 170 215
rect 162 208 165 210
rect 167 208 170 210
rect 162 191 170 208
rect 172 204 177 219
rect 186 207 191 219
rect 184 205 191 207
rect 172 202 179 204
rect 172 200 175 202
rect 177 200 179 202
rect 172 195 179 200
rect 172 193 175 195
rect 177 193 179 195
rect 184 203 186 205
rect 188 203 191 205
rect 184 198 191 203
rect 184 196 186 198
rect 188 196 191 198
rect 184 194 191 196
rect 193 217 202 219
rect 193 215 197 217
rect 199 215 202 217
rect 284 220 291 222
rect 284 219 286 220
rect 225 217 239 219
rect 225 216 232 217
rect 193 207 202 215
rect 209 207 214 216
rect 193 194 204 207
rect 206 198 214 207
rect 206 196 209 198
rect 211 196 214 198
rect 206 194 214 196
rect 172 191 179 193
rect 209 191 214 194
rect 216 191 221 216
rect 223 215 232 216
rect 234 215 239 217
rect 223 210 239 215
rect 223 208 232 210
rect 234 208 239 210
rect 223 191 239 208
rect 241 209 249 219
rect 241 207 244 209
rect 246 207 249 209
rect 241 202 249 207
rect 241 200 244 202
rect 246 200 249 202
rect 241 191 249 200
rect 251 217 259 219
rect 251 215 254 217
rect 256 215 259 217
rect 251 210 259 215
rect 251 208 254 210
rect 256 208 259 210
rect 251 191 259 208
rect 261 204 266 219
rect 275 213 280 219
rect 273 211 280 213
rect 273 209 275 211
rect 277 209 280 211
rect 273 204 280 209
rect 261 202 268 204
rect 261 200 264 202
rect 266 200 268 202
rect 273 202 275 204
rect 277 202 280 204
rect 273 200 280 202
rect 261 195 268 200
rect 261 193 264 195
rect 266 193 268 195
rect 261 191 268 193
rect 275 191 280 200
rect 282 218 286 219
rect 288 219 291 220
rect 288 218 293 219
rect 282 191 293 218
rect 295 191 300 219
rect 302 213 307 219
rect 302 211 309 213
rect 302 209 305 211
rect 307 209 309 211
rect 302 207 309 209
rect 321 210 328 212
rect 321 208 323 210
rect 325 208 328 210
rect 302 191 307 207
rect 321 199 328 208
rect 330 210 338 212
rect 330 208 333 210
rect 335 208 338 210
rect 330 203 338 208
rect 330 201 333 203
rect 335 201 338 203
rect 330 199 338 201
rect 340 210 346 212
rect 340 208 348 210
rect 340 206 343 208
rect 345 206 348 208
rect 340 199 348 206
rect 342 192 348 199
rect 350 205 355 210
rect 365 207 370 219
rect 363 205 370 207
rect 350 203 357 205
rect 350 201 353 203
rect 355 201 357 203
rect 350 196 357 201
rect 350 194 353 196
rect 355 194 357 196
rect 363 203 365 205
rect 367 203 370 205
rect 363 198 370 203
rect 363 196 365 198
rect 367 196 370 198
rect 363 194 370 196
rect 372 217 381 219
rect 372 215 376 217
rect 378 215 381 217
rect 404 217 418 219
rect 404 216 411 217
rect 372 207 381 215
rect 388 207 393 216
rect 372 194 383 207
rect 385 198 393 207
rect 385 196 388 198
rect 390 196 393 198
rect 385 194 393 196
rect 350 192 357 194
rect 388 191 393 194
rect 395 191 400 216
rect 402 215 411 216
rect 413 215 418 217
rect 402 210 418 215
rect 402 208 411 210
rect 413 208 418 210
rect 402 191 418 208
rect 420 209 428 219
rect 420 207 423 209
rect 425 207 428 209
rect 420 202 428 207
rect 420 200 423 202
rect 425 200 428 202
rect 420 191 428 200
rect 430 217 438 219
rect 430 215 433 217
rect 435 215 438 217
rect 430 210 438 215
rect 430 208 433 210
rect 435 208 438 210
rect 430 191 438 208
rect 440 204 445 219
rect 454 207 459 219
rect 452 205 459 207
rect 440 202 447 204
rect 440 200 443 202
rect 445 200 447 202
rect 440 195 447 200
rect 440 193 443 195
rect 445 193 447 195
rect 452 203 454 205
rect 456 203 459 205
rect 452 198 459 203
rect 452 196 454 198
rect 456 196 459 198
rect 452 194 459 196
rect 461 217 470 219
rect 461 215 465 217
rect 467 215 470 217
rect 552 220 559 222
rect 552 219 554 220
rect 493 217 507 219
rect 493 216 500 217
rect 461 207 470 215
rect 477 207 482 216
rect 461 194 472 207
rect 474 198 482 207
rect 474 196 477 198
rect 479 196 482 198
rect 474 194 482 196
rect 440 191 447 193
rect 477 191 482 194
rect 484 191 489 216
rect 491 215 500 216
rect 502 215 507 217
rect 491 210 507 215
rect 491 208 500 210
rect 502 208 507 210
rect 491 191 507 208
rect 509 209 517 219
rect 509 207 512 209
rect 514 207 517 209
rect 509 202 517 207
rect 509 200 512 202
rect 514 200 517 202
rect 509 191 517 200
rect 519 217 527 219
rect 519 215 522 217
rect 524 215 527 217
rect 519 210 527 215
rect 519 208 522 210
rect 524 208 527 210
rect 519 191 527 208
rect 529 204 534 219
rect 543 213 548 219
rect 541 211 548 213
rect 541 209 543 211
rect 545 209 548 211
rect 541 204 548 209
rect 529 202 536 204
rect 529 200 532 202
rect 534 200 536 202
rect 541 202 543 204
rect 545 202 548 204
rect 541 200 548 202
rect 529 195 536 200
rect 529 193 532 195
rect 534 193 536 195
rect 529 191 536 193
rect 543 191 548 200
rect 550 218 554 219
rect 556 219 559 220
rect 556 218 561 219
rect 550 191 561 218
rect 563 191 568 219
rect 570 213 575 219
rect 570 211 577 213
rect 570 209 573 211
rect 575 209 577 211
rect 570 207 577 209
rect 589 210 596 212
rect 589 208 591 210
rect 593 208 596 210
rect 570 191 575 207
rect 589 199 596 208
rect 598 210 606 212
rect 598 208 601 210
rect 603 208 606 210
rect 598 203 606 208
rect 598 201 601 203
rect 603 201 606 203
rect 598 199 606 201
rect 608 210 614 212
rect 608 208 616 210
rect 608 206 611 208
rect 613 206 616 208
rect 608 199 616 206
rect 610 192 616 199
rect 618 205 623 210
rect 632 207 637 219
rect 630 205 637 207
rect 618 203 625 205
rect 618 201 621 203
rect 623 201 625 203
rect 618 196 625 201
rect 618 194 621 196
rect 623 194 625 196
rect 630 203 632 205
rect 634 203 637 205
rect 630 198 637 203
rect 630 196 632 198
rect 634 196 637 198
rect 630 194 637 196
rect 639 217 648 219
rect 639 215 643 217
rect 645 215 648 217
rect 671 217 685 219
rect 671 216 678 217
rect 639 207 648 215
rect 655 207 660 216
rect 639 194 650 207
rect 652 198 660 207
rect 652 196 655 198
rect 657 196 660 198
rect 652 194 660 196
rect 618 192 625 194
rect 655 191 660 194
rect 662 191 667 216
rect 669 215 678 216
rect 680 215 685 217
rect 669 210 685 215
rect 669 208 678 210
rect 680 208 685 210
rect 669 191 685 208
rect 687 209 695 219
rect 687 207 690 209
rect 692 207 695 209
rect 687 202 695 207
rect 687 200 690 202
rect 692 200 695 202
rect 687 191 695 200
rect 697 217 705 219
rect 697 215 700 217
rect 702 215 705 217
rect 697 210 705 215
rect 697 208 700 210
rect 702 208 705 210
rect 697 191 705 208
rect 707 204 712 219
rect 721 207 726 219
rect 719 205 726 207
rect 707 202 714 204
rect 707 200 710 202
rect 712 200 714 202
rect 707 195 714 200
rect 707 193 710 195
rect 712 193 714 195
rect 719 203 721 205
rect 723 203 726 205
rect 719 198 726 203
rect 719 196 721 198
rect 723 196 726 198
rect 719 194 726 196
rect 728 217 737 219
rect 728 215 732 217
rect 734 215 737 217
rect 819 220 826 222
rect 819 219 821 220
rect 760 217 774 219
rect 760 216 767 217
rect 728 207 737 215
rect 744 207 749 216
rect 728 194 739 207
rect 741 198 749 207
rect 741 196 744 198
rect 746 196 749 198
rect 741 194 749 196
rect 707 191 714 193
rect 744 191 749 194
rect 751 191 756 216
rect 758 215 767 216
rect 769 215 774 217
rect 758 210 774 215
rect 758 208 767 210
rect 769 208 774 210
rect 758 191 774 208
rect 776 209 784 219
rect 776 207 779 209
rect 781 207 784 209
rect 776 202 784 207
rect 776 200 779 202
rect 781 200 784 202
rect 776 191 784 200
rect 786 217 794 219
rect 786 215 789 217
rect 791 215 794 217
rect 786 210 794 215
rect 786 208 789 210
rect 791 208 794 210
rect 786 191 794 208
rect 796 204 801 219
rect 810 213 815 219
rect 808 211 815 213
rect 808 209 810 211
rect 812 209 815 211
rect 808 204 815 209
rect 796 202 803 204
rect 796 200 799 202
rect 801 200 803 202
rect 808 202 810 204
rect 812 202 815 204
rect 808 200 815 202
rect 796 195 803 200
rect 796 193 799 195
rect 801 193 803 195
rect 796 191 803 193
rect 810 191 815 200
rect 817 218 821 219
rect 823 219 826 220
rect 823 218 828 219
rect 817 191 828 218
rect 830 191 835 219
rect 837 213 842 219
rect 837 211 844 213
rect 837 209 840 211
rect 842 209 844 211
rect 837 207 844 209
rect 837 191 842 207
rect 34 107 40 114
rect 13 98 20 107
rect 13 96 15 98
rect 17 96 20 98
rect 13 94 20 96
rect 22 105 30 107
rect 22 103 25 105
rect 27 103 30 105
rect 22 98 30 103
rect 22 96 25 98
rect 27 96 30 98
rect 22 94 30 96
rect 32 100 40 107
rect 32 98 35 100
rect 37 98 40 100
rect 32 96 40 98
rect 42 112 49 114
rect 42 110 45 112
rect 47 110 49 112
rect 42 105 49 110
rect 74 107 80 114
rect 42 103 45 105
rect 47 103 49 105
rect 42 101 49 103
rect 42 96 47 101
rect 53 98 60 107
rect 53 96 55 98
rect 57 96 60 98
rect 32 94 38 96
rect 53 94 60 96
rect 62 105 70 107
rect 62 103 65 105
rect 67 103 70 105
rect 62 98 70 103
rect 62 96 65 98
rect 67 96 70 98
rect 62 94 70 96
rect 72 100 80 107
rect 72 98 75 100
rect 77 98 80 100
rect 72 96 80 98
rect 82 112 89 114
rect 120 112 125 115
rect 82 110 85 112
rect 87 110 89 112
rect 82 105 89 110
rect 82 103 85 105
rect 87 103 89 105
rect 82 101 89 103
rect 95 110 102 112
rect 95 108 97 110
rect 99 108 102 110
rect 95 103 102 108
rect 95 101 97 103
rect 99 101 102 103
rect 82 96 87 101
rect 95 99 102 101
rect 72 94 78 96
rect 97 87 102 99
rect 104 99 115 112
rect 117 110 125 112
rect 117 108 120 110
rect 122 108 125 110
rect 117 99 125 108
rect 104 91 113 99
rect 104 89 108 91
rect 110 89 113 91
rect 120 90 125 99
rect 127 90 132 115
rect 134 98 150 115
rect 134 96 143 98
rect 145 96 150 98
rect 134 91 150 96
rect 134 90 143 91
rect 104 87 113 89
rect 136 89 143 90
rect 145 89 150 91
rect 136 87 150 89
rect 152 106 160 115
rect 152 104 155 106
rect 157 104 160 106
rect 152 99 160 104
rect 152 97 155 99
rect 157 97 160 99
rect 152 87 160 97
rect 162 98 170 115
rect 162 96 165 98
rect 167 96 170 98
rect 162 91 170 96
rect 162 89 165 91
rect 167 89 170 91
rect 162 87 170 89
rect 172 113 179 115
rect 172 111 175 113
rect 177 111 179 113
rect 209 112 214 115
rect 172 106 179 111
rect 172 104 175 106
rect 177 104 179 106
rect 172 102 179 104
rect 184 110 191 112
rect 184 108 186 110
rect 188 108 191 110
rect 184 103 191 108
rect 172 87 177 102
rect 184 101 186 103
rect 188 101 191 103
rect 184 99 191 101
rect 186 87 191 99
rect 193 99 204 112
rect 206 110 214 112
rect 206 108 209 110
rect 211 108 214 110
rect 206 99 214 108
rect 193 91 202 99
rect 193 89 197 91
rect 199 89 202 91
rect 209 90 214 99
rect 216 90 221 115
rect 223 98 239 115
rect 223 96 232 98
rect 234 96 239 98
rect 223 91 239 96
rect 223 90 232 91
rect 193 87 202 89
rect 225 89 232 90
rect 234 89 239 91
rect 225 87 239 89
rect 241 106 249 115
rect 241 104 244 106
rect 246 104 249 106
rect 241 99 249 104
rect 241 97 244 99
rect 246 97 249 99
rect 241 87 249 97
rect 251 98 259 115
rect 251 96 254 98
rect 256 96 259 98
rect 251 91 259 96
rect 251 89 254 91
rect 256 89 259 91
rect 251 87 259 89
rect 261 113 268 115
rect 261 111 264 113
rect 266 111 268 113
rect 261 106 268 111
rect 275 106 280 115
rect 261 104 264 106
rect 266 104 268 106
rect 261 102 268 104
rect 273 104 280 106
rect 273 102 275 104
rect 277 102 280 104
rect 261 87 266 102
rect 273 97 280 102
rect 273 95 275 97
rect 277 95 280 97
rect 273 93 280 95
rect 275 87 280 93
rect 282 88 293 115
rect 282 87 286 88
rect 284 86 286 87
rect 288 87 293 88
rect 295 87 300 115
rect 302 99 307 115
rect 342 107 348 114
rect 302 97 309 99
rect 302 95 305 97
rect 307 95 309 97
rect 302 93 309 95
rect 321 98 328 107
rect 321 96 323 98
rect 325 96 328 98
rect 321 94 328 96
rect 330 105 338 107
rect 330 103 333 105
rect 335 103 338 105
rect 330 98 338 103
rect 330 96 333 98
rect 335 96 338 98
rect 330 94 338 96
rect 340 100 348 107
rect 340 98 343 100
rect 345 98 348 100
rect 340 96 348 98
rect 350 112 357 114
rect 388 112 393 115
rect 350 110 353 112
rect 355 110 357 112
rect 350 105 357 110
rect 350 103 353 105
rect 355 103 357 105
rect 350 101 357 103
rect 363 110 370 112
rect 363 108 365 110
rect 367 108 370 110
rect 363 103 370 108
rect 363 101 365 103
rect 367 101 370 103
rect 350 96 355 101
rect 363 99 370 101
rect 340 94 346 96
rect 302 87 307 93
rect 288 86 291 87
rect 284 84 291 86
rect 365 87 370 99
rect 372 99 383 112
rect 385 110 393 112
rect 385 108 388 110
rect 390 108 393 110
rect 385 99 393 108
rect 372 91 381 99
rect 372 89 376 91
rect 378 89 381 91
rect 388 90 393 99
rect 395 90 400 115
rect 402 98 418 115
rect 402 96 411 98
rect 413 96 418 98
rect 402 91 418 96
rect 402 90 411 91
rect 372 87 381 89
rect 404 89 411 90
rect 413 89 418 91
rect 404 87 418 89
rect 420 106 428 115
rect 420 104 423 106
rect 425 104 428 106
rect 420 99 428 104
rect 420 97 423 99
rect 425 97 428 99
rect 420 87 428 97
rect 430 98 438 115
rect 430 96 433 98
rect 435 96 438 98
rect 430 91 438 96
rect 430 89 433 91
rect 435 89 438 91
rect 430 87 438 89
rect 440 113 447 115
rect 440 111 443 113
rect 445 111 447 113
rect 477 112 482 115
rect 440 106 447 111
rect 440 104 443 106
rect 445 104 447 106
rect 440 102 447 104
rect 452 110 459 112
rect 452 108 454 110
rect 456 108 459 110
rect 452 103 459 108
rect 440 87 445 102
rect 452 101 454 103
rect 456 101 459 103
rect 452 99 459 101
rect 454 87 459 99
rect 461 99 472 112
rect 474 110 482 112
rect 474 108 477 110
rect 479 108 482 110
rect 474 99 482 108
rect 461 91 470 99
rect 461 89 465 91
rect 467 89 470 91
rect 477 90 482 99
rect 484 90 489 115
rect 491 98 507 115
rect 491 96 500 98
rect 502 96 507 98
rect 491 91 507 96
rect 491 90 500 91
rect 461 87 470 89
rect 493 89 500 90
rect 502 89 507 91
rect 493 87 507 89
rect 509 106 517 115
rect 509 104 512 106
rect 514 104 517 106
rect 509 99 517 104
rect 509 97 512 99
rect 514 97 517 99
rect 509 87 517 97
rect 519 98 527 115
rect 519 96 522 98
rect 524 96 527 98
rect 519 91 527 96
rect 519 89 522 91
rect 524 89 527 91
rect 519 87 527 89
rect 529 113 536 115
rect 529 111 532 113
rect 534 111 536 113
rect 529 106 536 111
rect 543 106 548 115
rect 529 104 532 106
rect 534 104 536 106
rect 529 102 536 104
rect 541 104 548 106
rect 541 102 543 104
rect 545 102 548 104
rect 529 87 534 102
rect 541 97 548 102
rect 541 95 543 97
rect 545 95 548 97
rect 541 93 548 95
rect 543 87 548 93
rect 550 88 561 115
rect 550 87 554 88
rect 552 86 554 87
rect 556 87 561 88
rect 563 87 568 115
rect 570 99 575 115
rect 610 107 616 114
rect 570 97 577 99
rect 570 95 573 97
rect 575 95 577 97
rect 570 93 577 95
rect 589 98 596 107
rect 589 96 591 98
rect 593 96 596 98
rect 589 94 596 96
rect 598 105 606 107
rect 598 103 601 105
rect 603 103 606 105
rect 598 98 606 103
rect 598 96 601 98
rect 603 96 606 98
rect 598 94 606 96
rect 608 100 616 107
rect 608 98 611 100
rect 613 98 616 100
rect 608 96 616 98
rect 618 112 625 114
rect 655 112 660 115
rect 618 110 621 112
rect 623 110 625 112
rect 618 105 625 110
rect 618 103 621 105
rect 623 103 625 105
rect 618 101 625 103
rect 630 110 637 112
rect 630 108 632 110
rect 634 108 637 110
rect 630 103 637 108
rect 630 101 632 103
rect 634 101 637 103
rect 618 96 623 101
rect 630 99 637 101
rect 608 94 614 96
rect 570 87 575 93
rect 556 86 559 87
rect 552 84 559 86
rect 632 87 637 99
rect 639 99 650 112
rect 652 110 660 112
rect 652 108 655 110
rect 657 108 660 110
rect 652 99 660 108
rect 639 91 648 99
rect 639 89 643 91
rect 645 89 648 91
rect 655 90 660 99
rect 662 90 667 115
rect 669 98 685 115
rect 669 96 678 98
rect 680 96 685 98
rect 669 91 685 96
rect 669 90 678 91
rect 639 87 648 89
rect 671 89 678 90
rect 680 89 685 91
rect 671 87 685 89
rect 687 106 695 115
rect 687 104 690 106
rect 692 104 695 106
rect 687 99 695 104
rect 687 97 690 99
rect 692 97 695 99
rect 687 87 695 97
rect 697 98 705 115
rect 697 96 700 98
rect 702 96 705 98
rect 697 91 705 96
rect 697 89 700 91
rect 702 89 705 91
rect 697 87 705 89
rect 707 113 714 115
rect 707 111 710 113
rect 712 111 714 113
rect 744 112 749 115
rect 707 106 714 111
rect 707 104 710 106
rect 712 104 714 106
rect 707 102 714 104
rect 719 110 726 112
rect 719 108 721 110
rect 723 108 726 110
rect 719 103 726 108
rect 707 87 712 102
rect 719 101 721 103
rect 723 101 726 103
rect 719 99 726 101
rect 721 87 726 99
rect 728 99 739 112
rect 741 110 749 112
rect 741 108 744 110
rect 746 108 749 110
rect 741 99 749 108
rect 728 91 737 99
rect 728 89 732 91
rect 734 89 737 91
rect 744 90 749 99
rect 751 90 756 115
rect 758 98 774 115
rect 758 96 767 98
rect 769 96 774 98
rect 758 91 774 96
rect 758 90 767 91
rect 728 87 737 89
rect 760 89 767 90
rect 769 89 774 91
rect 760 87 774 89
rect 776 106 784 115
rect 776 104 779 106
rect 781 104 784 106
rect 776 99 784 104
rect 776 97 779 99
rect 781 97 784 99
rect 776 87 784 97
rect 786 98 794 115
rect 786 96 789 98
rect 791 96 794 98
rect 786 91 794 96
rect 786 89 789 91
rect 791 89 794 91
rect 786 87 794 89
rect 796 113 803 115
rect 796 111 799 113
rect 801 111 803 113
rect 796 106 803 111
rect 810 106 815 115
rect 796 104 799 106
rect 801 104 803 106
rect 796 102 803 104
rect 808 104 815 106
rect 808 102 810 104
rect 812 102 815 104
rect 796 87 801 102
rect 808 97 815 102
rect 808 95 810 97
rect 812 95 815 97
rect 808 93 815 95
rect 810 87 815 93
rect 817 88 828 115
rect 817 87 821 88
rect 819 86 821 87
rect 823 87 828 88
rect 830 87 835 115
rect 837 99 842 115
rect 837 97 844 99
rect 837 95 840 97
rect 842 95 844 97
rect 837 93 844 95
rect 837 87 842 93
rect 823 86 826 87
rect 819 84 826 86
rect 13 66 20 68
rect 13 64 15 66
rect 17 64 20 66
rect 13 55 20 64
rect 22 66 30 68
rect 22 64 25 66
rect 27 64 30 66
rect 22 59 30 64
rect 22 57 25 59
rect 27 57 30 59
rect 22 55 30 57
rect 32 66 38 68
rect 53 66 60 68
rect 32 64 40 66
rect 32 62 35 64
rect 37 62 40 64
rect 32 55 40 62
rect 34 48 40 55
rect 42 61 47 66
rect 53 64 55 66
rect 57 64 60 66
rect 42 59 49 61
rect 42 57 45 59
rect 47 57 49 59
rect 42 52 49 57
rect 53 55 60 64
rect 62 66 70 68
rect 62 64 65 66
rect 67 64 70 66
rect 62 59 70 64
rect 62 57 65 59
rect 67 57 70 59
rect 62 55 70 57
rect 72 66 78 68
rect 72 64 80 66
rect 72 62 75 64
rect 77 62 80 64
rect 72 55 80 62
rect 42 50 45 52
rect 47 50 49 52
rect 42 48 49 50
rect 74 48 80 55
rect 82 61 87 66
rect 97 63 102 75
rect 95 61 102 63
rect 82 59 89 61
rect 82 57 85 59
rect 87 57 89 59
rect 82 52 89 57
rect 82 50 85 52
rect 87 50 89 52
rect 95 59 97 61
rect 99 59 102 61
rect 95 54 102 59
rect 95 52 97 54
rect 99 52 102 54
rect 95 50 102 52
rect 104 73 113 75
rect 104 71 108 73
rect 110 71 113 73
rect 136 73 150 75
rect 136 72 143 73
rect 104 63 113 71
rect 120 63 125 72
rect 104 50 115 63
rect 117 54 125 63
rect 117 52 120 54
rect 122 52 125 54
rect 117 50 125 52
rect 82 48 89 50
rect 120 47 125 50
rect 127 47 132 72
rect 134 71 143 72
rect 145 71 150 73
rect 134 66 150 71
rect 134 64 143 66
rect 145 64 150 66
rect 134 47 150 64
rect 152 65 160 75
rect 152 63 155 65
rect 157 63 160 65
rect 152 58 160 63
rect 152 56 155 58
rect 157 56 160 58
rect 152 47 160 56
rect 162 73 170 75
rect 162 71 165 73
rect 167 71 170 73
rect 162 66 170 71
rect 162 64 165 66
rect 167 64 170 66
rect 162 47 170 64
rect 172 60 177 75
rect 186 63 191 75
rect 184 61 191 63
rect 172 58 179 60
rect 172 56 175 58
rect 177 56 179 58
rect 172 51 179 56
rect 172 49 175 51
rect 177 49 179 51
rect 184 59 186 61
rect 188 59 191 61
rect 184 54 191 59
rect 184 52 186 54
rect 188 52 191 54
rect 184 50 191 52
rect 193 73 202 75
rect 193 71 197 73
rect 199 71 202 73
rect 284 76 291 78
rect 284 75 286 76
rect 225 73 239 75
rect 225 72 232 73
rect 193 63 202 71
rect 209 63 214 72
rect 193 50 204 63
rect 206 54 214 63
rect 206 52 209 54
rect 211 52 214 54
rect 206 50 214 52
rect 172 47 179 49
rect 209 47 214 50
rect 216 47 221 72
rect 223 71 232 72
rect 234 71 239 73
rect 223 66 239 71
rect 223 64 232 66
rect 234 64 239 66
rect 223 47 239 64
rect 241 65 249 75
rect 241 63 244 65
rect 246 63 249 65
rect 241 58 249 63
rect 241 56 244 58
rect 246 56 249 58
rect 241 47 249 56
rect 251 73 259 75
rect 251 71 254 73
rect 256 71 259 73
rect 251 66 259 71
rect 251 64 254 66
rect 256 64 259 66
rect 251 47 259 64
rect 261 60 266 75
rect 275 69 280 75
rect 273 67 280 69
rect 273 65 275 67
rect 277 65 280 67
rect 273 60 280 65
rect 261 58 268 60
rect 261 56 264 58
rect 266 56 268 58
rect 273 58 275 60
rect 277 58 280 60
rect 273 56 280 58
rect 261 51 268 56
rect 261 49 264 51
rect 266 49 268 51
rect 261 47 268 49
rect 275 47 280 56
rect 282 74 286 75
rect 288 75 291 76
rect 288 74 293 75
rect 282 47 293 74
rect 295 47 300 75
rect 302 69 307 75
rect 302 67 309 69
rect 302 65 305 67
rect 307 65 309 67
rect 302 63 309 65
rect 321 66 328 68
rect 321 64 323 66
rect 325 64 328 66
rect 302 47 307 63
rect 321 55 328 64
rect 330 66 338 68
rect 330 64 333 66
rect 335 64 338 66
rect 330 59 338 64
rect 330 57 333 59
rect 335 57 338 59
rect 330 55 338 57
rect 340 66 346 68
rect 340 64 348 66
rect 340 62 343 64
rect 345 62 348 64
rect 340 55 348 62
rect 342 48 348 55
rect 350 61 355 66
rect 365 63 370 75
rect 363 61 370 63
rect 350 59 357 61
rect 350 57 353 59
rect 355 57 357 59
rect 350 52 357 57
rect 350 50 353 52
rect 355 50 357 52
rect 363 59 365 61
rect 367 59 370 61
rect 363 54 370 59
rect 363 52 365 54
rect 367 52 370 54
rect 363 50 370 52
rect 372 73 381 75
rect 372 71 376 73
rect 378 71 381 73
rect 404 73 418 75
rect 404 72 411 73
rect 372 63 381 71
rect 388 63 393 72
rect 372 50 383 63
rect 385 54 393 63
rect 385 52 388 54
rect 390 52 393 54
rect 385 50 393 52
rect 350 48 357 50
rect 388 47 393 50
rect 395 47 400 72
rect 402 71 411 72
rect 413 71 418 73
rect 402 66 418 71
rect 402 64 411 66
rect 413 64 418 66
rect 402 47 418 64
rect 420 65 428 75
rect 420 63 423 65
rect 425 63 428 65
rect 420 58 428 63
rect 420 56 423 58
rect 425 56 428 58
rect 420 47 428 56
rect 430 73 438 75
rect 430 71 433 73
rect 435 71 438 73
rect 430 66 438 71
rect 430 64 433 66
rect 435 64 438 66
rect 430 47 438 64
rect 440 60 445 75
rect 454 63 459 75
rect 452 61 459 63
rect 440 58 447 60
rect 440 56 443 58
rect 445 56 447 58
rect 440 51 447 56
rect 440 49 443 51
rect 445 49 447 51
rect 452 59 454 61
rect 456 59 459 61
rect 452 54 459 59
rect 452 52 454 54
rect 456 52 459 54
rect 452 50 459 52
rect 461 73 470 75
rect 461 71 465 73
rect 467 71 470 73
rect 552 76 559 78
rect 552 75 554 76
rect 493 73 507 75
rect 493 72 500 73
rect 461 63 470 71
rect 477 63 482 72
rect 461 50 472 63
rect 474 54 482 63
rect 474 52 477 54
rect 479 52 482 54
rect 474 50 482 52
rect 440 47 447 49
rect 477 47 482 50
rect 484 47 489 72
rect 491 71 500 72
rect 502 71 507 73
rect 491 66 507 71
rect 491 64 500 66
rect 502 64 507 66
rect 491 47 507 64
rect 509 65 517 75
rect 509 63 512 65
rect 514 63 517 65
rect 509 58 517 63
rect 509 56 512 58
rect 514 56 517 58
rect 509 47 517 56
rect 519 73 527 75
rect 519 71 522 73
rect 524 71 527 73
rect 519 66 527 71
rect 519 64 522 66
rect 524 64 527 66
rect 519 47 527 64
rect 529 60 534 75
rect 543 69 548 75
rect 541 67 548 69
rect 541 65 543 67
rect 545 65 548 67
rect 541 60 548 65
rect 529 58 536 60
rect 529 56 532 58
rect 534 56 536 58
rect 541 58 543 60
rect 545 58 548 60
rect 541 56 548 58
rect 529 51 536 56
rect 529 49 532 51
rect 534 49 536 51
rect 529 47 536 49
rect 543 47 548 56
rect 550 74 554 75
rect 556 75 559 76
rect 556 74 561 75
rect 550 47 561 74
rect 563 47 568 75
rect 570 69 575 75
rect 570 67 577 69
rect 570 65 573 67
rect 575 65 577 67
rect 570 63 577 65
rect 589 66 596 68
rect 589 64 591 66
rect 593 64 596 66
rect 570 47 575 63
rect 589 55 596 64
rect 598 66 606 68
rect 598 64 601 66
rect 603 64 606 66
rect 598 59 606 64
rect 598 57 601 59
rect 603 57 606 59
rect 598 55 606 57
rect 608 66 614 68
rect 608 64 616 66
rect 608 62 611 64
rect 613 62 616 64
rect 608 55 616 62
rect 610 48 616 55
rect 618 61 623 66
rect 632 63 637 75
rect 630 61 637 63
rect 618 59 625 61
rect 618 57 621 59
rect 623 57 625 59
rect 618 52 625 57
rect 618 50 621 52
rect 623 50 625 52
rect 630 59 632 61
rect 634 59 637 61
rect 630 54 637 59
rect 630 52 632 54
rect 634 52 637 54
rect 630 50 637 52
rect 639 73 648 75
rect 639 71 643 73
rect 645 71 648 73
rect 671 73 685 75
rect 671 72 678 73
rect 639 63 648 71
rect 655 63 660 72
rect 639 50 650 63
rect 652 54 660 63
rect 652 52 655 54
rect 657 52 660 54
rect 652 50 660 52
rect 618 48 625 50
rect 655 47 660 50
rect 662 47 667 72
rect 669 71 678 72
rect 680 71 685 73
rect 669 66 685 71
rect 669 64 678 66
rect 680 64 685 66
rect 669 47 685 64
rect 687 65 695 75
rect 687 63 690 65
rect 692 63 695 65
rect 687 58 695 63
rect 687 56 690 58
rect 692 56 695 58
rect 687 47 695 56
rect 697 73 705 75
rect 697 71 700 73
rect 702 71 705 73
rect 697 66 705 71
rect 697 64 700 66
rect 702 64 705 66
rect 697 47 705 64
rect 707 60 712 75
rect 721 63 726 75
rect 719 61 726 63
rect 707 58 714 60
rect 707 56 710 58
rect 712 56 714 58
rect 707 51 714 56
rect 707 49 710 51
rect 712 49 714 51
rect 719 59 721 61
rect 723 59 726 61
rect 719 54 726 59
rect 719 52 721 54
rect 723 52 726 54
rect 719 50 726 52
rect 728 73 737 75
rect 728 71 732 73
rect 734 71 737 73
rect 819 76 826 78
rect 819 75 821 76
rect 760 73 774 75
rect 760 72 767 73
rect 728 63 737 71
rect 744 63 749 72
rect 728 50 739 63
rect 741 54 749 63
rect 741 52 744 54
rect 746 52 749 54
rect 741 50 749 52
rect 707 47 714 49
rect 744 47 749 50
rect 751 47 756 72
rect 758 71 767 72
rect 769 71 774 73
rect 758 66 774 71
rect 758 64 767 66
rect 769 64 774 66
rect 758 47 774 64
rect 776 65 784 75
rect 776 63 779 65
rect 781 63 784 65
rect 776 58 784 63
rect 776 56 779 58
rect 781 56 784 58
rect 776 47 784 56
rect 786 73 794 75
rect 786 71 789 73
rect 791 71 794 73
rect 786 66 794 71
rect 786 64 789 66
rect 791 64 794 66
rect 786 47 794 64
rect 796 60 801 75
rect 810 69 815 75
rect 808 67 815 69
rect 808 65 810 67
rect 812 65 815 67
rect 808 60 815 65
rect 796 58 803 60
rect 796 56 799 58
rect 801 56 803 58
rect 808 58 810 60
rect 812 58 815 60
rect 808 56 815 58
rect 796 51 803 56
rect 796 49 799 51
rect 801 49 803 51
rect 796 47 803 49
rect 810 47 815 56
rect 817 74 821 75
rect 823 75 826 76
rect 823 74 828 75
rect 817 47 828 74
rect 830 47 835 75
rect 837 69 842 75
rect 837 67 844 69
rect 837 65 840 67
rect 842 65 844 67
rect 837 63 844 65
rect 837 47 842 63
<< alu1 >>
rect 12 305 838 306
rect 12 303 25 305
rect 27 303 59 305
rect 61 303 318 305
rect 320 303 595 305
rect 597 303 838 305
rect 12 302 838 303
rect 0 292 848 297
rect 0 290 34 292
rect 36 290 44 292
rect 46 290 74 292
rect 76 290 84 292
rect 86 290 144 292
rect 146 290 302 292
rect 304 290 342 292
rect 344 290 352 292
rect 354 290 570 292
rect 572 290 610 292
rect 612 290 620 292
rect 622 290 837 292
rect 839 290 848 292
rect 0 289 848 290
rect 0 161 4 289
rect 20 275 25 276
rect 20 273 22 275
rect 24 273 25 275
rect 20 267 25 273
rect 37 280 49 284
rect 37 278 45 280
rect 47 278 49 280
rect 20 266 34 267
rect 20 264 28 266
rect 30 264 34 266
rect 20 263 34 264
rect 13 258 26 259
rect 13 256 18 258
rect 20 256 26 258
rect 13 255 26 256
rect 13 249 17 255
rect 45 274 49 278
rect 45 272 46 274
rect 48 272 49 274
rect 45 258 49 272
rect 60 267 65 276
rect 77 280 89 284
rect 77 278 85 280
rect 87 278 89 280
rect 60 266 74 267
rect 60 264 62 266
rect 64 264 68 266
rect 70 264 74 266
rect 60 263 74 264
rect 13 247 14 249
rect 16 247 17 249
rect 13 246 17 247
rect 44 256 49 258
rect 44 254 45 256
rect 47 254 49 256
rect 44 249 49 254
rect 44 247 45 249
rect 47 247 49 249
rect 44 245 49 247
rect 53 258 66 259
rect 53 256 54 258
rect 56 256 58 258
rect 60 256 66 258
rect 53 255 66 256
rect 53 246 57 255
rect 85 262 89 278
rect 85 260 86 262
rect 88 260 89 262
rect 85 258 89 260
rect 84 256 89 258
rect 84 254 85 256
rect 87 254 89 256
rect 84 249 89 254
rect 84 247 85 249
rect 87 247 89 249
rect 84 245 89 247
rect 95 282 100 284
rect 95 280 97 282
rect 99 280 100 282
rect 95 278 100 280
rect 95 266 99 278
rect 158 282 180 283
rect 158 280 175 282
rect 177 280 180 282
rect 158 279 180 280
rect 143 274 147 276
rect 143 272 144 274
rect 146 272 147 274
rect 95 264 96 266
rect 98 264 99 266
rect 95 256 99 264
rect 95 254 100 256
rect 95 252 97 254
rect 99 252 100 254
rect 95 247 100 252
rect 123 266 131 268
rect 143 267 147 272
rect 176 274 180 279
rect 176 272 177 274
rect 179 272 180 274
rect 123 264 124 266
rect 126 264 131 266
rect 123 262 131 264
rect 141 266 156 267
rect 141 264 143 266
rect 145 264 150 266
rect 152 264 156 266
rect 141 263 156 264
rect 126 259 131 262
rect 126 258 164 259
rect 126 256 128 258
rect 130 256 164 258
rect 126 255 164 256
rect 176 259 180 272
rect 174 257 180 259
rect 174 255 175 257
rect 177 255 180 257
rect 174 250 180 255
rect 174 248 175 250
rect 177 248 180 250
rect 95 245 97 247
rect 99 245 100 247
rect 95 243 100 245
rect 174 246 180 248
rect 184 282 189 284
rect 184 280 186 282
rect 188 280 189 282
rect 184 278 189 280
rect 184 256 188 278
rect 247 282 269 283
rect 247 280 264 282
rect 266 280 269 282
rect 247 279 269 280
rect 184 254 189 256
rect 184 252 186 254
rect 188 252 189 254
rect 184 247 189 252
rect 212 266 220 268
rect 232 267 236 276
rect 212 264 213 266
rect 215 264 216 266
rect 218 264 220 266
rect 212 262 220 264
rect 230 266 245 267
rect 230 264 232 266
rect 234 264 236 266
rect 238 264 239 266
rect 241 264 245 266
rect 230 263 245 264
rect 215 259 220 262
rect 215 255 253 259
rect 265 260 269 279
rect 265 259 266 260
rect 263 258 266 259
rect 268 258 269 260
rect 263 257 269 258
rect 263 255 264 257
rect 266 255 269 257
rect 263 250 269 255
rect 263 248 264 250
rect 266 248 269 250
rect 184 245 186 247
rect 188 245 189 247
rect 184 243 189 245
rect 263 246 269 248
rect 273 282 278 284
rect 273 280 275 282
rect 277 280 278 282
rect 273 275 278 280
rect 273 273 275 275
rect 277 273 278 275
rect 273 271 278 273
rect 328 275 333 276
rect 328 273 330 275
rect 332 273 333 275
rect 273 248 277 271
rect 289 266 301 268
rect 289 264 292 266
rect 294 264 301 266
rect 289 262 301 264
rect 289 259 293 262
rect 289 257 290 259
rect 292 257 293 259
rect 289 254 293 257
rect 305 266 309 268
rect 307 264 309 266
rect 305 261 309 264
rect 328 267 333 273
rect 345 280 357 284
rect 345 278 353 280
rect 355 278 357 280
rect 328 266 342 267
rect 328 264 336 266
rect 338 264 342 266
rect 328 263 342 264
rect 305 259 306 261
rect 308 259 309 261
rect 305 252 309 259
rect 273 246 275 248
rect 273 244 277 246
rect 95 239 108 243
rect 184 242 197 243
rect 184 240 186 242
rect 188 240 197 242
rect 184 239 197 240
rect 273 242 285 244
rect 273 241 278 242
rect 273 239 275 241
rect 277 240 278 241
rect 280 240 285 242
rect 277 239 285 240
rect 273 238 285 239
rect 297 246 309 252
rect 321 258 334 259
rect 321 256 326 258
rect 328 256 334 258
rect 321 255 334 256
rect 321 250 325 255
rect 353 274 357 278
rect 353 272 354 274
rect 356 272 357 274
rect 353 258 357 272
rect 321 248 322 250
rect 324 248 325 250
rect 321 246 325 248
rect 352 256 357 258
rect 352 254 353 256
rect 355 254 357 256
rect 352 249 357 254
rect 352 247 353 249
rect 355 247 357 249
rect 352 245 357 247
rect 363 282 368 284
rect 363 280 365 282
rect 367 280 368 282
rect 363 278 368 280
rect 363 266 367 278
rect 426 282 448 283
rect 426 280 443 282
rect 445 280 448 282
rect 426 279 448 280
rect 411 274 415 276
rect 411 272 412 274
rect 414 272 415 274
rect 363 264 364 266
rect 366 264 367 266
rect 363 256 367 264
rect 363 254 368 256
rect 363 252 365 254
rect 367 252 368 254
rect 363 247 368 252
rect 391 266 399 268
rect 411 267 415 272
rect 444 274 448 279
rect 444 272 445 274
rect 447 272 448 274
rect 391 264 392 266
rect 394 264 399 266
rect 391 262 399 264
rect 409 266 424 267
rect 409 264 411 266
rect 413 264 418 266
rect 420 264 424 266
rect 409 263 424 264
rect 394 259 399 262
rect 394 258 432 259
rect 394 256 396 258
rect 398 256 432 258
rect 394 255 432 256
rect 444 259 448 272
rect 442 257 448 259
rect 442 255 443 257
rect 445 255 448 257
rect 442 250 448 255
rect 442 248 443 250
rect 445 248 448 250
rect 363 245 365 247
rect 367 245 368 247
rect 363 243 368 245
rect 442 246 448 248
rect 452 282 457 284
rect 452 280 454 282
rect 456 280 457 282
rect 452 278 457 280
rect 452 256 456 278
rect 515 282 537 283
rect 515 280 532 282
rect 534 280 537 282
rect 515 279 537 280
rect 452 254 457 256
rect 452 252 454 254
rect 456 252 457 254
rect 452 247 457 252
rect 480 266 488 268
rect 500 267 504 276
rect 480 264 481 266
rect 483 264 484 266
rect 486 264 488 266
rect 480 262 488 264
rect 498 266 513 267
rect 498 264 500 266
rect 502 264 504 266
rect 506 264 507 266
rect 509 264 513 266
rect 498 263 513 264
rect 483 259 488 262
rect 483 255 521 259
rect 533 260 537 279
rect 533 259 534 260
rect 531 258 534 259
rect 536 258 537 260
rect 531 257 537 258
rect 531 255 532 257
rect 534 255 537 257
rect 531 250 537 255
rect 531 248 532 250
rect 534 248 537 250
rect 452 245 454 247
rect 456 245 457 247
rect 452 243 457 245
rect 531 246 537 248
rect 541 282 546 284
rect 541 280 543 282
rect 545 280 546 282
rect 541 275 546 280
rect 541 273 543 275
rect 545 273 546 275
rect 541 271 546 273
rect 596 275 601 276
rect 596 273 598 275
rect 600 273 601 275
rect 541 248 545 271
rect 557 266 569 268
rect 557 264 560 266
rect 562 264 569 266
rect 557 262 569 264
rect 557 259 561 262
rect 557 257 558 259
rect 560 257 561 259
rect 557 254 561 257
rect 573 266 577 268
rect 575 264 577 266
rect 573 261 577 264
rect 596 267 601 273
rect 613 280 625 284
rect 613 278 621 280
rect 623 278 625 280
rect 596 266 610 267
rect 596 264 604 266
rect 606 264 610 266
rect 596 263 610 264
rect 573 259 574 261
rect 576 259 577 261
rect 573 252 577 259
rect 541 246 543 248
rect 541 244 545 246
rect 363 239 376 243
rect 452 242 465 243
rect 452 240 454 242
rect 456 240 465 242
rect 452 239 465 240
rect 541 241 553 244
rect 541 239 543 241
rect 545 239 546 241
rect 548 239 553 241
rect 541 238 553 239
rect 565 246 577 252
rect 589 258 602 259
rect 589 256 590 258
rect 592 256 594 258
rect 596 256 602 258
rect 589 255 602 256
rect 589 246 593 255
rect 621 274 625 278
rect 621 272 622 274
rect 624 272 625 274
rect 621 258 625 272
rect 620 256 625 258
rect 620 254 621 256
rect 623 254 625 256
rect 620 249 625 254
rect 620 247 621 249
rect 623 247 625 249
rect 620 245 625 247
rect 630 282 635 284
rect 630 280 632 282
rect 634 280 635 282
rect 630 278 635 280
rect 630 266 634 278
rect 693 282 715 283
rect 693 280 710 282
rect 712 280 715 282
rect 693 279 715 280
rect 678 274 682 276
rect 678 272 679 274
rect 681 272 682 274
rect 630 264 631 266
rect 633 264 634 266
rect 630 256 634 264
rect 630 254 635 256
rect 630 252 632 254
rect 634 252 635 254
rect 630 247 635 252
rect 658 266 666 268
rect 678 267 682 272
rect 711 274 715 279
rect 711 272 712 274
rect 714 272 715 274
rect 658 264 659 266
rect 661 264 666 266
rect 658 262 666 264
rect 676 266 691 267
rect 676 264 678 266
rect 680 264 685 266
rect 687 264 691 266
rect 676 263 691 264
rect 661 259 666 262
rect 661 258 699 259
rect 661 256 663 258
rect 665 256 699 258
rect 661 255 699 256
rect 711 259 715 272
rect 709 257 715 259
rect 709 255 710 257
rect 712 255 715 257
rect 709 250 715 255
rect 709 248 710 250
rect 712 248 715 250
rect 630 245 632 247
rect 634 245 635 247
rect 630 243 635 245
rect 709 246 715 248
rect 719 282 724 284
rect 719 280 721 282
rect 723 280 724 282
rect 719 278 724 280
rect 719 256 723 278
rect 782 282 804 283
rect 782 280 799 282
rect 801 280 804 282
rect 782 279 804 280
rect 719 254 724 256
rect 719 252 721 254
rect 723 252 724 254
rect 719 247 724 252
rect 747 266 755 268
rect 767 267 771 276
rect 747 264 748 266
rect 750 264 751 266
rect 753 264 755 266
rect 747 262 755 264
rect 765 266 780 267
rect 765 264 767 266
rect 769 264 771 266
rect 773 264 774 266
rect 776 264 780 266
rect 765 263 780 264
rect 750 259 755 262
rect 750 255 788 259
rect 800 260 804 279
rect 800 259 801 260
rect 798 258 801 259
rect 803 258 804 260
rect 798 257 804 258
rect 798 255 799 257
rect 801 255 804 257
rect 798 250 804 255
rect 798 248 799 250
rect 801 248 804 250
rect 719 245 721 247
rect 723 245 724 247
rect 719 243 724 245
rect 798 246 804 248
rect 808 282 813 284
rect 808 280 810 282
rect 812 280 813 282
rect 808 275 813 280
rect 808 273 810 275
rect 812 273 813 275
rect 808 271 813 273
rect 808 248 812 271
rect 824 266 836 268
rect 824 264 827 266
rect 829 264 836 266
rect 824 262 836 264
rect 824 259 828 262
rect 824 257 825 259
rect 827 257 828 259
rect 824 254 828 257
rect 840 266 844 268
rect 842 264 844 266
rect 840 261 844 264
rect 840 259 841 261
rect 843 259 844 261
rect 840 252 844 259
rect 808 246 810 248
rect 808 244 812 246
rect 630 239 643 243
rect 719 242 732 243
rect 719 240 721 242
rect 723 240 732 242
rect 719 239 732 240
rect 808 242 820 244
rect 808 241 813 242
rect 808 239 810 241
rect 812 240 813 241
rect 815 240 820 242
rect 812 239 820 240
rect 808 238 820 239
rect 832 246 844 252
rect 9 232 857 233
rect 9 230 44 232
rect 46 230 84 232
rect 86 230 286 232
rect 288 230 352 232
rect 354 230 554 232
rect 556 230 620 232
rect 622 230 821 232
rect 823 230 857 232
rect 9 220 857 230
rect 9 218 44 220
rect 46 218 84 220
rect 86 218 286 220
rect 288 218 352 220
rect 354 218 554 220
rect 556 218 620 220
rect 622 218 821 220
rect 823 218 857 220
rect 9 217 857 218
rect 13 203 17 204
rect 13 201 14 203
rect 16 201 17 203
rect 13 195 17 201
rect 44 203 49 205
rect 13 194 26 195
rect 13 192 18 194
rect 20 192 26 194
rect 13 191 26 192
rect 20 186 34 187
rect 20 184 28 186
rect 30 184 34 186
rect 20 183 34 184
rect 44 201 45 203
rect 47 201 49 203
rect 44 196 49 201
rect 44 194 45 196
rect 47 194 49 196
rect 44 192 49 194
rect 20 177 25 183
rect 20 175 22 177
rect 24 175 25 177
rect 20 174 25 175
rect 45 178 49 192
rect 53 195 57 204
rect 95 207 108 211
rect 184 210 197 211
rect 184 208 186 210
rect 188 208 197 210
rect 184 207 197 208
rect 273 211 285 212
rect 273 209 275 211
rect 277 210 285 211
rect 277 209 278 210
rect 273 208 278 209
rect 280 208 285 210
rect 95 205 100 207
rect 84 203 89 205
rect 53 194 66 195
rect 53 192 54 194
rect 56 192 58 194
rect 60 192 66 194
rect 53 191 66 192
rect 45 176 46 178
rect 48 176 49 178
rect 45 172 49 176
rect 60 186 74 187
rect 60 184 62 186
rect 64 184 68 186
rect 70 184 74 186
rect 60 183 74 184
rect 84 201 85 203
rect 87 201 89 203
rect 84 196 89 201
rect 84 194 85 196
rect 87 194 89 196
rect 84 192 89 194
rect 60 174 65 183
rect 85 190 89 192
rect 85 188 86 190
rect 88 188 89 190
rect 37 170 45 172
rect 47 170 49 172
rect 85 172 89 188
rect 37 166 49 170
rect 77 170 85 172
rect 87 170 89 172
rect 77 166 89 170
rect 95 203 97 205
rect 99 203 100 205
rect 184 205 189 207
rect 95 198 100 203
rect 95 196 97 198
rect 99 196 100 198
rect 95 194 100 196
rect 95 186 99 194
rect 95 184 96 186
rect 98 184 99 186
rect 126 194 164 195
rect 126 192 128 194
rect 130 192 164 194
rect 126 191 164 192
rect 95 172 99 184
rect 126 188 131 191
rect 123 186 131 188
rect 123 184 124 186
rect 126 184 131 186
rect 123 182 131 184
rect 141 186 156 187
rect 141 184 143 186
rect 145 184 150 186
rect 152 184 156 186
rect 141 183 156 184
rect 95 170 100 172
rect 143 178 147 183
rect 174 202 180 204
rect 174 200 175 202
rect 177 200 180 202
rect 174 195 180 200
rect 174 193 175 195
rect 177 193 180 195
rect 174 191 180 193
rect 143 176 144 178
rect 146 176 147 178
rect 143 174 147 176
rect 176 178 180 191
rect 176 176 177 178
rect 179 176 180 178
rect 176 171 180 176
rect 95 168 97 170
rect 99 168 100 170
rect 95 166 100 168
rect 158 170 180 171
rect 158 168 175 170
rect 177 168 180 170
rect 158 167 180 168
rect 184 203 186 205
rect 188 203 189 205
rect 273 206 285 208
rect 273 204 277 206
rect 184 198 189 203
rect 184 196 186 198
rect 188 196 189 198
rect 184 194 189 196
rect 184 172 188 194
rect 215 191 253 195
rect 215 188 220 191
rect 212 186 220 188
rect 212 184 213 186
rect 215 184 216 186
rect 218 184 220 186
rect 212 182 220 184
rect 230 186 245 187
rect 230 184 232 186
rect 234 184 236 186
rect 238 184 239 186
rect 241 184 245 186
rect 230 183 245 184
rect 184 170 189 172
rect 232 174 236 183
rect 263 202 269 204
rect 263 200 264 202
rect 266 200 269 202
rect 263 195 269 200
rect 263 193 264 195
rect 266 193 269 195
rect 263 192 269 193
rect 263 191 266 192
rect 265 190 266 191
rect 268 190 269 192
rect 265 171 269 190
rect 184 168 186 170
rect 188 168 189 170
rect 184 166 189 168
rect 247 170 269 171
rect 247 168 264 170
rect 266 168 269 170
rect 247 167 269 168
rect 273 202 275 204
rect 273 179 277 202
rect 297 198 309 204
rect 273 177 278 179
rect 273 175 275 177
rect 277 175 278 177
rect 273 170 278 175
rect 289 193 293 196
rect 289 191 290 193
rect 292 191 293 193
rect 289 188 293 191
rect 289 186 301 188
rect 289 184 292 186
rect 294 184 301 186
rect 289 182 301 184
rect 305 191 309 198
rect 321 203 325 204
rect 321 201 322 203
rect 324 201 325 203
rect 321 195 325 201
rect 363 207 376 211
rect 452 210 465 211
rect 452 208 454 210
rect 456 208 465 210
rect 452 207 465 208
rect 541 211 553 212
rect 541 209 543 211
rect 545 210 553 211
rect 545 209 546 210
rect 541 208 546 209
rect 548 208 553 210
rect 363 205 368 207
rect 352 203 357 205
rect 321 194 334 195
rect 321 192 326 194
rect 328 192 334 194
rect 321 191 334 192
rect 305 189 306 191
rect 308 189 309 191
rect 305 186 309 189
rect 307 184 309 186
rect 305 182 309 184
rect 328 186 342 187
rect 328 184 336 186
rect 338 184 342 186
rect 328 183 342 184
rect 352 201 353 203
rect 355 201 357 203
rect 352 196 357 201
rect 352 194 353 196
rect 355 194 357 196
rect 352 192 357 194
rect 328 177 333 183
rect 328 175 330 177
rect 332 175 333 177
rect 328 174 333 175
rect 353 178 357 192
rect 353 176 354 178
rect 356 176 357 178
rect 273 168 275 170
rect 277 168 278 170
rect 273 166 278 168
rect 353 172 357 176
rect 345 170 353 172
rect 355 170 357 172
rect 345 166 357 170
rect 363 203 365 205
rect 367 203 368 205
rect 452 205 457 207
rect 363 198 368 203
rect 363 196 365 198
rect 367 196 368 198
rect 363 194 368 196
rect 363 186 367 194
rect 363 184 364 186
rect 366 184 367 186
rect 394 194 432 195
rect 394 192 396 194
rect 398 192 432 194
rect 394 191 432 192
rect 363 172 367 184
rect 394 188 399 191
rect 391 186 399 188
rect 391 184 392 186
rect 394 184 399 186
rect 391 182 399 184
rect 409 186 424 187
rect 409 184 411 186
rect 413 184 418 186
rect 420 184 424 186
rect 409 183 424 184
rect 363 170 368 172
rect 411 178 415 183
rect 442 202 448 204
rect 442 200 443 202
rect 445 200 448 202
rect 442 195 448 200
rect 442 193 443 195
rect 445 193 448 195
rect 442 191 448 193
rect 411 176 412 178
rect 414 176 415 178
rect 411 174 415 176
rect 444 178 448 191
rect 444 176 445 178
rect 447 176 448 178
rect 444 171 448 176
rect 363 168 365 170
rect 367 168 368 170
rect 363 166 368 168
rect 426 170 448 171
rect 426 168 443 170
rect 445 168 448 170
rect 426 167 448 168
rect 452 203 454 205
rect 456 203 457 205
rect 541 206 553 208
rect 541 204 545 206
rect 452 198 457 203
rect 452 196 454 198
rect 456 196 457 198
rect 452 194 457 196
rect 452 172 456 194
rect 483 191 521 195
rect 483 188 488 191
rect 480 186 488 188
rect 480 184 481 186
rect 483 184 484 186
rect 486 184 488 186
rect 480 182 488 184
rect 498 186 513 187
rect 498 184 500 186
rect 502 184 504 186
rect 506 184 507 186
rect 509 184 513 186
rect 498 183 513 184
rect 452 170 457 172
rect 500 174 504 183
rect 531 202 537 204
rect 531 200 532 202
rect 534 200 537 202
rect 531 195 537 200
rect 531 193 532 195
rect 534 193 537 195
rect 531 192 537 193
rect 531 191 534 192
rect 533 190 534 191
rect 536 190 537 192
rect 533 171 537 190
rect 452 168 454 170
rect 456 168 457 170
rect 452 166 457 168
rect 515 170 537 171
rect 515 168 532 170
rect 534 168 537 170
rect 515 167 537 168
rect 541 202 543 204
rect 541 179 545 202
rect 565 198 577 204
rect 541 177 546 179
rect 541 175 543 177
rect 545 175 546 177
rect 541 170 546 175
rect 557 193 561 196
rect 557 191 558 193
rect 560 191 561 193
rect 557 188 561 191
rect 557 186 569 188
rect 557 184 560 186
rect 562 184 569 186
rect 557 182 569 184
rect 573 191 577 198
rect 589 203 593 204
rect 589 201 590 203
rect 592 201 593 203
rect 589 195 593 201
rect 630 207 643 211
rect 719 210 732 211
rect 719 208 721 210
rect 723 208 732 210
rect 719 207 732 208
rect 808 211 820 212
rect 808 209 810 211
rect 812 210 820 211
rect 812 209 813 210
rect 808 208 813 209
rect 815 208 820 210
rect 630 205 635 207
rect 620 203 625 205
rect 589 194 602 195
rect 589 192 594 194
rect 596 192 602 194
rect 589 191 602 192
rect 573 189 574 191
rect 576 189 577 191
rect 573 186 577 189
rect 575 184 577 186
rect 573 182 577 184
rect 596 186 610 187
rect 596 184 604 186
rect 606 184 610 186
rect 596 183 610 184
rect 620 201 621 203
rect 623 201 625 203
rect 620 196 625 201
rect 620 194 621 196
rect 623 194 625 196
rect 620 192 625 194
rect 596 177 601 183
rect 596 175 598 177
rect 600 175 601 177
rect 596 174 601 175
rect 621 178 625 192
rect 621 176 622 178
rect 624 176 625 178
rect 541 168 543 170
rect 545 168 546 170
rect 541 166 546 168
rect 621 172 625 176
rect 613 170 621 172
rect 623 170 625 172
rect 613 166 625 170
rect 630 203 632 205
rect 634 203 635 205
rect 719 205 724 207
rect 630 198 635 203
rect 630 196 632 198
rect 634 196 635 198
rect 630 194 635 196
rect 630 186 634 194
rect 630 184 631 186
rect 633 184 634 186
rect 661 194 699 195
rect 661 192 663 194
rect 665 192 699 194
rect 661 191 699 192
rect 630 172 634 184
rect 661 188 666 191
rect 658 186 666 188
rect 658 184 659 186
rect 661 184 666 186
rect 658 182 666 184
rect 676 186 691 187
rect 676 184 678 186
rect 680 184 685 186
rect 687 184 691 186
rect 676 183 691 184
rect 630 170 635 172
rect 678 178 682 183
rect 709 202 715 204
rect 709 200 710 202
rect 712 200 715 202
rect 709 195 715 200
rect 709 193 710 195
rect 712 193 715 195
rect 709 191 715 193
rect 678 176 679 178
rect 681 176 682 178
rect 678 174 682 176
rect 711 178 715 191
rect 711 176 712 178
rect 714 176 715 178
rect 711 171 715 176
rect 630 168 632 170
rect 634 168 635 170
rect 630 166 635 168
rect 693 170 715 171
rect 693 168 710 170
rect 712 168 715 170
rect 693 167 715 168
rect 719 203 721 205
rect 723 203 724 205
rect 808 206 820 208
rect 808 204 812 206
rect 719 198 724 203
rect 719 196 721 198
rect 723 196 724 198
rect 719 194 724 196
rect 719 172 723 194
rect 750 191 788 195
rect 750 188 755 191
rect 747 186 755 188
rect 747 184 748 186
rect 750 184 751 186
rect 753 184 755 186
rect 747 182 755 184
rect 765 186 780 187
rect 765 184 767 186
rect 769 184 771 186
rect 773 184 774 186
rect 776 184 780 186
rect 765 183 780 184
rect 719 170 724 172
rect 767 174 771 183
rect 798 202 804 204
rect 798 200 799 202
rect 801 200 804 202
rect 798 195 804 200
rect 798 193 799 195
rect 801 193 804 195
rect 798 192 804 193
rect 798 191 801 192
rect 800 190 801 191
rect 803 190 804 192
rect 800 171 804 190
rect 719 168 721 170
rect 723 168 724 170
rect 719 166 724 168
rect 782 170 804 171
rect 782 168 799 170
rect 801 168 804 170
rect 782 167 804 168
rect 808 202 810 204
rect 808 179 812 202
rect 832 198 844 204
rect 808 177 813 179
rect 808 175 810 177
rect 812 175 813 177
rect 808 170 813 175
rect 824 193 828 196
rect 824 191 825 193
rect 827 191 828 193
rect 824 188 828 191
rect 824 186 836 188
rect 824 184 827 186
rect 829 184 836 186
rect 824 182 836 184
rect 840 191 844 198
rect 840 189 841 191
rect 843 189 844 191
rect 840 186 844 189
rect 842 184 844 186
rect 840 182 844 184
rect 808 168 810 170
rect 812 168 813 170
rect 808 166 813 168
rect 0 160 848 161
rect 0 158 34 160
rect 36 158 44 160
rect 46 158 74 160
rect 76 158 84 160
rect 86 158 302 160
rect 304 158 342 160
rect 344 158 352 160
rect 354 158 570 160
rect 572 158 610 160
rect 612 158 620 160
rect 622 158 837 160
rect 839 158 848 160
rect 0 148 848 158
rect 0 146 34 148
rect 36 146 44 148
rect 46 146 74 148
rect 76 146 84 148
rect 86 146 302 148
rect 304 146 342 148
rect 344 146 352 148
rect 354 146 570 148
rect 572 146 610 148
rect 612 146 620 148
rect 622 146 837 148
rect 839 146 848 148
rect 0 145 848 146
rect 0 17 4 145
rect 20 131 25 132
rect 20 129 22 131
rect 24 129 25 131
rect 20 123 25 129
rect 37 136 49 140
rect 37 134 45 136
rect 47 134 49 136
rect 20 122 34 123
rect 20 120 28 122
rect 30 120 34 122
rect 20 119 34 120
rect 13 114 26 115
rect 13 112 18 114
rect 20 112 21 114
rect 23 112 26 114
rect 13 111 26 112
rect 13 102 17 111
rect 45 130 49 134
rect 45 128 46 130
rect 48 128 49 130
rect 45 114 49 128
rect 60 123 65 132
rect 77 136 89 140
rect 77 134 85 136
rect 87 134 89 136
rect 60 122 74 123
rect 60 120 62 122
rect 64 120 68 122
rect 70 120 74 122
rect 60 119 74 120
rect 44 112 49 114
rect 44 110 45 112
rect 47 110 49 112
rect 44 105 49 110
rect 44 103 45 105
rect 47 103 49 105
rect 44 101 49 103
rect 53 114 66 115
rect 53 112 54 114
rect 56 112 58 114
rect 60 112 66 114
rect 53 111 66 112
rect 53 102 57 111
rect 85 118 89 134
rect 85 116 86 118
rect 88 116 89 118
rect 85 114 89 116
rect 84 112 89 114
rect 84 110 85 112
rect 87 110 89 112
rect 84 105 89 110
rect 84 103 85 105
rect 87 103 89 105
rect 84 101 89 103
rect 95 138 100 140
rect 95 136 97 138
rect 99 136 100 138
rect 95 134 100 136
rect 95 122 99 134
rect 158 138 180 139
rect 158 136 175 138
rect 177 136 180 138
rect 158 135 180 136
rect 143 130 147 132
rect 143 128 144 130
rect 146 128 147 130
rect 95 120 96 122
rect 98 120 99 122
rect 95 112 99 120
rect 95 110 100 112
rect 95 108 97 110
rect 99 108 100 110
rect 95 103 100 108
rect 123 122 131 124
rect 143 123 147 128
rect 176 130 180 135
rect 176 128 177 130
rect 179 128 180 130
rect 123 120 124 122
rect 126 120 131 122
rect 123 118 131 120
rect 141 122 156 123
rect 141 120 143 122
rect 145 120 150 122
rect 152 120 156 122
rect 141 119 156 120
rect 126 115 131 118
rect 126 114 164 115
rect 126 112 128 114
rect 130 112 164 114
rect 126 111 164 112
rect 176 115 180 128
rect 174 113 180 115
rect 174 111 175 113
rect 177 111 180 113
rect 174 106 180 111
rect 174 104 175 106
rect 177 104 180 106
rect 95 101 97 103
rect 99 101 100 103
rect 95 99 100 101
rect 174 102 180 104
rect 184 138 189 140
rect 184 136 186 138
rect 188 136 189 138
rect 184 134 189 136
rect 184 112 188 134
rect 247 138 269 139
rect 247 136 264 138
rect 266 136 269 138
rect 247 135 269 136
rect 184 110 189 112
rect 184 108 186 110
rect 188 108 189 110
rect 184 103 189 108
rect 212 122 220 124
rect 232 123 236 132
rect 212 120 213 122
rect 215 120 216 122
rect 218 120 220 122
rect 212 118 220 120
rect 230 122 245 123
rect 230 120 232 122
rect 234 120 236 122
rect 238 120 239 122
rect 241 120 245 122
rect 230 119 245 120
rect 215 115 220 118
rect 215 111 253 115
rect 265 116 269 135
rect 265 115 266 116
rect 263 114 266 115
rect 268 114 269 116
rect 263 113 269 114
rect 263 111 264 113
rect 266 111 269 113
rect 263 106 269 111
rect 263 104 264 106
rect 266 104 269 106
rect 184 101 186 103
rect 188 101 189 103
rect 184 99 189 101
rect 263 102 269 104
rect 273 138 278 140
rect 273 136 275 138
rect 277 136 278 138
rect 273 131 278 136
rect 273 129 275 131
rect 277 129 278 131
rect 273 127 278 129
rect 328 130 333 132
rect 328 128 329 130
rect 331 128 333 130
rect 273 104 277 127
rect 289 122 301 124
rect 289 120 292 122
rect 294 120 301 122
rect 289 118 301 120
rect 289 115 293 118
rect 289 113 290 115
rect 292 113 293 115
rect 289 110 293 113
rect 305 122 309 124
rect 307 120 309 122
rect 305 117 309 120
rect 328 123 333 128
rect 345 136 357 140
rect 345 134 353 136
rect 355 134 357 136
rect 328 122 342 123
rect 328 120 336 122
rect 338 120 342 122
rect 328 119 342 120
rect 305 115 306 117
rect 308 115 309 117
rect 305 108 309 115
rect 273 102 275 104
rect 273 100 277 102
rect 95 95 108 99
rect 184 98 197 99
rect 184 96 186 98
rect 188 96 197 98
rect 184 95 197 96
rect 273 98 285 100
rect 273 97 278 98
rect 273 95 275 97
rect 277 96 278 97
rect 280 96 285 98
rect 277 95 285 96
rect 273 94 285 95
rect 297 102 309 108
rect 321 114 334 115
rect 321 112 326 114
rect 328 112 334 114
rect 321 111 334 112
rect 321 105 325 111
rect 353 130 357 134
rect 353 128 354 130
rect 356 128 357 130
rect 353 114 357 128
rect 321 103 322 105
rect 324 103 325 105
rect 321 102 325 103
rect 352 112 357 114
rect 352 110 353 112
rect 355 110 357 112
rect 352 105 357 110
rect 352 103 353 105
rect 355 103 357 105
rect 352 101 357 103
rect 363 138 368 140
rect 363 136 365 138
rect 367 136 368 138
rect 363 134 368 136
rect 363 122 367 134
rect 426 138 448 139
rect 426 136 443 138
rect 445 136 448 138
rect 426 135 448 136
rect 411 130 415 132
rect 411 128 412 130
rect 414 128 415 130
rect 363 120 364 122
rect 366 120 367 122
rect 363 112 367 120
rect 363 110 368 112
rect 363 108 365 110
rect 367 108 368 110
rect 363 103 368 108
rect 391 122 399 124
rect 411 123 415 128
rect 444 130 448 135
rect 444 128 445 130
rect 447 128 448 130
rect 391 120 392 122
rect 394 120 399 122
rect 391 118 399 120
rect 409 122 424 123
rect 409 120 411 122
rect 413 120 418 122
rect 420 120 424 122
rect 409 119 424 120
rect 394 115 399 118
rect 394 114 432 115
rect 394 112 396 114
rect 398 112 432 114
rect 394 111 432 112
rect 444 115 448 128
rect 442 113 448 115
rect 442 111 443 113
rect 445 111 448 113
rect 442 106 448 111
rect 442 104 443 106
rect 445 104 448 106
rect 363 101 365 103
rect 367 101 368 103
rect 363 99 368 101
rect 442 102 448 104
rect 452 138 457 140
rect 452 136 454 138
rect 456 136 457 138
rect 452 134 457 136
rect 452 112 456 134
rect 515 138 537 139
rect 515 136 532 138
rect 534 136 537 138
rect 515 135 537 136
rect 452 110 457 112
rect 452 108 454 110
rect 456 108 457 110
rect 452 103 457 108
rect 480 122 488 124
rect 500 123 504 132
rect 480 120 481 122
rect 483 120 484 122
rect 486 120 488 122
rect 480 118 488 120
rect 498 122 513 123
rect 498 120 500 122
rect 502 120 504 122
rect 506 120 507 122
rect 509 120 513 122
rect 498 119 513 120
rect 483 115 488 118
rect 483 111 521 115
rect 533 116 537 135
rect 533 115 534 116
rect 531 114 534 115
rect 536 114 537 116
rect 531 113 537 114
rect 531 111 532 113
rect 534 111 537 113
rect 531 106 537 111
rect 531 104 532 106
rect 534 104 537 106
rect 452 101 454 103
rect 456 101 457 103
rect 452 99 457 101
rect 531 102 537 104
rect 541 138 546 140
rect 541 136 543 138
rect 545 136 546 138
rect 541 131 546 136
rect 541 129 543 131
rect 545 129 546 131
rect 541 127 546 129
rect 596 131 601 132
rect 596 129 598 131
rect 600 129 601 131
rect 541 104 545 127
rect 557 122 569 124
rect 557 120 560 122
rect 562 120 569 122
rect 557 118 569 120
rect 557 115 561 118
rect 557 113 558 115
rect 560 113 561 115
rect 557 110 561 113
rect 573 122 577 124
rect 575 120 577 122
rect 573 117 577 120
rect 596 123 601 129
rect 613 136 625 140
rect 613 134 621 136
rect 623 134 625 136
rect 596 122 610 123
rect 596 120 604 122
rect 606 120 610 122
rect 596 119 610 120
rect 573 115 574 117
rect 576 115 577 117
rect 573 108 577 115
rect 541 102 543 104
rect 541 100 545 102
rect 363 95 376 99
rect 452 98 465 99
rect 452 96 454 98
rect 456 96 465 98
rect 452 95 465 96
rect 541 98 553 100
rect 541 97 546 98
rect 541 95 543 97
rect 545 96 546 97
rect 548 96 553 98
rect 545 95 553 96
rect 541 94 553 95
rect 565 102 577 108
rect 589 114 602 115
rect 589 112 594 114
rect 596 112 602 114
rect 589 111 602 112
rect 589 105 593 111
rect 621 130 625 134
rect 621 128 622 130
rect 624 128 625 130
rect 621 114 625 128
rect 589 103 590 105
rect 592 103 593 105
rect 589 102 593 103
rect 620 112 625 114
rect 620 110 621 112
rect 623 110 625 112
rect 620 105 625 110
rect 620 103 621 105
rect 623 103 625 105
rect 620 101 625 103
rect 630 138 635 140
rect 630 136 632 138
rect 634 136 635 138
rect 630 134 635 136
rect 630 122 634 134
rect 693 138 715 139
rect 693 136 710 138
rect 712 136 715 138
rect 693 135 715 136
rect 678 130 682 132
rect 678 128 679 130
rect 681 128 682 130
rect 630 120 631 122
rect 633 120 634 122
rect 630 112 634 120
rect 630 110 635 112
rect 630 108 632 110
rect 634 108 635 110
rect 630 103 635 108
rect 658 122 666 124
rect 678 123 682 128
rect 711 130 715 135
rect 711 128 712 130
rect 714 128 715 130
rect 658 120 659 122
rect 661 120 666 122
rect 658 118 666 120
rect 676 122 691 123
rect 676 120 678 122
rect 680 120 685 122
rect 687 120 691 122
rect 676 119 691 120
rect 661 115 666 118
rect 661 114 699 115
rect 661 112 663 114
rect 665 112 699 114
rect 661 111 699 112
rect 711 115 715 128
rect 709 113 715 115
rect 709 111 710 113
rect 712 111 715 113
rect 709 106 715 111
rect 709 104 710 106
rect 712 104 715 106
rect 630 101 632 103
rect 634 101 635 103
rect 630 99 635 101
rect 709 102 715 104
rect 719 138 724 140
rect 719 136 721 138
rect 723 136 724 138
rect 719 134 724 136
rect 719 112 723 134
rect 782 138 804 139
rect 782 136 799 138
rect 801 136 804 138
rect 782 135 804 136
rect 719 110 724 112
rect 719 108 721 110
rect 723 108 724 110
rect 719 103 724 108
rect 747 122 755 124
rect 767 123 771 132
rect 747 120 748 122
rect 750 120 751 122
rect 753 120 755 122
rect 747 118 755 120
rect 765 122 780 123
rect 765 120 767 122
rect 769 120 771 122
rect 773 120 774 122
rect 776 120 780 122
rect 765 119 780 120
rect 750 115 755 118
rect 750 111 788 115
rect 800 116 804 135
rect 800 115 801 116
rect 798 114 801 115
rect 803 114 804 116
rect 798 113 804 114
rect 798 111 799 113
rect 801 111 804 113
rect 798 106 804 111
rect 798 104 799 106
rect 801 104 804 106
rect 719 101 721 103
rect 723 101 724 103
rect 719 99 724 101
rect 798 102 804 104
rect 808 138 813 140
rect 808 136 810 138
rect 812 136 813 138
rect 808 131 813 136
rect 808 129 810 131
rect 812 129 813 131
rect 808 127 813 129
rect 808 104 812 127
rect 824 122 836 124
rect 824 120 827 122
rect 829 120 836 122
rect 824 118 836 120
rect 824 115 828 118
rect 824 113 825 115
rect 827 113 828 115
rect 824 110 828 113
rect 840 122 844 124
rect 842 120 844 122
rect 840 117 844 120
rect 840 115 841 117
rect 843 115 844 117
rect 840 108 844 115
rect 808 102 810 104
rect 808 100 812 102
rect 630 95 643 99
rect 719 98 732 99
rect 719 96 721 98
rect 723 96 732 98
rect 719 95 732 96
rect 808 98 820 100
rect 808 97 813 98
rect 808 95 810 97
rect 812 96 813 97
rect 815 96 820 98
rect 812 95 820 96
rect 808 94 820 95
rect 832 102 844 108
rect 9 88 848 89
rect 853 88 857 217
rect 9 86 44 88
rect 46 86 84 88
rect 86 86 286 88
rect 288 86 352 88
rect 354 86 554 88
rect 556 86 620 88
rect 622 86 821 88
rect 823 86 857 88
rect 9 76 857 86
rect 9 74 44 76
rect 46 74 84 76
rect 86 74 286 76
rect 288 74 352 76
rect 354 74 554 76
rect 556 74 620 76
rect 622 74 821 76
rect 823 74 857 76
rect 9 73 857 74
rect 13 59 17 60
rect 13 57 14 59
rect 16 57 17 59
rect 13 51 17 57
rect 44 59 49 61
rect 13 50 26 51
rect 13 48 18 50
rect 20 48 26 50
rect 13 47 26 48
rect 20 42 34 43
rect 20 40 28 42
rect 30 40 34 42
rect 20 39 34 40
rect 44 57 45 59
rect 47 57 49 59
rect 44 52 49 57
rect 44 50 45 52
rect 47 50 49 52
rect 44 48 49 50
rect 20 33 25 39
rect 20 31 22 33
rect 24 31 25 33
rect 20 30 25 31
rect 45 34 49 48
rect 53 51 57 60
rect 95 63 108 67
rect 184 66 197 67
rect 184 64 186 66
rect 188 64 197 66
rect 184 63 197 64
rect 273 67 285 68
rect 273 65 275 67
rect 277 66 285 67
rect 277 65 278 66
rect 273 64 278 65
rect 280 64 285 66
rect 95 61 100 63
rect 84 59 89 61
rect 53 50 66 51
rect 53 48 54 50
rect 56 48 58 50
rect 60 48 66 50
rect 53 47 66 48
rect 45 32 46 34
rect 48 32 49 34
rect 45 28 49 32
rect 60 42 74 43
rect 60 40 62 42
rect 64 40 68 42
rect 70 40 74 42
rect 60 39 74 40
rect 84 57 85 59
rect 87 57 89 59
rect 84 52 89 57
rect 84 50 85 52
rect 87 50 89 52
rect 84 48 89 50
rect 60 30 65 39
rect 85 46 89 48
rect 85 44 86 46
rect 88 44 89 46
rect 37 26 45 28
rect 47 26 49 28
rect 85 28 89 44
rect 37 22 49 26
rect 77 26 85 28
rect 87 26 89 28
rect 77 22 89 26
rect 95 59 97 61
rect 99 59 100 61
rect 184 61 189 63
rect 95 54 100 59
rect 95 52 97 54
rect 99 52 100 54
rect 95 50 100 52
rect 95 42 99 50
rect 95 40 96 42
rect 98 40 99 42
rect 126 50 164 51
rect 126 48 128 50
rect 130 48 164 50
rect 126 47 164 48
rect 95 28 99 40
rect 126 44 131 47
rect 123 42 131 44
rect 123 40 124 42
rect 126 40 131 42
rect 123 38 131 40
rect 141 42 156 43
rect 141 40 143 42
rect 145 40 150 42
rect 152 40 156 42
rect 141 39 156 40
rect 95 26 100 28
rect 143 34 147 39
rect 174 58 180 60
rect 174 56 175 58
rect 177 56 180 58
rect 174 51 180 56
rect 174 49 175 51
rect 177 49 180 51
rect 174 47 180 49
rect 143 32 144 34
rect 146 32 147 34
rect 143 30 147 32
rect 176 34 180 47
rect 176 32 177 34
rect 179 32 180 34
rect 176 27 180 32
rect 95 24 97 26
rect 99 24 100 26
rect 95 22 100 24
rect 158 26 180 27
rect 158 24 175 26
rect 177 24 180 26
rect 158 23 180 24
rect 184 59 186 61
rect 188 59 189 61
rect 273 62 285 64
rect 273 60 277 62
rect 184 54 189 59
rect 184 52 186 54
rect 188 52 189 54
rect 184 50 189 52
rect 184 28 188 50
rect 215 47 253 51
rect 215 44 220 47
rect 212 42 220 44
rect 212 40 213 42
rect 215 40 216 42
rect 218 40 220 42
rect 212 38 220 40
rect 230 42 245 43
rect 230 40 232 42
rect 234 40 236 42
rect 238 40 239 42
rect 241 40 245 42
rect 230 39 245 40
rect 184 26 189 28
rect 232 30 236 39
rect 263 58 269 60
rect 263 56 264 58
rect 266 56 269 58
rect 263 51 269 56
rect 263 49 264 51
rect 266 49 269 51
rect 263 48 269 49
rect 263 47 266 48
rect 265 46 266 47
rect 268 46 269 48
rect 265 27 269 46
rect 184 24 186 26
rect 188 24 189 26
rect 184 22 189 24
rect 247 26 269 27
rect 247 24 264 26
rect 266 24 269 26
rect 247 23 269 24
rect 273 58 275 60
rect 273 35 277 58
rect 297 54 309 60
rect 273 33 278 35
rect 273 31 275 33
rect 277 31 278 33
rect 273 26 278 31
rect 289 49 293 52
rect 289 47 290 49
rect 292 47 293 49
rect 289 44 293 47
rect 289 42 301 44
rect 289 40 292 42
rect 294 40 301 42
rect 289 38 301 40
rect 305 47 309 54
rect 321 59 325 60
rect 321 57 322 59
rect 324 57 325 59
rect 321 51 325 57
rect 363 63 376 67
rect 452 66 465 67
rect 452 64 454 66
rect 456 64 465 66
rect 452 63 465 64
rect 541 67 553 68
rect 541 65 543 67
rect 545 66 553 67
rect 545 65 546 66
rect 541 64 546 65
rect 548 64 553 66
rect 363 61 368 63
rect 352 59 357 61
rect 321 50 334 51
rect 321 48 326 50
rect 328 48 334 50
rect 321 47 334 48
rect 305 45 306 47
rect 308 45 309 47
rect 305 42 309 45
rect 307 40 309 42
rect 305 38 309 40
rect 328 42 342 43
rect 328 40 336 42
rect 338 40 339 42
rect 341 40 342 42
rect 328 39 342 40
rect 352 57 353 59
rect 355 57 357 59
rect 352 52 357 57
rect 352 50 353 52
rect 355 50 357 52
rect 352 48 357 50
rect 328 30 333 39
rect 353 34 357 48
rect 353 32 354 34
rect 356 32 357 34
rect 273 24 275 26
rect 277 24 278 26
rect 273 22 278 24
rect 353 28 357 32
rect 345 26 353 28
rect 355 26 357 28
rect 345 22 357 26
rect 363 59 365 61
rect 367 59 368 61
rect 452 61 457 63
rect 363 54 368 59
rect 363 52 365 54
rect 367 52 368 54
rect 363 50 368 52
rect 363 42 367 50
rect 363 40 364 42
rect 366 40 367 42
rect 394 50 432 51
rect 394 48 396 50
rect 398 48 432 50
rect 394 47 432 48
rect 363 28 367 40
rect 394 44 399 47
rect 391 42 399 44
rect 391 40 392 42
rect 394 40 399 42
rect 391 38 399 40
rect 409 42 424 43
rect 409 40 411 42
rect 413 40 418 42
rect 420 40 424 42
rect 409 39 424 40
rect 363 26 368 28
rect 411 34 415 39
rect 442 58 448 60
rect 442 56 443 58
rect 445 56 448 58
rect 442 51 448 56
rect 442 49 443 51
rect 445 49 448 51
rect 442 47 448 49
rect 411 32 412 34
rect 414 32 415 34
rect 411 30 415 32
rect 444 34 448 47
rect 444 32 445 34
rect 447 32 448 34
rect 444 27 448 32
rect 363 24 365 26
rect 367 24 368 26
rect 363 22 368 24
rect 426 26 448 27
rect 426 24 443 26
rect 445 24 448 26
rect 426 23 448 24
rect 452 59 454 61
rect 456 59 457 61
rect 541 62 553 64
rect 541 60 545 62
rect 452 54 457 59
rect 452 52 454 54
rect 456 52 457 54
rect 452 50 457 52
rect 452 28 456 50
rect 483 47 521 51
rect 483 44 488 47
rect 480 42 488 44
rect 480 40 481 42
rect 483 40 484 42
rect 486 40 488 42
rect 480 38 488 40
rect 498 42 513 43
rect 498 40 500 42
rect 502 40 504 42
rect 506 40 507 42
rect 509 40 513 42
rect 498 39 513 40
rect 452 26 457 28
rect 500 30 504 39
rect 531 58 537 60
rect 531 56 532 58
rect 534 56 537 58
rect 531 51 537 56
rect 531 49 532 51
rect 534 49 537 51
rect 531 48 537 49
rect 531 47 534 48
rect 533 46 534 47
rect 536 46 537 48
rect 533 27 537 46
rect 452 24 454 26
rect 456 24 457 26
rect 452 22 457 24
rect 515 26 537 27
rect 515 24 532 26
rect 534 24 537 26
rect 515 23 537 24
rect 541 58 543 60
rect 541 35 545 58
rect 565 54 577 60
rect 541 33 546 35
rect 541 31 543 33
rect 545 31 546 33
rect 541 26 546 31
rect 557 49 561 52
rect 557 47 558 49
rect 560 47 561 49
rect 557 44 561 47
rect 557 42 569 44
rect 557 40 560 42
rect 562 40 569 42
rect 557 38 569 40
rect 573 47 577 54
rect 589 59 593 60
rect 589 57 590 59
rect 592 57 593 59
rect 589 51 593 57
rect 630 63 643 67
rect 719 66 732 67
rect 719 64 721 66
rect 723 64 732 66
rect 719 63 732 64
rect 808 67 820 68
rect 808 65 810 67
rect 812 66 820 67
rect 812 65 813 66
rect 808 64 813 65
rect 815 64 820 66
rect 630 61 635 63
rect 620 59 625 61
rect 589 50 602 51
rect 589 48 594 50
rect 596 48 602 50
rect 589 47 602 48
rect 573 45 574 47
rect 576 45 577 47
rect 573 42 577 45
rect 575 40 577 42
rect 573 38 577 40
rect 596 42 610 43
rect 596 40 604 42
rect 606 40 607 42
rect 609 40 610 42
rect 596 39 610 40
rect 620 57 621 59
rect 623 57 625 59
rect 620 52 625 57
rect 620 50 621 52
rect 623 50 625 52
rect 620 48 625 50
rect 596 30 601 39
rect 621 34 625 48
rect 621 32 622 34
rect 624 32 625 34
rect 541 24 543 26
rect 545 24 546 26
rect 541 22 546 24
rect 621 28 625 32
rect 613 26 621 28
rect 623 26 625 28
rect 613 22 625 26
rect 630 59 632 61
rect 634 59 635 61
rect 719 61 724 63
rect 630 54 635 59
rect 630 52 632 54
rect 634 52 635 54
rect 630 50 635 52
rect 630 42 634 50
rect 630 40 631 42
rect 633 40 634 42
rect 661 50 699 51
rect 661 48 663 50
rect 665 48 699 50
rect 661 47 699 48
rect 630 28 634 40
rect 661 44 666 47
rect 658 42 666 44
rect 658 40 659 42
rect 661 40 666 42
rect 658 38 666 40
rect 676 42 691 43
rect 676 40 678 42
rect 680 40 685 42
rect 687 40 691 42
rect 676 39 691 40
rect 630 26 635 28
rect 678 34 682 39
rect 709 58 715 60
rect 709 56 710 58
rect 712 56 715 58
rect 709 51 715 56
rect 709 49 710 51
rect 712 49 715 51
rect 709 47 715 49
rect 678 32 679 34
rect 681 32 682 34
rect 678 30 682 32
rect 711 34 715 47
rect 711 32 712 34
rect 714 32 715 34
rect 711 27 715 32
rect 630 24 632 26
rect 634 24 635 26
rect 630 22 635 24
rect 693 26 715 27
rect 693 24 710 26
rect 712 24 715 26
rect 693 23 715 24
rect 719 59 721 61
rect 723 59 724 61
rect 808 62 820 64
rect 808 60 812 62
rect 719 54 724 59
rect 719 52 721 54
rect 723 52 724 54
rect 719 50 724 52
rect 719 28 723 50
rect 750 47 788 51
rect 750 44 755 47
rect 747 42 755 44
rect 747 40 748 42
rect 750 40 751 42
rect 753 40 755 42
rect 747 38 755 40
rect 765 42 780 43
rect 765 40 767 42
rect 769 40 771 42
rect 773 40 774 42
rect 776 40 780 42
rect 765 39 780 40
rect 719 26 724 28
rect 767 30 771 39
rect 798 58 804 60
rect 798 56 799 58
rect 801 56 804 58
rect 798 51 804 56
rect 798 49 799 51
rect 801 49 804 51
rect 798 48 804 49
rect 798 47 801 48
rect 800 46 801 47
rect 803 46 804 48
rect 800 27 804 46
rect 719 24 721 26
rect 723 24 724 26
rect 719 22 724 24
rect 782 26 804 27
rect 782 24 799 26
rect 801 24 804 26
rect 782 23 804 24
rect 808 58 810 60
rect 808 35 812 58
rect 832 54 844 60
rect 808 33 813 35
rect 808 31 810 33
rect 812 31 813 33
rect 808 26 813 31
rect 824 49 828 52
rect 824 47 825 49
rect 827 47 828 49
rect 824 44 828 47
rect 824 42 836 44
rect 824 40 827 42
rect 829 40 836 42
rect 824 38 836 40
rect 840 47 844 54
rect 840 45 841 47
rect 843 45 844 47
rect 840 42 844 45
rect 842 40 844 42
rect 840 38 844 40
rect 808 24 810 26
rect 812 24 813 26
rect 808 22 813 24
rect 0 16 848 17
rect 0 14 34 16
rect 36 14 44 16
rect 46 14 74 16
rect 76 14 84 16
rect 86 14 302 16
rect 304 15 342 16
rect 304 14 308 15
rect 0 13 308 14
rect 310 14 342 15
rect 344 14 352 16
rect 354 14 570 16
rect 572 15 610 16
rect 572 14 576 15
rect 310 13 576 14
rect 578 14 610 15
rect 612 14 620 16
rect 622 14 837 16
rect 839 15 848 16
rect 839 14 843 15
rect 578 13 843 14
rect 845 13 848 15
rect 0 9 848 13
rect 3 3 852 4
rect 3 1 12 3
rect 14 1 57 3
rect 59 1 330 3
rect 332 1 595 3
rect 597 1 852 3
rect 3 0 852 1
<< alu2 >>
rect 20 305 28 306
rect 20 303 21 305
rect 23 303 25 305
rect 27 303 28 305
rect 20 302 28 303
rect 58 305 66 306
rect 58 303 59 305
rect 61 303 63 305
rect 65 303 66 305
rect 58 302 66 303
rect 317 305 325 306
rect 317 303 318 305
rect 320 303 322 305
rect 324 303 325 305
rect 317 302 325 303
rect 594 305 602 306
rect 594 303 595 305
rect 597 303 599 305
rect 601 303 602 305
rect 594 302 602 303
rect 11 300 16 301
rect 11 298 12 300
rect 14 298 16 300
rect 11 297 16 298
rect 32 297 54 301
rect 70 300 313 301
rect 70 298 306 300
rect 308 298 313 300
rect 70 297 313 298
rect 329 297 590 301
rect 606 300 838 301
rect 606 298 614 300
rect 616 298 838 300
rect 606 297 838 298
rect 11 293 36 297
rect 50 293 74 297
rect 309 293 333 297
rect 586 293 610 297
rect 5 275 25 276
rect 5 273 22 275
rect 24 273 25 275
rect 5 271 25 273
rect 5 204 9 271
rect 31 259 36 293
rect 143 292 147 293
rect 143 290 144 292
rect 146 290 147 292
rect 85 275 89 288
rect 45 274 89 275
rect 45 272 46 274
rect 48 272 89 274
rect 45 271 89 272
rect 143 274 147 290
rect 328 275 333 276
rect 589 275 601 276
rect 143 272 144 274
rect 146 272 147 274
rect 143 271 147 272
rect 176 274 309 275
rect 176 272 177 274
rect 179 272 309 274
rect 176 271 309 272
rect 49 266 65 267
rect 49 264 50 266
rect 52 264 62 266
rect 64 264 65 266
rect 49 263 65 264
rect 95 266 219 267
rect 95 264 96 266
rect 98 264 216 266
rect 218 264 219 266
rect 95 263 219 264
rect 235 266 239 267
rect 235 264 236 266
rect 238 264 239 266
rect 85 262 89 263
rect 85 260 86 262
rect 88 260 89 262
rect 85 259 89 260
rect 31 255 49 259
rect 53 258 66 259
rect 53 256 54 258
rect 56 256 63 258
rect 65 256 66 258
rect 53 255 66 256
rect 85 258 131 259
rect 85 256 128 258
rect 130 256 131 258
rect 85 255 131 256
rect 13 249 36 250
rect 13 247 14 249
rect 16 247 36 249
rect 13 246 36 247
rect 5 203 17 204
rect 5 201 14 203
rect 16 201 17 203
rect 5 200 17 201
rect 5 132 9 200
rect 20 185 25 187
rect 20 183 21 185
rect 23 183 25 185
rect 20 177 25 183
rect 20 175 22 177
rect 24 175 25 177
rect 20 174 25 175
rect 5 131 25 132
rect 5 129 22 131
rect 24 129 25 131
rect 5 127 25 129
rect 5 60 9 127
rect 14 114 24 115
rect 14 112 15 114
rect 17 112 21 114
rect 23 112 24 114
rect 14 111 24 112
rect 5 59 17 60
rect 5 57 14 59
rect 16 57 17 59
rect 5 56 17 57
rect 32 43 36 246
rect 44 226 49 255
rect 235 244 239 264
rect 305 261 309 271
rect 328 273 330 275
rect 332 273 333 275
rect 328 267 333 273
rect 353 274 415 275
rect 353 272 354 274
rect 356 272 412 274
rect 414 272 415 274
rect 353 271 415 272
rect 444 274 577 275
rect 444 272 445 274
rect 447 272 577 274
rect 444 271 577 272
rect 589 274 598 275
rect 589 272 590 274
rect 592 273 598 274
rect 600 273 601 275
rect 592 272 601 273
rect 589 271 601 272
rect 621 274 682 275
rect 621 272 622 274
rect 624 272 679 274
rect 681 272 682 274
rect 621 271 682 272
rect 711 274 844 275
rect 711 272 712 274
rect 714 272 844 274
rect 711 271 844 272
rect 328 266 342 267
rect 328 264 331 266
rect 333 264 342 266
rect 328 263 342 264
rect 363 266 487 267
rect 363 264 364 266
rect 366 264 484 266
rect 486 264 487 266
rect 363 263 487 264
rect 503 266 507 267
rect 503 264 504 266
rect 506 264 507 266
rect 265 260 293 261
rect 265 258 266 260
rect 268 259 293 260
rect 268 258 290 259
rect 265 257 290 258
rect 292 257 293 259
rect 265 256 293 257
rect 305 259 306 261
rect 308 259 309 261
rect 305 256 309 259
rect 352 258 399 259
rect 352 256 396 258
rect 398 256 399 258
rect 321 254 325 256
rect 321 252 322 254
rect 324 252 325 254
rect 321 250 325 252
rect 321 248 322 250
rect 324 248 325 250
rect 321 247 325 248
rect 352 255 399 256
rect 185 242 189 243
rect 185 240 186 242
rect 188 240 189 242
rect 185 231 189 240
rect 235 242 236 244
rect 238 242 239 244
rect 352 243 356 255
rect 503 244 507 264
rect 573 261 577 271
rect 630 266 754 267
rect 630 264 631 266
rect 633 264 751 266
rect 753 264 754 266
rect 630 263 754 264
rect 770 266 774 267
rect 770 264 771 266
rect 773 264 774 266
rect 533 260 561 261
rect 533 258 534 260
rect 536 259 561 260
rect 536 258 558 259
rect 533 257 558 258
rect 560 257 561 259
rect 533 256 561 257
rect 573 259 574 261
rect 576 259 577 261
rect 573 256 577 259
rect 589 258 602 259
rect 589 256 590 258
rect 592 256 599 258
rect 601 256 602 258
rect 589 255 602 256
rect 631 258 666 259
rect 631 256 663 258
rect 665 256 666 258
rect 631 255 666 256
rect 235 235 239 242
rect 275 242 356 243
rect 275 240 278 242
rect 280 240 356 242
rect 275 238 356 240
rect 453 242 457 243
rect 453 240 454 242
rect 456 240 457 242
rect 453 231 457 240
rect 503 242 504 244
rect 506 242 507 244
rect 631 242 635 255
rect 770 244 774 264
rect 840 261 844 271
rect 800 260 828 261
rect 800 258 801 260
rect 803 259 828 260
rect 803 258 825 259
rect 800 257 825 258
rect 827 257 828 259
rect 800 256 828 257
rect 840 259 841 261
rect 843 259 844 261
rect 840 256 844 259
rect 503 235 507 242
rect 543 241 635 242
rect 543 239 546 241
rect 548 239 635 241
rect 543 238 635 239
rect 720 242 724 243
rect 720 240 721 242
rect 723 240 724 242
rect 720 231 724 240
rect 770 242 771 244
rect 773 242 774 244
rect 770 235 774 242
rect 810 242 854 243
rect 810 240 813 242
rect 815 240 854 242
rect 810 238 854 240
rect 185 227 356 231
rect 453 227 636 231
rect 720 227 859 231
rect 44 222 74 226
rect 49 194 57 195
rect 49 192 50 194
rect 52 192 54 194
rect 56 192 57 194
rect 49 191 57 192
rect 70 187 74 222
rect 185 219 346 223
rect 185 210 189 219
rect 185 208 186 210
rect 188 208 189 210
rect 185 207 189 208
rect 235 202 239 215
rect 275 210 317 212
rect 275 208 278 210
rect 280 208 312 210
rect 314 208 317 210
rect 275 207 317 208
rect 321 203 325 204
rect 235 198 317 202
rect 85 194 131 195
rect 85 192 128 194
rect 130 192 131 194
rect 85 191 131 192
rect 85 190 89 191
rect 85 188 86 190
rect 88 188 89 190
rect 85 187 89 188
rect 60 186 74 187
rect 60 184 62 186
rect 64 184 74 186
rect 60 183 74 184
rect 95 186 219 187
rect 95 184 96 186
rect 98 184 216 186
rect 218 184 219 186
rect 95 183 219 184
rect 235 186 239 198
rect 265 193 293 194
rect 265 192 290 193
rect 265 190 266 192
rect 268 191 290 192
rect 292 191 293 193
rect 268 190 293 191
rect 265 189 293 190
rect 305 191 309 194
rect 305 189 306 191
rect 308 189 309 191
rect 235 184 236 186
rect 238 184 239 186
rect 235 183 239 184
rect 305 179 309 189
rect 45 178 147 179
rect 45 176 46 178
rect 48 176 144 178
rect 146 176 147 178
rect 45 175 147 176
rect 176 178 309 179
rect 176 176 177 178
rect 179 176 309 178
rect 176 175 309 176
rect 45 130 147 131
rect 45 128 46 130
rect 48 128 144 130
rect 146 128 147 130
rect 45 127 147 128
rect 176 130 309 131
rect 176 128 177 130
rect 179 128 309 130
rect 176 127 309 128
rect 49 122 65 123
rect 49 120 50 122
rect 52 120 62 122
rect 64 120 65 122
rect 49 119 65 120
rect 95 122 219 123
rect 95 120 96 122
rect 98 120 216 122
rect 218 120 219 122
rect 95 119 219 120
rect 235 122 239 123
rect 235 120 236 122
rect 238 120 239 122
rect 85 118 89 119
rect 85 116 86 118
rect 88 116 89 118
rect 85 115 89 116
rect 53 114 66 115
rect 53 112 54 114
rect 56 112 61 114
rect 63 112 66 114
rect 53 111 66 112
rect 85 114 131 115
rect 85 112 128 114
rect 130 112 131 114
rect 85 111 131 112
rect 235 99 239 120
rect 305 117 309 127
rect 265 116 293 117
rect 265 114 266 116
rect 268 115 293 116
rect 268 114 290 115
rect 265 113 290 114
rect 292 113 293 115
rect 265 112 293 113
rect 305 115 306 117
rect 308 115 309 117
rect 305 112 309 115
rect 313 99 317 198
rect 321 201 322 203
rect 324 201 325 203
rect 321 195 325 201
rect 321 194 334 195
rect 321 192 331 194
rect 333 192 334 194
rect 321 191 334 192
rect 321 178 333 179
rect 321 176 322 178
rect 324 177 333 178
rect 324 176 330 177
rect 321 175 330 176
rect 332 175 333 177
rect 321 174 333 175
rect 328 130 333 132
rect 328 128 329 130
rect 331 128 333 130
rect 328 123 333 128
rect 328 122 335 123
rect 328 120 331 122
rect 333 120 335 122
rect 328 119 335 120
rect 342 115 346 219
rect 352 195 356 227
rect 453 219 611 223
rect 453 210 457 219
rect 453 208 454 210
rect 456 208 457 210
rect 453 207 457 208
rect 503 202 507 215
rect 543 210 583 212
rect 543 208 546 210
rect 548 208 580 210
rect 582 208 583 210
rect 543 207 583 208
rect 589 203 593 204
rect 503 198 585 202
rect 352 194 399 195
rect 352 192 396 194
rect 398 192 399 194
rect 352 191 399 192
rect 363 186 487 187
rect 363 184 364 186
rect 366 184 484 186
rect 486 184 487 186
rect 363 183 487 184
rect 503 186 507 198
rect 533 193 561 194
rect 533 192 558 193
rect 533 190 534 192
rect 536 191 558 192
rect 560 191 561 193
rect 536 190 561 191
rect 533 189 561 190
rect 573 191 577 194
rect 573 189 574 191
rect 576 189 577 191
rect 503 184 504 186
rect 506 184 507 186
rect 503 183 507 184
rect 573 179 577 189
rect 353 178 415 179
rect 353 176 354 178
rect 356 176 412 178
rect 414 176 415 178
rect 353 175 415 176
rect 444 178 577 179
rect 444 176 445 178
rect 447 176 577 178
rect 444 175 577 176
rect 353 130 415 131
rect 353 128 354 130
rect 356 128 412 130
rect 414 128 415 130
rect 353 127 415 128
rect 444 130 577 131
rect 444 128 445 130
rect 447 128 577 130
rect 444 127 577 128
rect 363 122 487 123
rect 363 120 364 122
rect 366 120 484 122
rect 486 120 487 122
rect 363 119 487 120
rect 503 122 507 123
rect 503 120 504 122
rect 506 120 507 122
rect 342 114 399 115
rect 321 111 325 113
rect 321 109 322 111
rect 324 109 325 111
rect 342 112 396 114
rect 398 112 399 114
rect 342 111 399 112
rect 342 110 346 111
rect 321 105 325 109
rect 321 103 322 105
rect 324 103 325 105
rect 321 102 325 103
rect 503 99 507 120
rect 573 117 577 127
rect 533 116 561 117
rect 533 114 534 116
rect 536 115 561 116
rect 536 114 558 115
rect 533 113 558 114
rect 560 113 561 115
rect 533 112 561 113
rect 573 115 574 117
rect 576 115 577 117
rect 573 112 577 115
rect 581 99 585 198
rect 589 201 590 203
rect 592 201 593 203
rect 589 195 593 201
rect 589 193 590 195
rect 592 193 593 195
rect 589 191 593 193
rect 596 186 601 187
rect 596 184 598 186
rect 600 184 601 186
rect 596 179 601 184
rect 589 177 601 179
rect 589 175 598 177
rect 600 175 601 177
rect 589 174 601 175
rect 589 131 601 132
rect 589 129 590 131
rect 592 129 598 131
rect 600 129 601 131
rect 589 127 601 129
rect 607 115 611 219
rect 630 195 636 227
rect 720 219 859 223
rect 720 210 724 219
rect 720 208 721 210
rect 723 208 724 210
rect 720 207 724 208
rect 770 202 774 215
rect 810 210 855 212
rect 810 208 813 210
rect 815 208 847 210
rect 849 208 855 210
rect 810 207 855 208
rect 770 198 852 202
rect 630 194 666 195
rect 630 192 663 194
rect 665 192 666 194
rect 630 191 666 192
rect 630 186 754 187
rect 630 184 631 186
rect 633 184 751 186
rect 753 184 754 186
rect 630 183 754 184
rect 770 186 774 198
rect 800 193 828 194
rect 800 192 825 193
rect 800 190 801 192
rect 803 191 825 192
rect 827 191 828 193
rect 803 190 828 191
rect 800 189 828 190
rect 840 191 844 194
rect 840 189 841 191
rect 843 189 844 191
rect 770 184 771 186
rect 773 184 774 186
rect 770 183 774 184
rect 840 179 844 189
rect 621 178 682 179
rect 621 176 622 178
rect 624 176 679 178
rect 681 176 682 178
rect 621 175 682 176
rect 711 178 844 179
rect 711 176 712 178
rect 714 176 844 178
rect 711 175 844 176
rect 621 130 682 131
rect 621 128 622 130
rect 624 128 679 130
rect 681 128 682 130
rect 621 127 682 128
rect 711 130 844 131
rect 711 128 712 130
rect 714 128 844 130
rect 711 127 844 128
rect 630 122 754 123
rect 630 120 631 122
rect 633 120 751 122
rect 753 120 754 122
rect 630 119 754 120
rect 770 122 774 123
rect 770 120 771 122
rect 773 120 774 122
rect 589 114 602 115
rect 589 112 599 114
rect 601 112 602 114
rect 589 111 602 112
rect 607 114 666 115
rect 607 112 663 114
rect 665 112 666 114
rect 607 111 666 112
rect 589 105 593 111
rect 607 110 611 111
rect 589 103 590 105
rect 592 103 593 105
rect 589 102 593 103
rect 770 99 774 120
rect 840 117 844 127
rect 800 116 828 117
rect 800 114 801 116
rect 803 115 828 116
rect 803 114 825 115
rect 800 113 825 114
rect 827 113 828 115
rect 800 112 828 113
rect 840 115 841 117
rect 843 115 844 117
rect 840 112 844 115
rect 848 99 852 198
rect 185 98 189 99
rect 185 96 186 98
rect 188 96 189 98
rect 185 87 189 96
rect 235 97 236 99
rect 238 97 239 99
rect 235 91 239 97
rect 275 98 317 99
rect 275 96 278 98
rect 280 96 317 98
rect 275 94 317 96
rect 453 98 457 99
rect 453 96 454 98
rect 456 96 457 98
rect 453 87 457 96
rect 503 97 504 99
rect 506 97 507 99
rect 503 91 507 97
rect 543 98 585 99
rect 543 96 546 98
rect 548 96 585 98
rect 543 94 585 96
rect 720 98 724 99
rect 720 96 721 98
rect 723 96 724 98
rect 720 87 724 96
rect 770 97 771 99
rect 773 97 774 99
rect 770 91 774 97
rect 810 98 852 99
rect 810 96 813 98
rect 815 96 852 98
rect 810 94 852 96
rect 185 83 361 87
rect 453 83 637 87
rect 720 83 859 87
rect 185 75 317 79
rect 185 66 189 75
rect 185 64 186 66
rect 188 64 189 66
rect 185 63 189 64
rect 235 59 239 71
rect 275 66 313 68
rect 275 64 278 66
rect 280 64 310 66
rect 312 64 313 66
rect 275 63 313 64
rect 321 59 325 60
rect 235 54 317 59
rect 49 50 57 51
rect 49 48 50 50
rect 52 48 54 50
rect 56 48 57 50
rect 49 47 57 48
rect 85 50 131 51
rect 85 48 128 50
rect 130 48 131 50
rect 85 47 131 48
rect 85 46 89 47
rect 85 44 86 46
rect 88 44 89 46
rect 85 43 89 44
rect 32 42 65 43
rect 32 40 62 42
rect 64 40 65 42
rect 32 39 65 40
rect 95 42 219 43
rect 95 40 96 42
rect 98 40 216 42
rect 218 40 219 42
rect 95 39 219 40
rect 235 42 239 54
rect 265 49 293 50
rect 265 48 290 49
rect 265 46 266 48
rect 268 47 290 48
rect 292 47 293 49
rect 268 46 293 47
rect 265 45 293 46
rect 305 47 309 50
rect 305 45 306 47
rect 308 45 309 47
rect 235 40 236 42
rect 238 40 239 42
rect 235 39 239 40
rect 16 33 25 35
rect 16 31 17 33
rect 19 31 22 33
rect 24 31 25 33
rect 16 30 25 31
rect 3 9 28 13
rect 3 4 7 9
rect 24 8 28 9
rect 32 8 36 39
rect 305 35 309 45
rect 45 34 147 35
rect 45 32 46 34
rect 48 32 144 34
rect 146 32 147 34
rect 45 31 147 32
rect 176 34 309 35
rect 176 32 177 34
rect 179 32 309 34
rect 176 31 309 32
rect 313 27 317 54
rect 321 57 322 59
rect 324 57 325 59
rect 321 51 325 57
rect 356 51 361 83
rect 453 75 585 79
rect 453 66 457 75
rect 453 64 454 66
rect 456 64 457 66
rect 453 63 457 64
rect 503 59 507 71
rect 543 66 581 68
rect 543 64 546 66
rect 548 64 578 66
rect 580 64 581 66
rect 543 63 581 64
rect 589 59 593 60
rect 503 54 585 59
rect 321 50 334 51
rect 321 48 331 50
rect 333 48 334 50
rect 321 47 334 48
rect 356 50 399 51
rect 356 48 396 50
rect 398 48 399 50
rect 356 47 399 48
rect 306 23 317 27
rect 338 42 342 43
rect 338 40 339 42
rect 341 40 342 42
rect 306 15 311 23
rect 306 13 308 15
rect 310 13 311 15
rect 48 8 72 13
rect 306 12 311 13
rect 338 12 342 40
rect 363 42 487 43
rect 363 40 364 42
rect 366 40 484 42
rect 486 40 487 42
rect 363 39 487 40
rect 503 42 507 54
rect 533 49 561 50
rect 533 48 558 49
rect 533 46 534 48
rect 536 47 558 48
rect 560 47 561 49
rect 536 46 561 47
rect 533 45 561 46
rect 573 47 577 50
rect 573 45 574 47
rect 576 45 577 47
rect 503 40 504 42
rect 506 40 507 42
rect 503 39 507 40
rect 573 35 577 45
rect 353 34 415 35
rect 353 32 354 34
rect 356 32 412 34
rect 414 32 415 34
rect 353 31 415 32
rect 444 34 577 35
rect 444 32 445 34
rect 447 32 577 34
rect 444 31 577 32
rect 581 21 585 54
rect 589 57 590 59
rect 592 57 593 59
rect 589 50 593 57
rect 589 48 590 50
rect 592 48 593 50
rect 589 47 593 48
rect 630 51 637 83
rect 720 75 859 79
rect 720 66 724 75
rect 720 64 721 66
rect 723 64 724 66
rect 720 63 724 64
rect 770 59 774 71
rect 810 66 855 68
rect 810 64 813 66
rect 815 64 845 66
rect 847 64 855 66
rect 810 63 855 64
rect 770 54 852 59
rect 630 50 666 51
rect 630 48 663 50
rect 665 48 666 50
rect 630 47 666 48
rect 575 17 585 21
rect 606 42 610 43
rect 606 40 607 42
rect 609 40 610 42
rect 574 15 579 17
rect 574 13 576 15
rect 578 13 579 15
rect 574 12 579 13
rect 606 12 610 40
rect 630 42 754 43
rect 630 40 631 42
rect 633 40 751 42
rect 753 40 754 42
rect 630 39 754 40
rect 770 42 774 54
rect 800 49 828 50
rect 800 48 825 49
rect 800 46 801 48
rect 803 47 825 48
rect 827 47 828 49
rect 803 46 828 47
rect 800 45 828 46
rect 840 47 844 50
rect 840 45 841 47
rect 843 45 844 47
rect 770 40 771 42
rect 773 40 774 42
rect 770 39 774 40
rect 840 35 844 45
rect 621 34 682 35
rect 621 32 622 34
rect 624 32 679 34
rect 681 32 682 34
rect 621 31 682 32
rect 711 34 844 35
rect 711 32 712 34
rect 714 32 844 34
rect 711 31 844 32
rect 848 17 852 54
rect 841 15 852 17
rect 841 13 843 15
rect 845 13 852 15
rect 841 12 852 13
rect 317 8 342 12
rect 586 8 610 12
rect 24 4 52 8
rect 68 4 321 8
rect 337 4 590 8
rect 606 4 852 8
rect 11 3 20 4
rect 11 1 12 3
rect 14 1 17 3
rect 19 1 20 3
rect 11 0 20 1
rect 56 3 64 4
rect 56 1 57 3
rect 59 1 61 3
rect 63 1 64 3
rect 56 0 64 1
rect 325 3 333 4
rect 325 1 326 3
rect 328 1 330 3
rect 332 1 333 3
rect 325 0 333 1
rect 594 3 602 4
rect 594 1 595 3
rect 597 1 599 3
rect 601 1 602 3
rect 594 0 602 1
<< alu3 >>
rect 20 305 24 306
rect 20 303 21 305
rect 23 303 24 305
rect 11 300 15 301
rect 11 298 12 300
rect 14 298 15 300
rect 11 115 15 298
rect 20 185 24 303
rect 62 305 66 306
rect 62 303 63 305
rect 65 303 66 305
rect 20 183 21 185
rect 23 183 24 185
rect 20 181 24 183
rect 49 266 53 298
rect 49 264 50 266
rect 52 264 53 266
rect 49 194 53 264
rect 62 258 66 303
rect 321 305 325 306
rect 321 303 322 305
rect 324 303 325 305
rect 302 300 316 301
rect 302 298 306 300
rect 308 298 316 300
rect 302 297 316 298
rect 62 256 63 258
rect 65 256 66 258
rect 62 255 66 256
rect 235 244 239 245
rect 235 242 236 244
rect 238 242 239 244
rect 235 217 239 242
rect 311 237 316 297
rect 321 254 325 303
rect 598 305 602 306
rect 598 303 599 305
rect 601 303 602 305
rect 321 252 322 254
rect 324 252 325 254
rect 321 251 325 252
rect 330 266 334 298
rect 330 264 331 266
rect 333 264 334 266
rect 311 232 326 237
rect 235 213 315 217
rect 311 210 315 213
rect 311 208 312 210
rect 314 208 315 210
rect 311 207 315 208
rect 49 192 50 194
rect 52 192 53 194
rect 49 122 53 192
rect 321 178 326 232
rect 321 176 322 178
rect 324 176 326 178
rect 321 174 326 176
rect 330 194 334 264
rect 589 274 593 299
rect 589 272 590 274
rect 592 272 593 274
rect 503 244 507 245
rect 503 242 504 244
rect 506 242 507 244
rect 503 217 507 242
rect 503 213 583 217
rect 579 210 583 213
rect 579 208 580 210
rect 582 208 583 210
rect 579 207 583 208
rect 330 192 331 194
rect 333 192 334 194
rect 49 120 50 122
rect 52 120 53 122
rect 11 114 20 115
rect 11 112 15 114
rect 17 112 20 114
rect 11 111 20 112
rect 49 50 53 120
rect 330 122 334 192
rect 330 120 331 122
rect 333 120 334 122
rect 49 48 50 50
rect 52 48 53 50
rect 49 35 53 48
rect 60 114 64 115
rect 60 112 61 114
rect 63 112 64 114
rect 16 33 20 35
rect 16 31 17 33
rect 19 31 20 33
rect 16 3 20 31
rect 16 1 17 3
rect 19 1 20 3
rect 16 0 20 1
rect 60 3 64 112
rect 321 111 325 113
rect 321 109 322 111
rect 324 109 325 111
rect 235 99 239 100
rect 235 97 236 99
rect 238 97 239 99
rect 235 73 239 97
rect 235 69 313 73
rect 309 66 313 69
rect 309 64 310 66
rect 312 64 313 66
rect 309 63 313 64
rect 321 13 325 109
rect 330 50 334 120
rect 589 195 593 272
rect 598 258 602 303
rect 598 256 599 258
rect 601 256 602 258
rect 598 255 602 256
rect 613 300 617 301
rect 613 298 614 300
rect 616 298 617 300
rect 613 247 617 298
rect 589 193 590 195
rect 592 193 593 195
rect 589 131 593 193
rect 597 243 617 247
rect 770 244 774 245
rect 597 186 601 243
rect 770 242 771 244
rect 773 242 774 244
rect 770 217 774 242
rect 770 213 850 217
rect 846 210 850 213
rect 846 208 847 210
rect 849 208 850 210
rect 846 207 850 208
rect 597 184 598 186
rect 600 184 601 186
rect 597 179 601 184
rect 589 129 590 131
rect 592 129 593 131
rect 503 99 507 100
rect 503 97 504 99
rect 506 97 507 99
rect 503 73 507 97
rect 503 69 581 73
rect 577 66 581 69
rect 577 64 578 66
rect 580 64 581 66
rect 577 63 581 64
rect 330 48 331 50
rect 333 48 334 50
rect 330 17 334 48
rect 589 50 593 129
rect 589 48 590 50
rect 592 48 593 50
rect 589 17 593 48
rect 598 114 602 115
rect 598 112 599 114
rect 601 112 602 114
rect 321 9 329 13
rect 60 1 61 3
rect 63 1 64 3
rect 60 0 64 1
rect 325 3 329 9
rect 325 1 326 3
rect 328 1 329 3
rect 325 0 329 1
rect 598 3 602 112
rect 770 99 774 100
rect 770 97 771 99
rect 773 97 774 99
rect 770 73 774 97
rect 770 69 848 73
rect 844 66 848 69
rect 844 64 845 66
rect 847 64 848 66
rect 844 63 848 64
rect 598 1 599 3
rect 601 1 602 3
rect 598 0 602 1
<< alu4 >>
rect 48 4 52 12
rect 11 0 20 4
<< ptie >>
rect 42 292 48 294
rect 42 290 44 292
rect 46 290 48 292
rect 42 288 48 290
rect 82 292 88 294
rect 82 290 84 292
rect 86 290 88 292
rect 82 288 88 290
rect 298 292 308 294
rect 298 290 302 292
rect 304 290 308 292
rect 298 288 308 290
rect 350 292 356 294
rect 350 290 352 292
rect 354 290 356 292
rect 350 288 356 290
rect 566 292 576 294
rect 566 290 570 292
rect 572 290 576 292
rect 566 288 576 290
rect 618 292 624 294
rect 618 290 620 292
rect 622 290 624 292
rect 618 288 624 290
rect 833 292 843 294
rect 833 290 837 292
rect 839 290 843 292
rect 833 288 843 290
rect 42 160 48 162
rect 42 158 44 160
rect 46 158 48 160
rect 42 156 48 158
rect 82 160 88 162
rect 82 158 84 160
rect 86 158 88 160
rect 82 156 88 158
rect 298 160 308 162
rect 298 158 302 160
rect 304 158 308 160
rect 298 156 308 158
rect 350 160 356 162
rect 350 158 352 160
rect 354 158 356 160
rect 350 156 356 158
rect 566 160 576 162
rect 566 158 570 160
rect 572 158 576 160
rect 566 156 576 158
rect 618 160 624 162
rect 618 158 620 160
rect 622 158 624 160
rect 618 156 624 158
rect 833 160 843 162
rect 833 158 837 160
rect 839 158 843 160
rect 833 156 843 158
rect 42 148 48 150
rect 42 146 44 148
rect 46 146 48 148
rect 42 144 48 146
rect 82 148 88 150
rect 82 146 84 148
rect 86 146 88 148
rect 82 144 88 146
rect 298 148 308 150
rect 298 146 302 148
rect 304 146 308 148
rect 298 144 308 146
rect 350 148 356 150
rect 350 146 352 148
rect 354 146 356 148
rect 350 144 356 146
rect 566 148 576 150
rect 566 146 570 148
rect 572 146 576 148
rect 566 144 576 146
rect 618 148 624 150
rect 618 146 620 148
rect 622 146 624 148
rect 618 144 624 146
rect 833 148 843 150
rect 833 146 837 148
rect 839 146 843 148
rect 833 144 843 146
rect 42 16 48 18
rect 42 14 44 16
rect 46 14 48 16
rect 42 12 48 14
rect 82 16 88 18
rect 82 14 84 16
rect 86 14 88 16
rect 82 12 88 14
rect 298 16 308 18
rect 298 14 302 16
rect 304 14 308 16
rect 298 12 308 14
rect 350 16 356 18
rect 350 14 352 16
rect 354 14 356 16
rect 350 12 356 14
rect 566 16 576 18
rect 566 14 570 16
rect 572 14 576 16
rect 566 12 576 14
rect 618 16 624 18
rect 618 14 620 16
rect 622 14 624 16
rect 618 12 624 14
rect 833 16 843 18
rect 833 14 837 16
rect 839 14 843 16
rect 833 12 843 14
<< ntie >>
rect 42 232 48 234
rect 42 230 44 232
rect 46 230 48 232
rect 42 228 48 230
rect 82 232 88 234
rect 82 230 84 232
rect 86 230 88 232
rect 82 228 88 230
rect 350 232 356 234
rect 350 230 352 232
rect 354 230 356 232
rect 350 228 356 230
rect 618 232 624 234
rect 618 230 620 232
rect 622 230 624 232
rect 618 228 624 230
rect 42 220 48 222
rect 42 218 44 220
rect 46 218 48 220
rect 42 216 48 218
rect 82 220 88 222
rect 82 218 84 220
rect 86 218 88 220
rect 82 216 88 218
rect 350 220 356 222
rect 350 218 352 220
rect 354 218 356 220
rect 350 216 356 218
rect 618 220 624 222
rect 618 218 620 220
rect 622 218 624 220
rect 618 216 624 218
rect 42 88 48 90
rect 42 86 44 88
rect 46 86 48 88
rect 42 84 48 86
rect 82 88 88 90
rect 82 86 84 88
rect 86 86 88 88
rect 82 84 88 86
rect 350 88 356 90
rect 350 86 352 88
rect 354 86 356 88
rect 350 84 356 86
rect 618 88 624 90
rect 618 86 620 88
rect 622 86 624 88
rect 618 84 624 86
rect 42 76 48 78
rect 42 74 44 76
rect 46 74 48 76
rect 42 72 48 74
rect 82 76 88 78
rect 82 74 84 76
rect 86 74 88 76
rect 82 72 88 74
rect 350 76 356 78
rect 350 74 352 76
rect 354 74 356 76
rect 350 72 356 74
rect 618 76 624 78
rect 618 74 620 76
rect 622 74 624 76
rect 618 72 624 74
<< nmos >>
rect 20 273 22 284
rect 27 273 29 284
rect 40 273 42 282
rect 60 273 62 284
rect 67 273 69 284
rect 80 273 82 282
rect 102 278 104 291
rect 112 278 114 288
rect 122 271 124 285
rect 132 271 134 285
rect 152 271 154 291
rect 159 271 161 291
rect 170 277 172 291
rect 191 278 193 291
rect 201 278 203 288
rect 211 271 213 285
rect 221 271 223 285
rect 241 271 243 291
rect 248 271 250 291
rect 259 277 261 291
rect 280 271 282 285
rect 290 276 292 284
rect 300 274 302 282
rect 328 273 330 284
rect 335 273 337 284
rect 348 273 350 282
rect 370 278 372 291
rect 380 278 382 288
rect 390 271 392 285
rect 400 271 402 285
rect 420 271 422 291
rect 427 271 429 291
rect 438 277 440 291
rect 459 278 461 291
rect 469 278 471 288
rect 479 271 481 285
rect 489 271 491 285
rect 509 271 511 291
rect 516 271 518 291
rect 527 277 529 291
rect 548 271 550 285
rect 558 276 560 284
rect 568 274 570 282
rect 596 273 598 284
rect 603 273 605 284
rect 616 273 618 282
rect 637 278 639 291
rect 647 278 649 288
rect 657 271 659 285
rect 667 271 669 285
rect 687 271 689 291
rect 694 271 696 291
rect 705 277 707 291
rect 726 278 728 291
rect 736 278 738 288
rect 746 271 748 285
rect 756 271 758 285
rect 776 271 778 291
rect 783 271 785 291
rect 794 277 796 291
rect 815 271 817 285
rect 825 276 827 284
rect 835 274 837 282
rect 20 166 22 177
rect 27 166 29 177
rect 40 168 42 177
rect 60 166 62 177
rect 67 166 69 177
rect 80 168 82 177
rect 102 159 104 172
rect 112 162 114 172
rect 122 165 124 179
rect 132 165 134 179
rect 152 159 154 179
rect 159 159 161 179
rect 170 159 172 173
rect 191 159 193 172
rect 201 162 203 172
rect 211 165 213 179
rect 221 165 223 179
rect 241 159 243 179
rect 248 159 250 179
rect 259 159 261 173
rect 280 165 282 179
rect 290 166 292 174
rect 300 168 302 176
rect 328 166 330 177
rect 335 166 337 177
rect 348 168 350 177
rect 370 159 372 172
rect 380 162 382 172
rect 390 165 392 179
rect 400 165 402 179
rect 420 159 422 179
rect 427 159 429 179
rect 438 159 440 173
rect 459 159 461 172
rect 469 162 471 172
rect 479 165 481 179
rect 489 165 491 179
rect 509 159 511 179
rect 516 159 518 179
rect 527 159 529 173
rect 548 165 550 179
rect 558 166 560 174
rect 568 168 570 176
rect 596 166 598 177
rect 603 166 605 177
rect 616 168 618 177
rect 637 159 639 172
rect 647 162 649 172
rect 657 165 659 179
rect 667 165 669 179
rect 687 159 689 179
rect 694 159 696 179
rect 705 159 707 173
rect 726 159 728 172
rect 736 162 738 172
rect 746 165 748 179
rect 756 165 758 179
rect 776 159 778 179
rect 783 159 785 179
rect 794 159 796 173
rect 815 165 817 179
rect 825 166 827 174
rect 835 168 837 176
rect 20 129 22 140
rect 27 129 29 140
rect 40 129 42 138
rect 60 129 62 140
rect 67 129 69 140
rect 80 129 82 138
rect 102 134 104 147
rect 112 134 114 144
rect 122 127 124 141
rect 132 127 134 141
rect 152 127 154 147
rect 159 127 161 147
rect 170 133 172 147
rect 191 134 193 147
rect 201 134 203 144
rect 211 127 213 141
rect 221 127 223 141
rect 241 127 243 147
rect 248 127 250 147
rect 259 133 261 147
rect 280 127 282 141
rect 290 132 292 140
rect 300 130 302 138
rect 328 129 330 140
rect 335 129 337 140
rect 348 129 350 138
rect 370 134 372 147
rect 380 134 382 144
rect 390 127 392 141
rect 400 127 402 141
rect 420 127 422 147
rect 427 127 429 147
rect 438 133 440 147
rect 459 134 461 147
rect 469 134 471 144
rect 479 127 481 141
rect 489 127 491 141
rect 509 127 511 147
rect 516 127 518 147
rect 527 133 529 147
rect 548 127 550 141
rect 558 132 560 140
rect 568 130 570 138
rect 596 129 598 140
rect 603 129 605 140
rect 616 129 618 138
rect 637 134 639 147
rect 647 134 649 144
rect 657 127 659 141
rect 667 127 669 141
rect 687 127 689 147
rect 694 127 696 147
rect 705 133 707 147
rect 726 134 728 147
rect 736 134 738 144
rect 746 127 748 141
rect 756 127 758 141
rect 776 127 778 147
rect 783 127 785 147
rect 794 133 796 147
rect 815 127 817 141
rect 825 132 827 140
rect 835 130 837 138
rect 20 22 22 33
rect 27 22 29 33
rect 40 24 42 33
rect 60 22 62 33
rect 67 22 69 33
rect 80 24 82 33
rect 102 15 104 28
rect 112 18 114 28
rect 122 21 124 35
rect 132 21 134 35
rect 152 15 154 35
rect 159 15 161 35
rect 170 15 172 29
rect 191 15 193 28
rect 201 18 203 28
rect 211 21 213 35
rect 221 21 223 35
rect 241 15 243 35
rect 248 15 250 35
rect 259 15 261 29
rect 280 21 282 35
rect 290 22 292 30
rect 300 24 302 32
rect 328 22 330 33
rect 335 22 337 33
rect 348 24 350 33
rect 370 15 372 28
rect 380 18 382 28
rect 390 21 392 35
rect 400 21 402 35
rect 420 15 422 35
rect 427 15 429 35
rect 438 15 440 29
rect 459 15 461 28
rect 469 18 471 28
rect 479 21 481 35
rect 489 21 491 35
rect 509 15 511 35
rect 516 15 518 35
rect 527 15 529 29
rect 548 21 550 35
rect 558 22 560 30
rect 568 24 570 32
rect 596 22 598 33
rect 603 22 605 33
rect 616 24 618 33
rect 637 15 639 28
rect 647 18 649 28
rect 657 21 659 35
rect 667 21 669 35
rect 687 15 689 35
rect 694 15 696 35
rect 705 15 707 29
rect 726 15 728 28
rect 736 18 738 28
rect 746 21 748 35
rect 756 21 758 35
rect 776 15 778 35
rect 783 15 785 35
rect 794 15 796 29
rect 815 21 817 35
rect 825 22 827 30
rect 835 24 837 32
<< pmos >>
rect 20 238 22 251
rect 30 238 32 251
rect 40 240 42 258
rect 60 238 62 251
rect 70 238 72 251
rect 80 240 82 258
rect 102 231 104 256
rect 115 243 117 256
rect 125 234 127 259
rect 132 234 134 259
rect 150 231 152 259
rect 160 231 162 259
rect 170 231 172 259
rect 191 231 193 256
rect 204 243 206 256
rect 214 234 216 259
rect 221 234 223 259
rect 239 231 241 259
rect 249 231 251 259
rect 259 231 261 259
rect 280 231 282 259
rect 293 231 295 259
rect 300 231 302 259
rect 328 238 330 251
rect 338 238 340 251
rect 348 240 350 258
rect 370 231 372 256
rect 383 243 385 256
rect 393 234 395 259
rect 400 234 402 259
rect 418 231 420 259
rect 428 231 430 259
rect 438 231 440 259
rect 459 231 461 256
rect 472 243 474 256
rect 482 234 484 259
rect 489 234 491 259
rect 507 231 509 259
rect 517 231 519 259
rect 527 231 529 259
rect 548 231 550 259
rect 561 231 563 259
rect 568 231 570 259
rect 596 238 598 251
rect 606 238 608 251
rect 616 240 618 258
rect 637 231 639 256
rect 650 243 652 256
rect 660 234 662 259
rect 667 234 669 259
rect 685 231 687 259
rect 695 231 697 259
rect 705 231 707 259
rect 726 231 728 256
rect 739 243 741 256
rect 749 234 751 259
rect 756 234 758 259
rect 774 231 776 259
rect 784 231 786 259
rect 794 231 796 259
rect 815 231 817 259
rect 828 231 830 259
rect 835 231 837 259
rect 20 199 22 212
rect 30 199 32 212
rect 40 192 42 210
rect 60 199 62 212
rect 70 199 72 212
rect 80 192 82 210
rect 102 194 104 219
rect 115 194 117 207
rect 125 191 127 216
rect 132 191 134 216
rect 150 191 152 219
rect 160 191 162 219
rect 170 191 172 219
rect 191 194 193 219
rect 204 194 206 207
rect 214 191 216 216
rect 221 191 223 216
rect 239 191 241 219
rect 249 191 251 219
rect 259 191 261 219
rect 280 191 282 219
rect 293 191 295 219
rect 300 191 302 219
rect 328 199 330 212
rect 338 199 340 212
rect 348 192 350 210
rect 370 194 372 219
rect 383 194 385 207
rect 393 191 395 216
rect 400 191 402 216
rect 418 191 420 219
rect 428 191 430 219
rect 438 191 440 219
rect 459 194 461 219
rect 472 194 474 207
rect 482 191 484 216
rect 489 191 491 216
rect 507 191 509 219
rect 517 191 519 219
rect 527 191 529 219
rect 548 191 550 219
rect 561 191 563 219
rect 568 191 570 219
rect 596 199 598 212
rect 606 199 608 212
rect 616 192 618 210
rect 637 194 639 219
rect 650 194 652 207
rect 660 191 662 216
rect 667 191 669 216
rect 685 191 687 219
rect 695 191 697 219
rect 705 191 707 219
rect 726 194 728 219
rect 739 194 741 207
rect 749 191 751 216
rect 756 191 758 216
rect 774 191 776 219
rect 784 191 786 219
rect 794 191 796 219
rect 815 191 817 219
rect 828 191 830 219
rect 835 191 837 219
rect 20 94 22 107
rect 30 94 32 107
rect 40 96 42 114
rect 60 94 62 107
rect 70 94 72 107
rect 80 96 82 114
rect 102 87 104 112
rect 115 99 117 112
rect 125 90 127 115
rect 132 90 134 115
rect 150 87 152 115
rect 160 87 162 115
rect 170 87 172 115
rect 191 87 193 112
rect 204 99 206 112
rect 214 90 216 115
rect 221 90 223 115
rect 239 87 241 115
rect 249 87 251 115
rect 259 87 261 115
rect 280 87 282 115
rect 293 87 295 115
rect 300 87 302 115
rect 328 94 330 107
rect 338 94 340 107
rect 348 96 350 114
rect 370 87 372 112
rect 383 99 385 112
rect 393 90 395 115
rect 400 90 402 115
rect 418 87 420 115
rect 428 87 430 115
rect 438 87 440 115
rect 459 87 461 112
rect 472 99 474 112
rect 482 90 484 115
rect 489 90 491 115
rect 507 87 509 115
rect 517 87 519 115
rect 527 87 529 115
rect 548 87 550 115
rect 561 87 563 115
rect 568 87 570 115
rect 596 94 598 107
rect 606 94 608 107
rect 616 96 618 114
rect 637 87 639 112
rect 650 99 652 112
rect 660 90 662 115
rect 667 90 669 115
rect 685 87 687 115
rect 695 87 697 115
rect 705 87 707 115
rect 726 87 728 112
rect 739 99 741 112
rect 749 90 751 115
rect 756 90 758 115
rect 774 87 776 115
rect 784 87 786 115
rect 794 87 796 115
rect 815 87 817 115
rect 828 87 830 115
rect 835 87 837 115
rect 20 55 22 68
rect 30 55 32 68
rect 40 48 42 66
rect 60 55 62 68
rect 70 55 72 68
rect 80 48 82 66
rect 102 50 104 75
rect 115 50 117 63
rect 125 47 127 72
rect 132 47 134 72
rect 150 47 152 75
rect 160 47 162 75
rect 170 47 172 75
rect 191 50 193 75
rect 204 50 206 63
rect 214 47 216 72
rect 221 47 223 72
rect 239 47 241 75
rect 249 47 251 75
rect 259 47 261 75
rect 280 47 282 75
rect 293 47 295 75
rect 300 47 302 75
rect 328 55 330 68
rect 338 55 340 68
rect 348 48 350 66
rect 370 50 372 75
rect 383 50 385 63
rect 393 47 395 72
rect 400 47 402 72
rect 418 47 420 75
rect 428 47 430 75
rect 438 47 440 75
rect 459 50 461 75
rect 472 50 474 63
rect 482 47 484 72
rect 489 47 491 72
rect 507 47 509 75
rect 517 47 519 75
rect 527 47 529 75
rect 548 47 550 75
rect 561 47 563 75
rect 568 47 570 75
rect 596 55 598 68
rect 606 55 608 68
rect 616 48 618 66
rect 637 50 639 75
rect 650 50 652 63
rect 660 47 662 72
rect 667 47 669 72
rect 685 47 687 75
rect 695 47 697 75
rect 705 47 707 75
rect 726 50 728 75
rect 739 50 741 63
rect 749 47 751 72
rect 756 47 758 72
rect 774 47 776 75
rect 784 47 786 75
rect 794 47 796 75
rect 815 47 817 75
rect 828 47 830 75
rect 835 47 837 75
<< polyct0 >>
rect 38 264 40 266
rect 78 264 80 266
rect 104 271 106 273
rect 110 261 112 263
rect 193 271 195 273
rect 160 264 162 266
rect 170 264 172 266
rect 199 261 201 263
rect 249 264 251 266
rect 259 264 261 266
rect 282 264 284 266
rect 346 264 348 266
rect 372 271 374 273
rect 378 261 380 263
rect 461 271 463 273
rect 428 264 430 266
rect 438 264 440 266
rect 467 261 469 263
rect 517 264 519 266
rect 527 264 529 266
rect 550 264 552 266
rect 614 264 616 266
rect 639 271 641 273
rect 645 261 647 263
rect 728 271 730 273
rect 695 264 697 266
rect 705 264 707 266
rect 734 261 736 263
rect 784 264 786 266
rect 794 264 796 266
rect 817 264 819 266
rect 38 184 40 186
rect 78 184 80 186
rect 110 187 112 189
rect 104 177 106 179
rect 160 184 162 186
rect 170 184 172 186
rect 199 187 201 189
rect 193 177 195 179
rect 249 184 251 186
rect 259 184 261 186
rect 282 184 284 186
rect 346 184 348 186
rect 378 187 380 189
rect 372 177 374 179
rect 428 184 430 186
rect 438 184 440 186
rect 467 187 469 189
rect 461 177 463 179
rect 517 184 519 186
rect 527 184 529 186
rect 550 184 552 186
rect 614 184 616 186
rect 645 187 647 189
rect 639 177 641 179
rect 695 184 697 186
rect 705 184 707 186
rect 734 187 736 189
rect 728 177 730 179
rect 784 184 786 186
rect 794 184 796 186
rect 817 184 819 186
rect 38 120 40 122
rect 78 120 80 122
rect 104 127 106 129
rect 110 117 112 119
rect 193 127 195 129
rect 160 120 162 122
rect 170 120 172 122
rect 199 117 201 119
rect 249 120 251 122
rect 259 120 261 122
rect 282 120 284 122
rect 346 120 348 122
rect 372 127 374 129
rect 378 117 380 119
rect 461 127 463 129
rect 428 120 430 122
rect 438 120 440 122
rect 467 117 469 119
rect 517 120 519 122
rect 527 120 529 122
rect 550 120 552 122
rect 614 120 616 122
rect 639 127 641 129
rect 645 117 647 119
rect 728 127 730 129
rect 695 120 697 122
rect 705 120 707 122
rect 734 117 736 119
rect 784 120 786 122
rect 794 120 796 122
rect 817 120 819 122
rect 38 40 40 42
rect 78 40 80 42
rect 110 43 112 45
rect 104 33 106 35
rect 160 40 162 42
rect 170 40 172 42
rect 199 43 201 45
rect 193 33 195 35
rect 249 40 251 42
rect 259 40 261 42
rect 282 40 284 42
rect 346 40 348 42
rect 378 43 380 45
rect 372 33 374 35
rect 428 40 430 42
rect 438 40 440 42
rect 467 43 469 45
rect 461 33 463 35
rect 517 40 519 42
rect 527 40 529 42
rect 550 40 552 42
rect 614 40 616 42
rect 645 43 647 45
rect 639 33 641 35
rect 695 40 697 42
rect 705 40 707 42
rect 734 43 736 45
rect 728 33 730 35
rect 784 40 786 42
rect 794 40 796 42
rect 817 40 819 42
<< polyct1 >>
rect 28 264 30 266
rect 18 256 20 258
rect 68 264 70 266
rect 58 256 60 258
rect 124 264 126 266
rect 143 264 145 266
rect 150 264 152 266
rect 213 264 215 266
rect 232 264 234 266
rect 239 264 241 266
rect 292 264 294 266
rect 305 264 307 266
rect 336 264 338 266
rect 326 256 328 258
rect 392 264 394 266
rect 411 264 413 266
rect 418 264 420 266
rect 481 264 483 266
rect 500 264 502 266
rect 507 264 509 266
rect 560 264 562 266
rect 573 264 575 266
rect 604 264 606 266
rect 594 256 596 258
rect 659 264 661 266
rect 678 264 680 266
rect 685 264 687 266
rect 748 264 750 266
rect 767 264 769 266
rect 774 264 776 266
rect 827 264 829 266
rect 840 264 842 266
rect 18 192 20 194
rect 58 192 60 194
rect 28 184 30 186
rect 68 184 70 186
rect 124 184 126 186
rect 143 184 145 186
rect 150 184 152 186
rect 326 192 328 194
rect 213 184 215 186
rect 232 184 234 186
rect 239 184 241 186
rect 292 184 294 186
rect 305 184 307 186
rect 336 184 338 186
rect 392 184 394 186
rect 411 184 413 186
rect 418 184 420 186
rect 594 192 596 194
rect 481 184 483 186
rect 500 184 502 186
rect 507 184 509 186
rect 560 184 562 186
rect 573 184 575 186
rect 604 184 606 186
rect 659 184 661 186
rect 678 184 680 186
rect 685 184 687 186
rect 748 184 750 186
rect 767 184 769 186
rect 774 184 776 186
rect 827 184 829 186
rect 840 184 842 186
rect 28 120 30 122
rect 18 112 20 114
rect 68 120 70 122
rect 58 112 60 114
rect 124 120 126 122
rect 143 120 145 122
rect 150 120 152 122
rect 213 120 215 122
rect 232 120 234 122
rect 239 120 241 122
rect 292 120 294 122
rect 305 120 307 122
rect 336 120 338 122
rect 326 112 328 114
rect 392 120 394 122
rect 411 120 413 122
rect 418 120 420 122
rect 481 120 483 122
rect 500 120 502 122
rect 507 120 509 122
rect 560 120 562 122
rect 573 120 575 122
rect 604 120 606 122
rect 594 112 596 114
rect 659 120 661 122
rect 678 120 680 122
rect 685 120 687 122
rect 748 120 750 122
rect 767 120 769 122
rect 774 120 776 122
rect 827 120 829 122
rect 840 120 842 122
rect 18 48 20 50
rect 58 48 60 50
rect 28 40 30 42
rect 68 40 70 42
rect 124 40 126 42
rect 143 40 145 42
rect 150 40 152 42
rect 326 48 328 50
rect 213 40 215 42
rect 232 40 234 42
rect 239 40 241 42
rect 292 40 294 42
rect 305 40 307 42
rect 336 40 338 42
rect 392 40 394 42
rect 411 40 413 42
rect 418 40 420 42
rect 594 48 596 50
rect 481 40 483 42
rect 500 40 502 42
rect 507 40 509 42
rect 560 40 562 42
rect 573 40 575 42
rect 604 40 606 42
rect 659 40 661 42
rect 678 40 680 42
rect 685 40 687 42
rect 748 40 750 42
rect 767 40 769 42
rect 774 40 776 42
rect 827 40 829 42
rect 840 40 842 42
<< ndifct0 >>
rect 15 280 17 282
rect 55 280 57 282
rect 107 284 109 286
rect 117 281 119 283
rect 127 273 129 275
rect 137 280 139 282
rect 147 280 149 282
rect 137 273 139 275
rect 164 287 166 289
rect 196 284 198 286
rect 206 281 208 283
rect 216 273 218 275
rect 226 280 228 282
rect 236 280 238 282
rect 226 273 228 275
rect 253 287 255 289
rect 285 280 287 282
rect 295 278 297 280
rect 305 278 307 280
rect 323 280 325 282
rect 375 284 377 286
rect 385 281 387 283
rect 395 273 397 275
rect 405 280 407 282
rect 415 280 417 282
rect 405 273 407 275
rect 432 287 434 289
rect 464 284 466 286
rect 474 281 476 283
rect 484 273 486 275
rect 494 280 496 282
rect 504 280 506 282
rect 494 273 496 275
rect 521 287 523 289
rect 553 280 555 282
rect 563 278 565 280
rect 573 278 575 280
rect 591 280 593 282
rect 642 284 644 286
rect 652 281 654 283
rect 662 273 664 275
rect 672 280 674 282
rect 682 280 684 282
rect 672 273 674 275
rect 699 287 701 289
rect 731 284 733 286
rect 741 281 743 283
rect 751 273 753 275
rect 761 280 763 282
rect 771 280 773 282
rect 761 273 763 275
rect 788 287 790 289
rect 820 280 822 282
rect 830 278 832 280
rect 840 278 842 280
rect 15 168 17 170
rect 55 168 57 170
rect 107 164 109 166
rect 117 167 119 169
rect 127 175 129 177
rect 137 175 139 177
rect 137 168 139 170
rect 147 168 149 170
rect 164 161 166 163
rect 196 164 198 166
rect 206 167 208 169
rect 216 175 218 177
rect 226 175 228 177
rect 226 168 228 170
rect 236 168 238 170
rect 253 161 255 163
rect 285 168 287 170
rect 295 170 297 172
rect 305 170 307 172
rect 323 168 325 170
rect 375 164 377 166
rect 385 167 387 169
rect 395 175 397 177
rect 405 175 407 177
rect 405 168 407 170
rect 415 168 417 170
rect 432 161 434 163
rect 464 164 466 166
rect 474 167 476 169
rect 484 175 486 177
rect 494 175 496 177
rect 494 168 496 170
rect 504 168 506 170
rect 521 161 523 163
rect 553 168 555 170
rect 563 170 565 172
rect 573 170 575 172
rect 591 168 593 170
rect 642 164 644 166
rect 652 167 654 169
rect 662 175 664 177
rect 672 175 674 177
rect 672 168 674 170
rect 682 168 684 170
rect 699 161 701 163
rect 731 164 733 166
rect 741 167 743 169
rect 751 175 753 177
rect 761 175 763 177
rect 761 168 763 170
rect 771 168 773 170
rect 788 161 790 163
rect 820 168 822 170
rect 830 170 832 172
rect 840 170 842 172
rect 15 136 17 138
rect 55 136 57 138
rect 107 140 109 142
rect 117 137 119 139
rect 127 129 129 131
rect 137 136 139 138
rect 147 136 149 138
rect 137 129 139 131
rect 164 143 166 145
rect 196 140 198 142
rect 206 137 208 139
rect 216 129 218 131
rect 226 136 228 138
rect 236 136 238 138
rect 226 129 228 131
rect 253 143 255 145
rect 285 136 287 138
rect 295 134 297 136
rect 305 134 307 136
rect 323 136 325 138
rect 375 140 377 142
rect 385 137 387 139
rect 395 129 397 131
rect 405 136 407 138
rect 415 136 417 138
rect 405 129 407 131
rect 432 143 434 145
rect 464 140 466 142
rect 474 137 476 139
rect 484 129 486 131
rect 494 136 496 138
rect 504 136 506 138
rect 494 129 496 131
rect 521 143 523 145
rect 553 136 555 138
rect 563 134 565 136
rect 573 134 575 136
rect 591 136 593 138
rect 642 140 644 142
rect 652 137 654 139
rect 662 129 664 131
rect 672 136 674 138
rect 682 136 684 138
rect 672 129 674 131
rect 699 143 701 145
rect 731 140 733 142
rect 741 137 743 139
rect 751 129 753 131
rect 761 136 763 138
rect 771 136 773 138
rect 761 129 763 131
rect 788 143 790 145
rect 820 136 822 138
rect 830 134 832 136
rect 840 134 842 136
rect 15 24 17 26
rect 55 24 57 26
rect 107 20 109 22
rect 117 23 119 25
rect 127 31 129 33
rect 137 31 139 33
rect 137 24 139 26
rect 147 24 149 26
rect 164 17 166 19
rect 196 20 198 22
rect 206 23 208 25
rect 216 31 218 33
rect 226 31 228 33
rect 226 24 228 26
rect 236 24 238 26
rect 253 17 255 19
rect 285 24 287 26
rect 295 26 297 28
rect 305 26 307 28
rect 323 24 325 26
rect 375 20 377 22
rect 385 23 387 25
rect 395 31 397 33
rect 405 31 407 33
rect 405 24 407 26
rect 415 24 417 26
rect 432 17 434 19
rect 464 20 466 22
rect 474 23 476 25
rect 484 31 486 33
rect 494 31 496 33
rect 494 24 496 26
rect 504 24 506 26
rect 521 17 523 19
rect 553 24 555 26
rect 563 26 565 28
rect 573 26 575 28
rect 591 24 593 26
rect 642 20 644 22
rect 652 23 654 25
rect 662 31 664 33
rect 672 31 674 33
rect 672 24 674 26
rect 682 24 684 26
rect 699 17 701 19
rect 731 20 733 22
rect 741 23 743 25
rect 751 31 753 33
rect 761 31 763 33
rect 761 24 763 26
rect 771 24 773 26
rect 788 17 790 19
rect 820 24 822 26
rect 830 26 832 28
rect 840 26 842 28
<< ndifct1 >>
rect 34 290 36 292
rect 74 290 76 292
rect 45 278 47 280
rect 85 278 87 280
rect 97 280 99 282
rect 175 280 177 282
rect 186 280 188 282
rect 264 280 266 282
rect 275 280 277 282
rect 275 273 277 275
rect 342 290 344 292
rect 353 278 355 280
rect 365 280 367 282
rect 443 280 445 282
rect 454 280 456 282
rect 532 280 534 282
rect 543 280 545 282
rect 543 273 545 275
rect 610 290 612 292
rect 621 278 623 280
rect 632 280 634 282
rect 710 280 712 282
rect 721 280 723 282
rect 799 280 801 282
rect 810 280 812 282
rect 810 273 812 275
rect 45 170 47 172
rect 85 170 87 172
rect 97 168 99 170
rect 34 158 36 160
rect 74 158 76 160
rect 175 168 177 170
rect 186 168 188 170
rect 275 175 277 177
rect 264 168 266 170
rect 275 168 277 170
rect 353 170 355 172
rect 365 168 367 170
rect 342 158 344 160
rect 443 168 445 170
rect 454 168 456 170
rect 543 175 545 177
rect 532 168 534 170
rect 543 168 545 170
rect 621 170 623 172
rect 632 168 634 170
rect 610 158 612 160
rect 710 168 712 170
rect 721 168 723 170
rect 810 175 812 177
rect 799 168 801 170
rect 810 168 812 170
rect 34 146 36 148
rect 74 146 76 148
rect 45 134 47 136
rect 85 134 87 136
rect 97 136 99 138
rect 175 136 177 138
rect 186 136 188 138
rect 264 136 266 138
rect 275 136 277 138
rect 275 129 277 131
rect 342 146 344 148
rect 353 134 355 136
rect 365 136 367 138
rect 443 136 445 138
rect 454 136 456 138
rect 532 136 534 138
rect 543 136 545 138
rect 543 129 545 131
rect 610 146 612 148
rect 621 134 623 136
rect 632 136 634 138
rect 710 136 712 138
rect 721 136 723 138
rect 799 136 801 138
rect 810 136 812 138
rect 810 129 812 131
rect 45 26 47 28
rect 85 26 87 28
rect 97 24 99 26
rect 34 14 36 16
rect 74 14 76 16
rect 175 24 177 26
rect 186 24 188 26
rect 275 31 277 33
rect 264 24 266 26
rect 275 24 277 26
rect 353 26 355 28
rect 365 24 367 26
rect 342 14 344 16
rect 443 24 445 26
rect 454 24 456 26
rect 543 31 545 33
rect 532 24 534 26
rect 543 24 545 26
rect 621 26 623 28
rect 632 24 634 26
rect 610 14 612 16
rect 710 24 712 26
rect 721 24 723 26
rect 810 31 812 33
rect 799 24 801 26
rect 810 24 812 26
<< ntiect1 >>
rect 44 230 46 232
rect 84 230 86 232
rect 352 230 354 232
rect 620 230 622 232
rect 44 218 46 220
rect 84 218 86 220
rect 352 218 354 220
rect 620 218 622 220
rect 44 86 46 88
rect 84 86 86 88
rect 352 86 354 88
rect 620 86 622 88
rect 44 74 46 76
rect 84 74 86 76
rect 352 74 354 76
rect 620 74 622 76
<< ptiect1 >>
rect 44 290 46 292
rect 84 290 86 292
rect 302 290 304 292
rect 352 290 354 292
rect 570 290 572 292
rect 620 290 622 292
rect 837 290 839 292
rect 44 158 46 160
rect 84 158 86 160
rect 302 158 304 160
rect 352 158 354 160
rect 570 158 572 160
rect 620 158 622 160
rect 837 158 839 160
rect 44 146 46 148
rect 84 146 86 148
rect 302 146 304 148
rect 352 146 354 148
rect 570 146 572 148
rect 620 146 622 148
rect 837 146 839 148
rect 44 14 46 16
rect 84 14 86 16
rect 302 14 304 16
rect 352 14 354 16
rect 570 14 572 16
rect 620 14 622 16
rect 837 14 839 16
<< pdifct0 >>
rect 15 240 17 242
rect 25 247 27 249
rect 25 240 27 242
rect 35 242 37 244
rect 55 240 57 242
rect 65 247 67 249
rect 65 240 67 242
rect 75 242 77 244
rect 120 252 122 254
rect 108 233 110 235
rect 143 240 145 242
rect 143 233 145 235
rect 155 248 157 250
rect 155 241 157 243
rect 165 240 167 242
rect 165 233 167 235
rect 209 252 211 254
rect 197 233 199 235
rect 232 240 234 242
rect 232 233 234 235
rect 244 248 246 250
rect 244 241 246 243
rect 254 240 256 242
rect 254 233 256 235
rect 305 239 307 241
rect 323 240 325 242
rect 333 247 335 249
rect 333 240 335 242
rect 343 242 345 244
rect 388 252 390 254
rect 376 233 378 235
rect 411 240 413 242
rect 411 233 413 235
rect 423 248 425 250
rect 423 241 425 243
rect 433 240 435 242
rect 433 233 435 235
rect 477 252 479 254
rect 465 233 467 235
rect 500 240 502 242
rect 500 233 502 235
rect 512 248 514 250
rect 512 241 514 243
rect 522 240 524 242
rect 522 233 524 235
rect 573 239 575 241
rect 591 240 593 242
rect 601 247 603 249
rect 601 240 603 242
rect 611 242 613 244
rect 655 252 657 254
rect 643 233 645 235
rect 678 240 680 242
rect 678 233 680 235
rect 690 248 692 250
rect 690 241 692 243
rect 700 240 702 242
rect 700 233 702 235
rect 744 252 746 254
rect 732 233 734 235
rect 767 240 769 242
rect 767 233 769 235
rect 779 248 781 250
rect 779 241 781 243
rect 789 240 791 242
rect 789 233 791 235
rect 840 239 842 241
rect 15 208 17 210
rect 25 208 27 210
rect 25 201 27 203
rect 35 206 37 208
rect 55 208 57 210
rect 65 208 67 210
rect 65 201 67 203
rect 75 206 77 208
rect 108 215 110 217
rect 120 196 122 198
rect 143 215 145 217
rect 143 208 145 210
rect 155 207 157 209
rect 155 200 157 202
rect 165 215 167 217
rect 165 208 167 210
rect 197 215 199 217
rect 209 196 211 198
rect 232 215 234 217
rect 232 208 234 210
rect 244 207 246 209
rect 244 200 246 202
rect 254 215 256 217
rect 254 208 256 210
rect 305 209 307 211
rect 323 208 325 210
rect 333 208 335 210
rect 333 201 335 203
rect 343 206 345 208
rect 376 215 378 217
rect 388 196 390 198
rect 411 215 413 217
rect 411 208 413 210
rect 423 207 425 209
rect 423 200 425 202
rect 433 215 435 217
rect 433 208 435 210
rect 465 215 467 217
rect 477 196 479 198
rect 500 215 502 217
rect 500 208 502 210
rect 512 207 514 209
rect 512 200 514 202
rect 522 215 524 217
rect 522 208 524 210
rect 573 209 575 211
rect 591 208 593 210
rect 601 208 603 210
rect 601 201 603 203
rect 611 206 613 208
rect 643 215 645 217
rect 655 196 657 198
rect 678 215 680 217
rect 678 208 680 210
rect 690 207 692 209
rect 690 200 692 202
rect 700 215 702 217
rect 700 208 702 210
rect 732 215 734 217
rect 744 196 746 198
rect 767 215 769 217
rect 767 208 769 210
rect 779 207 781 209
rect 779 200 781 202
rect 789 215 791 217
rect 789 208 791 210
rect 840 209 842 211
rect 15 96 17 98
rect 25 103 27 105
rect 25 96 27 98
rect 35 98 37 100
rect 55 96 57 98
rect 65 103 67 105
rect 65 96 67 98
rect 75 98 77 100
rect 120 108 122 110
rect 108 89 110 91
rect 143 96 145 98
rect 143 89 145 91
rect 155 104 157 106
rect 155 97 157 99
rect 165 96 167 98
rect 165 89 167 91
rect 209 108 211 110
rect 197 89 199 91
rect 232 96 234 98
rect 232 89 234 91
rect 244 104 246 106
rect 244 97 246 99
rect 254 96 256 98
rect 254 89 256 91
rect 305 95 307 97
rect 323 96 325 98
rect 333 103 335 105
rect 333 96 335 98
rect 343 98 345 100
rect 388 108 390 110
rect 376 89 378 91
rect 411 96 413 98
rect 411 89 413 91
rect 423 104 425 106
rect 423 97 425 99
rect 433 96 435 98
rect 433 89 435 91
rect 477 108 479 110
rect 465 89 467 91
rect 500 96 502 98
rect 500 89 502 91
rect 512 104 514 106
rect 512 97 514 99
rect 522 96 524 98
rect 522 89 524 91
rect 573 95 575 97
rect 591 96 593 98
rect 601 103 603 105
rect 601 96 603 98
rect 611 98 613 100
rect 655 108 657 110
rect 643 89 645 91
rect 678 96 680 98
rect 678 89 680 91
rect 690 104 692 106
rect 690 97 692 99
rect 700 96 702 98
rect 700 89 702 91
rect 744 108 746 110
rect 732 89 734 91
rect 767 96 769 98
rect 767 89 769 91
rect 779 104 781 106
rect 779 97 781 99
rect 789 96 791 98
rect 789 89 791 91
rect 840 95 842 97
rect 15 64 17 66
rect 25 64 27 66
rect 25 57 27 59
rect 35 62 37 64
rect 55 64 57 66
rect 65 64 67 66
rect 65 57 67 59
rect 75 62 77 64
rect 108 71 110 73
rect 120 52 122 54
rect 143 71 145 73
rect 143 64 145 66
rect 155 63 157 65
rect 155 56 157 58
rect 165 71 167 73
rect 165 64 167 66
rect 197 71 199 73
rect 209 52 211 54
rect 232 71 234 73
rect 232 64 234 66
rect 244 63 246 65
rect 244 56 246 58
rect 254 71 256 73
rect 254 64 256 66
rect 305 65 307 67
rect 323 64 325 66
rect 333 64 335 66
rect 333 57 335 59
rect 343 62 345 64
rect 376 71 378 73
rect 388 52 390 54
rect 411 71 413 73
rect 411 64 413 66
rect 423 63 425 65
rect 423 56 425 58
rect 433 71 435 73
rect 433 64 435 66
rect 465 71 467 73
rect 477 52 479 54
rect 500 71 502 73
rect 500 64 502 66
rect 512 63 514 65
rect 512 56 514 58
rect 522 71 524 73
rect 522 64 524 66
rect 573 65 575 67
rect 591 64 593 66
rect 601 64 603 66
rect 601 57 603 59
rect 611 62 613 64
rect 643 71 645 73
rect 655 52 657 54
rect 678 71 680 73
rect 678 64 680 66
rect 690 63 692 65
rect 690 56 692 58
rect 700 71 702 73
rect 700 64 702 66
rect 732 71 734 73
rect 744 52 746 54
rect 767 71 769 73
rect 767 64 769 66
rect 779 63 781 65
rect 779 56 781 58
rect 789 71 791 73
rect 789 64 791 66
rect 840 65 842 67
<< pdifct1 >>
rect 45 254 47 256
rect 45 247 47 249
rect 85 254 87 256
rect 85 247 87 249
rect 97 252 99 254
rect 97 245 99 247
rect 175 255 177 257
rect 175 248 177 250
rect 186 252 188 254
rect 186 245 188 247
rect 264 255 266 257
rect 264 248 266 250
rect 275 246 277 248
rect 275 239 277 241
rect 286 230 288 232
rect 353 254 355 256
rect 353 247 355 249
rect 365 252 367 254
rect 365 245 367 247
rect 443 255 445 257
rect 443 248 445 250
rect 454 252 456 254
rect 454 245 456 247
rect 532 255 534 257
rect 532 248 534 250
rect 543 246 545 248
rect 543 239 545 241
rect 554 230 556 232
rect 621 254 623 256
rect 621 247 623 249
rect 632 252 634 254
rect 632 245 634 247
rect 710 255 712 257
rect 710 248 712 250
rect 721 252 723 254
rect 721 245 723 247
rect 799 255 801 257
rect 799 248 801 250
rect 810 246 812 248
rect 810 239 812 241
rect 821 230 823 232
rect 45 201 47 203
rect 45 194 47 196
rect 85 201 87 203
rect 85 194 87 196
rect 97 203 99 205
rect 97 196 99 198
rect 175 200 177 202
rect 175 193 177 195
rect 186 203 188 205
rect 186 196 188 198
rect 275 209 277 211
rect 264 200 266 202
rect 275 202 277 204
rect 264 193 266 195
rect 286 218 288 220
rect 353 201 355 203
rect 353 194 355 196
rect 365 203 367 205
rect 365 196 367 198
rect 443 200 445 202
rect 443 193 445 195
rect 454 203 456 205
rect 454 196 456 198
rect 543 209 545 211
rect 532 200 534 202
rect 543 202 545 204
rect 532 193 534 195
rect 554 218 556 220
rect 621 201 623 203
rect 621 194 623 196
rect 632 203 634 205
rect 632 196 634 198
rect 710 200 712 202
rect 710 193 712 195
rect 721 203 723 205
rect 721 196 723 198
rect 810 209 812 211
rect 799 200 801 202
rect 810 202 812 204
rect 799 193 801 195
rect 821 218 823 220
rect 45 110 47 112
rect 45 103 47 105
rect 85 110 87 112
rect 85 103 87 105
rect 97 108 99 110
rect 97 101 99 103
rect 175 111 177 113
rect 175 104 177 106
rect 186 108 188 110
rect 186 101 188 103
rect 264 111 266 113
rect 264 104 266 106
rect 275 102 277 104
rect 275 95 277 97
rect 286 86 288 88
rect 353 110 355 112
rect 353 103 355 105
rect 365 108 367 110
rect 365 101 367 103
rect 443 111 445 113
rect 443 104 445 106
rect 454 108 456 110
rect 454 101 456 103
rect 532 111 534 113
rect 532 104 534 106
rect 543 102 545 104
rect 543 95 545 97
rect 554 86 556 88
rect 621 110 623 112
rect 621 103 623 105
rect 632 108 634 110
rect 632 101 634 103
rect 710 111 712 113
rect 710 104 712 106
rect 721 108 723 110
rect 721 101 723 103
rect 799 111 801 113
rect 799 104 801 106
rect 810 102 812 104
rect 810 95 812 97
rect 821 86 823 88
rect 45 57 47 59
rect 45 50 47 52
rect 85 57 87 59
rect 85 50 87 52
rect 97 59 99 61
rect 97 52 99 54
rect 175 56 177 58
rect 175 49 177 51
rect 186 59 188 61
rect 186 52 188 54
rect 275 65 277 67
rect 264 56 266 58
rect 275 58 277 60
rect 264 49 266 51
rect 286 74 288 76
rect 353 57 355 59
rect 353 50 355 52
rect 365 59 367 61
rect 365 52 367 54
rect 443 56 445 58
rect 443 49 445 51
rect 454 59 456 61
rect 454 52 456 54
rect 543 65 545 67
rect 532 56 534 58
rect 543 58 545 60
rect 532 49 534 51
rect 554 74 556 76
rect 621 57 623 59
rect 621 50 623 52
rect 632 59 634 61
rect 632 52 634 54
rect 710 56 712 58
rect 710 49 712 51
rect 721 59 723 61
rect 721 52 723 54
rect 810 65 812 67
rect 799 56 801 58
rect 810 58 812 60
rect 799 49 801 51
rect 821 74 823 76
<< alu0 >>
rect 106 286 110 289
rect 162 287 164 289
rect 166 287 168 289
rect 162 286 168 287
rect 195 286 199 289
rect 251 287 253 289
rect 255 287 257 289
rect 251 286 257 287
rect 106 284 107 286
rect 109 284 110 286
rect 195 284 196 286
rect 198 284 199 286
rect 13 282 33 283
rect 13 280 15 282
rect 17 280 33 282
rect 13 279 33 280
rect 29 275 33 279
rect 53 282 73 283
rect 53 280 55 282
rect 57 280 73 282
rect 53 279 73 280
rect 44 276 45 278
rect 29 271 41 275
rect 37 266 41 271
rect 37 264 38 266
rect 40 264 41 266
rect 37 252 41 264
rect 69 275 73 279
rect 84 276 85 278
rect 69 271 81 275
rect 77 266 81 271
rect 77 264 78 266
rect 80 264 81 266
rect 24 249 41 252
rect 24 247 25 249
rect 27 248 41 249
rect 27 247 28 248
rect 13 242 19 243
rect 13 240 15 242
rect 17 240 19 242
rect 13 233 19 240
rect 24 242 28 247
rect 77 252 81 264
rect 64 249 81 252
rect 64 247 65 249
rect 67 248 81 249
rect 67 247 68 248
rect 24 240 25 242
rect 27 240 28 242
rect 24 238 28 240
rect 33 244 39 245
rect 33 242 35 244
rect 37 242 39 244
rect 33 233 39 242
rect 53 242 59 243
rect 53 240 55 242
rect 57 240 59 242
rect 53 233 59 240
rect 64 242 68 247
rect 106 282 110 284
rect 115 283 140 284
rect 115 281 117 283
rect 119 282 140 283
rect 119 281 137 282
rect 115 280 137 281
rect 139 280 140 282
rect 116 275 131 276
rect 116 274 127 275
rect 102 273 127 274
rect 129 273 131 275
rect 102 271 104 273
rect 106 272 131 273
rect 136 275 140 280
rect 145 282 155 283
rect 145 280 147 282
rect 149 280 155 282
rect 145 279 155 280
rect 136 273 137 275
rect 139 273 140 275
rect 106 271 120 272
rect 136 271 140 273
rect 102 270 120 271
rect 109 263 113 265
rect 109 261 110 263
rect 112 261 113 263
rect 109 251 113 261
rect 116 259 120 270
rect 151 275 155 279
rect 151 271 171 275
rect 167 268 171 271
rect 159 266 163 268
rect 159 264 160 266
rect 162 264 163 266
rect 159 259 163 264
rect 167 266 173 268
rect 167 264 170 266
rect 172 264 173 266
rect 167 262 173 264
rect 116 255 123 259
rect 119 254 123 255
rect 119 252 120 254
rect 122 252 123 254
rect 109 247 115 251
rect 119 250 123 252
rect 167 251 171 262
rect 131 250 171 251
rect 131 248 155 250
rect 157 248 171 250
rect 131 247 171 248
rect 64 240 65 242
rect 67 240 68 242
rect 64 238 68 240
rect 73 244 79 245
rect 73 242 75 244
rect 77 242 79 244
rect 73 233 79 242
rect 111 243 135 247
rect 154 243 158 247
rect 195 282 199 284
rect 204 283 229 284
rect 204 281 206 283
rect 208 282 229 283
rect 208 281 226 282
rect 204 280 226 281
rect 228 280 229 282
rect 205 275 220 276
rect 205 274 216 275
rect 191 273 216 274
rect 218 273 220 275
rect 191 271 193 273
rect 195 272 220 273
rect 225 275 229 280
rect 234 282 244 283
rect 234 280 236 282
rect 238 280 244 282
rect 234 279 244 280
rect 225 273 226 275
rect 228 273 229 275
rect 195 271 209 272
rect 225 271 229 273
rect 191 270 209 271
rect 198 263 202 265
rect 198 261 199 263
rect 201 261 202 263
rect 198 251 202 261
rect 205 259 209 270
rect 240 275 244 279
rect 240 271 260 275
rect 256 268 260 271
rect 248 266 252 268
rect 248 264 249 266
rect 251 264 252 266
rect 248 259 252 264
rect 256 266 262 268
rect 256 264 259 266
rect 261 264 262 266
rect 256 262 262 264
rect 205 255 212 259
rect 208 254 212 255
rect 208 252 209 254
rect 211 252 212 254
rect 198 247 204 251
rect 208 250 212 252
rect 256 251 260 262
rect 220 250 260 251
rect 220 248 244 250
rect 246 248 260 250
rect 220 247 260 248
rect 200 243 224 247
rect 243 243 247 247
rect 283 282 289 289
rect 283 280 285 282
rect 287 280 289 282
rect 283 279 289 280
rect 294 280 298 282
rect 294 278 295 280
rect 297 278 298 280
rect 294 276 298 278
rect 303 280 309 289
rect 374 286 378 289
rect 430 287 432 289
rect 434 287 436 289
rect 430 286 436 287
rect 463 286 467 289
rect 519 287 521 289
rect 523 287 525 289
rect 519 286 525 287
rect 374 284 375 286
rect 377 284 378 286
rect 463 284 464 286
rect 466 284 467 286
rect 303 278 305 280
rect 307 278 309 280
rect 321 282 341 283
rect 321 280 323 282
rect 325 280 341 282
rect 321 279 341 280
rect 303 277 309 278
rect 281 272 298 276
rect 281 266 285 272
rect 281 264 282 266
rect 284 264 285 266
rect 281 251 285 264
rect 304 252 305 268
rect 337 275 341 279
rect 352 276 353 278
rect 337 271 349 275
rect 345 266 349 271
rect 345 264 346 266
rect 348 264 349 266
rect 277 244 278 250
rect 281 247 293 251
rect 141 242 147 243
rect 141 240 143 242
rect 145 240 147 242
rect 106 235 112 236
rect 106 233 108 235
rect 110 233 112 235
rect 141 235 147 240
rect 154 241 155 243
rect 157 241 158 243
rect 154 239 158 241
rect 163 242 169 243
rect 163 240 165 242
rect 167 240 169 242
rect 141 233 143 235
rect 145 233 147 235
rect 163 235 169 240
rect 230 242 236 243
rect 230 240 232 242
rect 234 240 236 242
rect 163 233 165 235
rect 167 233 169 235
rect 195 235 201 236
rect 195 233 197 235
rect 199 233 201 235
rect 230 235 236 240
rect 243 241 244 243
rect 246 241 247 243
rect 243 239 247 241
rect 252 242 258 243
rect 252 240 254 242
rect 256 240 258 242
rect 230 233 232 235
rect 234 233 236 235
rect 252 235 258 240
rect 289 242 293 247
rect 345 252 349 264
rect 332 249 349 252
rect 332 247 333 249
rect 335 248 349 249
rect 335 247 336 248
rect 321 242 327 243
rect 289 241 309 242
rect 289 239 305 241
rect 307 239 309 241
rect 289 238 309 239
rect 321 240 323 242
rect 325 240 327 242
rect 252 233 254 235
rect 256 233 258 235
rect 321 233 327 240
rect 332 242 336 247
rect 374 282 378 284
rect 383 283 408 284
rect 383 281 385 283
rect 387 282 408 283
rect 387 281 405 282
rect 383 280 405 281
rect 407 280 408 282
rect 384 275 399 276
rect 384 274 395 275
rect 370 273 395 274
rect 397 273 399 275
rect 370 271 372 273
rect 374 272 399 273
rect 404 275 408 280
rect 413 282 423 283
rect 413 280 415 282
rect 417 280 423 282
rect 413 279 423 280
rect 404 273 405 275
rect 407 273 408 275
rect 374 271 388 272
rect 404 271 408 273
rect 370 270 388 271
rect 377 263 381 265
rect 377 261 378 263
rect 380 261 381 263
rect 377 251 381 261
rect 384 259 388 270
rect 419 275 423 279
rect 419 271 439 275
rect 435 268 439 271
rect 427 266 431 268
rect 427 264 428 266
rect 430 264 431 266
rect 427 259 431 264
rect 435 266 441 268
rect 435 264 438 266
rect 440 264 441 266
rect 435 262 441 264
rect 384 255 391 259
rect 387 254 391 255
rect 387 252 388 254
rect 390 252 391 254
rect 377 247 383 251
rect 387 250 391 252
rect 435 251 439 262
rect 399 250 439 251
rect 399 248 423 250
rect 425 248 439 250
rect 399 247 439 248
rect 332 240 333 242
rect 335 240 336 242
rect 332 238 336 240
rect 341 244 347 245
rect 341 242 343 244
rect 345 242 347 244
rect 341 233 347 242
rect 379 243 403 247
rect 422 243 426 247
rect 463 282 467 284
rect 472 283 497 284
rect 472 281 474 283
rect 476 282 497 283
rect 476 281 494 282
rect 472 280 494 281
rect 496 280 497 282
rect 473 275 488 276
rect 473 274 484 275
rect 459 273 484 274
rect 486 273 488 275
rect 459 271 461 273
rect 463 272 488 273
rect 493 275 497 280
rect 502 282 512 283
rect 502 280 504 282
rect 506 280 512 282
rect 502 279 512 280
rect 493 273 494 275
rect 496 273 497 275
rect 463 271 477 272
rect 493 271 497 273
rect 459 270 477 271
rect 466 263 470 265
rect 466 261 467 263
rect 469 261 470 263
rect 466 251 470 261
rect 473 259 477 270
rect 508 275 512 279
rect 508 271 528 275
rect 524 268 528 271
rect 516 266 520 268
rect 516 264 517 266
rect 519 264 520 266
rect 516 259 520 264
rect 524 266 530 268
rect 524 264 527 266
rect 529 264 530 266
rect 524 262 530 264
rect 473 255 480 259
rect 476 254 480 255
rect 476 252 477 254
rect 479 252 480 254
rect 466 247 472 251
rect 476 250 480 252
rect 524 251 528 262
rect 488 250 528 251
rect 488 248 512 250
rect 514 248 528 250
rect 488 247 528 248
rect 468 243 492 247
rect 511 243 515 247
rect 551 282 557 289
rect 551 280 553 282
rect 555 280 557 282
rect 551 279 557 280
rect 562 280 566 282
rect 562 278 563 280
rect 565 278 566 280
rect 562 276 566 278
rect 571 280 577 289
rect 641 286 645 289
rect 697 287 699 289
rect 701 287 703 289
rect 697 286 703 287
rect 730 286 734 289
rect 786 287 788 289
rect 790 287 792 289
rect 786 286 792 287
rect 641 284 642 286
rect 644 284 645 286
rect 730 284 731 286
rect 733 284 734 286
rect 571 278 573 280
rect 575 278 577 280
rect 589 282 609 283
rect 589 280 591 282
rect 593 280 609 282
rect 589 279 609 280
rect 571 277 577 278
rect 549 272 566 276
rect 549 266 553 272
rect 549 264 550 266
rect 552 264 553 266
rect 549 251 553 264
rect 572 252 573 268
rect 605 275 609 279
rect 620 276 621 278
rect 605 271 617 275
rect 613 266 617 271
rect 613 264 614 266
rect 616 264 617 266
rect 545 244 546 250
rect 549 247 561 251
rect 409 242 415 243
rect 409 240 411 242
rect 413 240 415 242
rect 374 235 380 236
rect 374 233 376 235
rect 378 233 380 235
rect 409 235 415 240
rect 422 241 423 243
rect 425 241 426 243
rect 422 239 426 241
rect 431 242 437 243
rect 431 240 433 242
rect 435 240 437 242
rect 409 233 411 235
rect 413 233 415 235
rect 431 235 437 240
rect 498 242 504 243
rect 498 240 500 242
rect 502 240 504 242
rect 431 233 433 235
rect 435 233 437 235
rect 463 235 469 236
rect 463 233 465 235
rect 467 233 469 235
rect 498 235 504 240
rect 511 241 512 243
rect 514 241 515 243
rect 511 239 515 241
rect 520 242 526 243
rect 520 240 522 242
rect 524 240 526 242
rect 498 233 500 235
rect 502 233 504 235
rect 520 235 526 240
rect 557 242 561 247
rect 613 252 617 264
rect 600 249 617 252
rect 600 247 601 249
rect 603 248 617 249
rect 603 247 604 248
rect 589 242 595 243
rect 557 241 577 242
rect 557 239 573 241
rect 575 239 577 241
rect 557 238 577 239
rect 589 240 591 242
rect 593 240 595 242
rect 520 233 522 235
rect 524 233 526 235
rect 589 233 595 240
rect 600 242 604 247
rect 641 282 645 284
rect 650 283 675 284
rect 650 281 652 283
rect 654 282 675 283
rect 654 281 672 282
rect 650 280 672 281
rect 674 280 675 282
rect 651 275 666 276
rect 651 274 662 275
rect 637 273 662 274
rect 664 273 666 275
rect 637 271 639 273
rect 641 272 666 273
rect 671 275 675 280
rect 680 282 690 283
rect 680 280 682 282
rect 684 280 690 282
rect 680 279 690 280
rect 671 273 672 275
rect 674 273 675 275
rect 641 271 655 272
rect 671 271 675 273
rect 637 270 655 271
rect 644 263 648 265
rect 644 261 645 263
rect 647 261 648 263
rect 644 251 648 261
rect 651 259 655 270
rect 686 275 690 279
rect 686 271 706 275
rect 702 268 706 271
rect 694 266 698 268
rect 694 264 695 266
rect 697 264 698 266
rect 694 259 698 264
rect 702 266 708 268
rect 702 264 705 266
rect 707 264 708 266
rect 702 262 708 264
rect 651 255 658 259
rect 654 254 658 255
rect 654 252 655 254
rect 657 252 658 254
rect 644 247 650 251
rect 654 250 658 252
rect 702 251 706 262
rect 666 250 706 251
rect 666 248 690 250
rect 692 248 706 250
rect 666 247 706 248
rect 600 240 601 242
rect 603 240 604 242
rect 600 238 604 240
rect 609 244 615 245
rect 609 242 611 244
rect 613 242 615 244
rect 609 233 615 242
rect 646 243 670 247
rect 689 243 693 247
rect 730 282 734 284
rect 739 283 764 284
rect 739 281 741 283
rect 743 282 764 283
rect 743 281 761 282
rect 739 280 761 281
rect 763 280 764 282
rect 740 275 755 276
rect 740 274 751 275
rect 726 273 751 274
rect 753 273 755 275
rect 726 271 728 273
rect 730 272 755 273
rect 760 275 764 280
rect 769 282 779 283
rect 769 280 771 282
rect 773 280 779 282
rect 769 279 779 280
rect 760 273 761 275
rect 763 273 764 275
rect 730 271 744 272
rect 760 271 764 273
rect 726 270 744 271
rect 733 263 737 265
rect 733 261 734 263
rect 736 261 737 263
rect 733 251 737 261
rect 740 259 744 270
rect 775 275 779 279
rect 775 271 795 275
rect 791 268 795 271
rect 783 266 787 268
rect 783 264 784 266
rect 786 264 787 266
rect 783 259 787 264
rect 791 266 797 268
rect 791 264 794 266
rect 796 264 797 266
rect 791 262 797 264
rect 740 255 747 259
rect 743 254 747 255
rect 743 252 744 254
rect 746 252 747 254
rect 733 247 739 251
rect 743 250 747 252
rect 791 251 795 262
rect 755 250 795 251
rect 755 248 779 250
rect 781 248 795 250
rect 755 247 795 248
rect 735 243 759 247
rect 778 243 782 247
rect 818 282 824 289
rect 818 280 820 282
rect 822 280 824 282
rect 818 279 824 280
rect 829 280 833 282
rect 829 278 830 280
rect 832 278 833 280
rect 829 276 833 278
rect 838 280 844 289
rect 838 278 840 280
rect 842 278 844 280
rect 838 277 844 278
rect 816 272 833 276
rect 816 266 820 272
rect 816 264 817 266
rect 819 264 820 266
rect 816 251 820 264
rect 839 252 840 268
rect 812 244 813 250
rect 816 247 828 251
rect 676 242 682 243
rect 676 240 678 242
rect 680 240 682 242
rect 641 235 647 236
rect 641 233 643 235
rect 645 233 647 235
rect 676 235 682 240
rect 689 241 690 243
rect 692 241 693 243
rect 689 239 693 241
rect 698 242 704 243
rect 698 240 700 242
rect 702 240 704 242
rect 676 233 678 235
rect 680 233 682 235
rect 698 235 704 240
rect 765 242 771 243
rect 765 240 767 242
rect 769 240 771 242
rect 698 233 700 235
rect 702 233 704 235
rect 730 235 736 236
rect 730 233 732 235
rect 734 233 736 235
rect 765 235 771 240
rect 778 241 779 243
rect 781 241 782 243
rect 778 239 782 241
rect 787 242 793 243
rect 787 240 789 242
rect 791 240 793 242
rect 765 233 767 235
rect 769 233 771 235
rect 787 235 793 240
rect 824 242 828 247
rect 824 241 844 242
rect 824 239 840 241
rect 842 239 844 241
rect 824 238 844 239
rect 787 233 789 235
rect 791 233 793 235
rect 13 210 19 217
rect 13 208 15 210
rect 17 208 19 210
rect 13 207 19 208
rect 24 210 28 212
rect 24 208 25 210
rect 27 208 28 210
rect 24 203 28 208
rect 33 208 39 217
rect 33 206 35 208
rect 37 206 39 208
rect 53 210 59 217
rect 53 208 55 210
rect 57 208 59 210
rect 53 207 59 208
rect 64 210 68 212
rect 64 208 65 210
rect 67 208 68 210
rect 33 205 39 206
rect 24 201 25 203
rect 27 202 28 203
rect 27 201 41 202
rect 24 198 41 201
rect 37 186 41 198
rect 37 184 38 186
rect 40 184 41 186
rect 37 179 41 184
rect 29 175 41 179
rect 64 203 68 208
rect 73 208 79 217
rect 106 215 108 217
rect 110 215 112 217
rect 106 214 112 215
rect 141 215 143 217
rect 145 215 147 217
rect 73 206 75 208
rect 77 206 79 208
rect 73 205 79 206
rect 141 210 147 215
rect 163 215 165 217
rect 167 215 169 217
rect 141 208 143 210
rect 145 208 147 210
rect 141 207 147 208
rect 154 209 158 211
rect 154 207 155 209
rect 157 207 158 209
rect 163 210 169 215
rect 195 215 197 217
rect 199 215 201 217
rect 195 214 201 215
rect 230 215 232 217
rect 234 215 236 217
rect 163 208 165 210
rect 167 208 169 210
rect 163 207 169 208
rect 230 210 236 215
rect 252 215 254 217
rect 256 215 258 217
rect 230 208 232 210
rect 234 208 236 210
rect 230 207 236 208
rect 243 209 247 211
rect 243 207 244 209
rect 246 207 247 209
rect 252 210 258 215
rect 252 208 254 210
rect 256 208 258 210
rect 252 207 258 208
rect 64 201 65 203
rect 67 202 68 203
rect 67 201 81 202
rect 64 198 81 201
rect 29 171 33 175
rect 44 172 45 174
rect 77 186 81 198
rect 77 184 78 186
rect 80 184 81 186
rect 77 179 81 184
rect 69 175 81 179
rect 13 170 33 171
rect 13 168 15 170
rect 17 168 33 170
rect 13 167 33 168
rect 69 171 73 175
rect 84 172 85 174
rect 53 170 73 171
rect 53 168 55 170
rect 57 168 73 170
rect 53 167 73 168
rect 111 203 135 207
rect 154 203 158 207
rect 109 199 115 203
rect 131 202 171 203
rect 131 200 155 202
rect 157 200 171 202
rect 109 189 113 199
rect 119 198 123 200
rect 131 199 171 200
rect 119 196 120 198
rect 122 196 123 198
rect 119 195 123 196
rect 109 187 110 189
rect 112 187 113 189
rect 109 185 113 187
rect 116 191 123 195
rect 116 180 120 191
rect 159 186 163 191
rect 159 184 160 186
rect 162 184 163 186
rect 102 179 120 180
rect 102 177 104 179
rect 106 178 120 179
rect 106 177 131 178
rect 102 176 127 177
rect 116 175 127 176
rect 129 175 131 177
rect 116 174 131 175
rect 136 177 140 179
rect 136 175 137 177
rect 139 175 140 177
rect 136 170 140 175
rect 159 182 163 184
rect 167 188 171 199
rect 167 186 173 188
rect 167 184 170 186
rect 172 184 173 186
rect 167 182 173 184
rect 167 179 171 182
rect 151 175 171 179
rect 151 171 155 175
rect 115 169 137 170
rect 106 166 110 168
rect 115 167 117 169
rect 119 168 137 169
rect 139 168 140 170
rect 119 167 140 168
rect 145 170 155 171
rect 145 168 147 170
rect 149 168 155 170
rect 145 167 155 168
rect 200 203 224 207
rect 243 203 247 207
rect 289 211 309 212
rect 289 209 305 211
rect 307 209 309 211
rect 289 208 309 209
rect 321 210 327 217
rect 321 208 323 210
rect 325 208 327 210
rect 198 199 204 203
rect 220 202 260 203
rect 220 200 244 202
rect 246 200 260 202
rect 198 189 202 199
rect 208 198 212 200
rect 220 199 260 200
rect 208 196 209 198
rect 211 196 212 198
rect 208 195 212 196
rect 198 187 199 189
rect 201 187 202 189
rect 198 185 202 187
rect 205 191 212 195
rect 205 180 209 191
rect 248 186 252 191
rect 248 184 249 186
rect 251 184 252 186
rect 191 179 209 180
rect 191 177 193 179
rect 195 178 209 179
rect 195 177 220 178
rect 191 176 216 177
rect 205 175 216 176
rect 218 175 220 177
rect 205 174 220 175
rect 225 177 229 179
rect 225 175 226 177
rect 228 175 229 177
rect 225 170 229 175
rect 248 182 252 184
rect 256 188 260 199
rect 256 186 262 188
rect 256 184 259 186
rect 261 184 262 186
rect 256 182 262 184
rect 256 179 260 182
rect 240 175 260 179
rect 240 171 244 175
rect 204 169 226 170
rect 115 166 140 167
rect 195 166 199 168
rect 204 167 206 169
rect 208 168 226 169
rect 228 168 229 170
rect 208 167 229 168
rect 234 170 244 171
rect 234 168 236 170
rect 238 168 244 170
rect 234 167 244 168
rect 277 200 278 206
rect 289 203 293 208
rect 321 207 327 208
rect 332 210 336 212
rect 332 208 333 210
rect 335 208 336 210
rect 281 199 293 203
rect 281 186 285 199
rect 281 184 282 186
rect 284 184 285 186
rect 281 178 285 184
rect 304 182 305 198
rect 332 203 336 208
rect 341 208 347 217
rect 374 215 376 217
rect 378 215 380 217
rect 374 214 380 215
rect 409 215 411 217
rect 413 215 415 217
rect 341 206 343 208
rect 345 206 347 208
rect 341 205 347 206
rect 409 210 415 215
rect 431 215 433 217
rect 435 215 437 217
rect 409 208 411 210
rect 413 208 415 210
rect 409 207 415 208
rect 422 209 426 211
rect 422 207 423 209
rect 425 207 426 209
rect 431 210 437 215
rect 463 215 465 217
rect 467 215 469 217
rect 463 214 469 215
rect 498 215 500 217
rect 502 215 504 217
rect 431 208 433 210
rect 435 208 437 210
rect 431 207 437 208
rect 498 210 504 215
rect 520 215 522 217
rect 524 215 526 217
rect 498 208 500 210
rect 502 208 504 210
rect 498 207 504 208
rect 511 209 515 211
rect 511 207 512 209
rect 514 207 515 209
rect 520 210 526 215
rect 520 208 522 210
rect 524 208 526 210
rect 520 207 526 208
rect 332 201 333 203
rect 335 202 336 203
rect 335 201 349 202
rect 332 198 349 201
rect 345 186 349 198
rect 345 184 346 186
rect 348 184 349 186
rect 281 174 298 178
rect 345 179 349 184
rect 337 175 349 179
rect 294 172 298 174
rect 204 166 229 167
rect 283 170 289 171
rect 283 168 285 170
rect 287 168 289 170
rect 294 170 295 172
rect 297 170 298 172
rect 294 168 298 170
rect 303 172 309 173
rect 303 170 305 172
rect 307 170 309 172
rect 337 171 341 175
rect 352 172 353 174
rect 106 164 107 166
rect 109 164 110 166
rect 195 164 196 166
rect 198 164 199 166
rect 106 161 110 164
rect 162 163 168 164
rect 162 161 164 163
rect 166 161 168 163
rect 195 161 199 164
rect 251 163 257 164
rect 251 161 253 163
rect 255 161 257 163
rect 283 161 289 168
rect 303 161 309 170
rect 321 170 341 171
rect 321 168 323 170
rect 325 168 341 170
rect 321 167 341 168
rect 379 203 403 207
rect 422 203 426 207
rect 377 199 383 203
rect 399 202 439 203
rect 399 200 423 202
rect 425 200 439 202
rect 377 189 381 199
rect 387 198 391 200
rect 399 199 439 200
rect 387 196 388 198
rect 390 196 391 198
rect 387 195 391 196
rect 377 187 378 189
rect 380 187 381 189
rect 377 185 381 187
rect 384 191 391 195
rect 384 180 388 191
rect 427 186 431 191
rect 427 184 428 186
rect 430 184 431 186
rect 370 179 388 180
rect 370 177 372 179
rect 374 178 388 179
rect 374 177 399 178
rect 370 176 395 177
rect 384 175 395 176
rect 397 175 399 177
rect 384 174 399 175
rect 404 177 408 179
rect 404 175 405 177
rect 407 175 408 177
rect 404 170 408 175
rect 427 182 431 184
rect 435 188 439 199
rect 435 186 441 188
rect 435 184 438 186
rect 440 184 441 186
rect 435 182 441 184
rect 435 179 439 182
rect 419 175 439 179
rect 419 171 423 175
rect 383 169 405 170
rect 374 166 378 168
rect 383 167 385 169
rect 387 168 405 169
rect 407 168 408 170
rect 387 167 408 168
rect 413 170 423 171
rect 413 168 415 170
rect 417 168 423 170
rect 413 167 423 168
rect 468 203 492 207
rect 511 203 515 207
rect 557 211 577 212
rect 557 209 573 211
rect 575 209 577 211
rect 557 208 577 209
rect 589 210 595 217
rect 589 208 591 210
rect 593 208 595 210
rect 466 199 472 203
rect 488 202 528 203
rect 488 200 512 202
rect 514 200 528 202
rect 466 189 470 199
rect 476 198 480 200
rect 488 199 528 200
rect 476 196 477 198
rect 479 196 480 198
rect 476 195 480 196
rect 466 187 467 189
rect 469 187 470 189
rect 466 185 470 187
rect 473 191 480 195
rect 473 180 477 191
rect 516 186 520 191
rect 516 184 517 186
rect 519 184 520 186
rect 459 179 477 180
rect 459 177 461 179
rect 463 178 477 179
rect 463 177 488 178
rect 459 176 484 177
rect 473 175 484 176
rect 486 175 488 177
rect 473 174 488 175
rect 493 177 497 179
rect 493 175 494 177
rect 496 175 497 177
rect 493 170 497 175
rect 516 182 520 184
rect 524 188 528 199
rect 524 186 530 188
rect 524 184 527 186
rect 529 184 530 186
rect 524 182 530 184
rect 524 179 528 182
rect 508 175 528 179
rect 508 171 512 175
rect 472 169 494 170
rect 383 166 408 167
rect 463 166 467 168
rect 472 167 474 169
rect 476 168 494 169
rect 496 168 497 170
rect 476 167 497 168
rect 502 170 512 171
rect 502 168 504 170
rect 506 168 512 170
rect 502 167 512 168
rect 545 200 546 206
rect 557 203 561 208
rect 589 207 595 208
rect 600 210 604 212
rect 600 208 601 210
rect 603 208 604 210
rect 549 199 561 203
rect 549 186 553 199
rect 549 184 550 186
rect 552 184 553 186
rect 549 178 553 184
rect 572 182 573 198
rect 600 203 604 208
rect 609 208 615 217
rect 641 215 643 217
rect 645 215 647 217
rect 641 214 647 215
rect 676 215 678 217
rect 680 215 682 217
rect 609 206 611 208
rect 613 206 615 208
rect 609 205 615 206
rect 676 210 682 215
rect 698 215 700 217
rect 702 215 704 217
rect 676 208 678 210
rect 680 208 682 210
rect 676 207 682 208
rect 689 209 693 211
rect 689 207 690 209
rect 692 207 693 209
rect 698 210 704 215
rect 730 215 732 217
rect 734 215 736 217
rect 730 214 736 215
rect 765 215 767 217
rect 769 215 771 217
rect 698 208 700 210
rect 702 208 704 210
rect 698 207 704 208
rect 765 210 771 215
rect 787 215 789 217
rect 791 215 793 217
rect 765 208 767 210
rect 769 208 771 210
rect 765 207 771 208
rect 778 209 782 211
rect 778 207 779 209
rect 781 207 782 209
rect 787 210 793 215
rect 787 208 789 210
rect 791 208 793 210
rect 787 207 793 208
rect 600 201 601 203
rect 603 202 604 203
rect 603 201 617 202
rect 600 198 617 201
rect 613 186 617 198
rect 613 184 614 186
rect 616 184 617 186
rect 549 174 566 178
rect 613 179 617 184
rect 605 175 617 179
rect 562 172 566 174
rect 472 166 497 167
rect 551 170 557 171
rect 551 168 553 170
rect 555 168 557 170
rect 562 170 563 172
rect 565 170 566 172
rect 562 168 566 170
rect 571 172 577 173
rect 571 170 573 172
rect 575 170 577 172
rect 605 171 609 175
rect 620 172 621 174
rect 374 164 375 166
rect 377 164 378 166
rect 463 164 464 166
rect 466 164 467 166
rect 374 161 378 164
rect 430 163 436 164
rect 430 161 432 163
rect 434 161 436 163
rect 463 161 467 164
rect 519 163 525 164
rect 519 161 521 163
rect 523 161 525 163
rect 551 161 557 168
rect 571 161 577 170
rect 589 170 609 171
rect 589 168 591 170
rect 593 168 609 170
rect 589 167 609 168
rect 646 203 670 207
rect 689 203 693 207
rect 644 199 650 203
rect 666 202 706 203
rect 666 200 690 202
rect 692 200 706 202
rect 644 189 648 199
rect 654 198 658 200
rect 666 199 706 200
rect 654 196 655 198
rect 657 196 658 198
rect 654 195 658 196
rect 644 187 645 189
rect 647 187 648 189
rect 644 185 648 187
rect 651 191 658 195
rect 651 180 655 191
rect 694 186 698 191
rect 694 184 695 186
rect 697 184 698 186
rect 637 179 655 180
rect 637 177 639 179
rect 641 178 655 179
rect 641 177 666 178
rect 637 176 662 177
rect 651 175 662 176
rect 664 175 666 177
rect 651 174 666 175
rect 671 177 675 179
rect 671 175 672 177
rect 674 175 675 177
rect 671 170 675 175
rect 694 182 698 184
rect 702 188 706 199
rect 702 186 708 188
rect 702 184 705 186
rect 707 184 708 186
rect 702 182 708 184
rect 702 179 706 182
rect 686 175 706 179
rect 686 171 690 175
rect 650 169 672 170
rect 641 166 645 168
rect 650 167 652 169
rect 654 168 672 169
rect 674 168 675 170
rect 654 167 675 168
rect 680 170 690 171
rect 680 168 682 170
rect 684 168 690 170
rect 680 167 690 168
rect 735 203 759 207
rect 778 203 782 207
rect 824 211 844 212
rect 824 209 840 211
rect 842 209 844 211
rect 824 208 844 209
rect 733 199 739 203
rect 755 202 795 203
rect 755 200 779 202
rect 781 200 795 202
rect 733 189 737 199
rect 743 198 747 200
rect 755 199 795 200
rect 743 196 744 198
rect 746 196 747 198
rect 743 195 747 196
rect 733 187 734 189
rect 736 187 737 189
rect 733 185 737 187
rect 740 191 747 195
rect 740 180 744 191
rect 783 186 787 191
rect 783 184 784 186
rect 786 184 787 186
rect 726 179 744 180
rect 726 177 728 179
rect 730 178 744 179
rect 730 177 755 178
rect 726 176 751 177
rect 740 175 751 176
rect 753 175 755 177
rect 740 174 755 175
rect 760 177 764 179
rect 760 175 761 177
rect 763 175 764 177
rect 760 170 764 175
rect 783 182 787 184
rect 791 188 795 199
rect 791 186 797 188
rect 791 184 794 186
rect 796 184 797 186
rect 791 182 797 184
rect 791 179 795 182
rect 775 175 795 179
rect 775 171 779 175
rect 739 169 761 170
rect 650 166 675 167
rect 730 166 734 168
rect 739 167 741 169
rect 743 168 761 169
rect 763 168 764 170
rect 743 167 764 168
rect 769 170 779 171
rect 769 168 771 170
rect 773 168 779 170
rect 769 167 779 168
rect 812 200 813 206
rect 824 203 828 208
rect 816 199 828 203
rect 816 186 820 199
rect 816 184 817 186
rect 819 184 820 186
rect 816 178 820 184
rect 839 182 840 198
rect 816 174 833 178
rect 829 172 833 174
rect 739 166 764 167
rect 818 170 824 171
rect 818 168 820 170
rect 822 168 824 170
rect 829 170 830 172
rect 832 170 833 172
rect 829 168 833 170
rect 838 172 844 173
rect 838 170 840 172
rect 842 170 844 172
rect 641 164 642 166
rect 644 164 645 166
rect 730 164 731 166
rect 733 164 734 166
rect 641 161 645 164
rect 697 163 703 164
rect 697 161 699 163
rect 701 161 703 163
rect 730 161 734 164
rect 786 163 792 164
rect 786 161 788 163
rect 790 161 792 163
rect 818 161 824 168
rect 838 161 844 170
rect 106 142 110 145
rect 162 143 164 145
rect 166 143 168 145
rect 162 142 168 143
rect 195 142 199 145
rect 251 143 253 145
rect 255 143 257 145
rect 251 142 257 143
rect 106 140 107 142
rect 109 140 110 142
rect 195 140 196 142
rect 198 140 199 142
rect 13 138 33 139
rect 13 136 15 138
rect 17 136 33 138
rect 13 135 33 136
rect 29 131 33 135
rect 53 138 73 139
rect 53 136 55 138
rect 57 136 73 138
rect 53 135 73 136
rect 44 132 45 134
rect 29 127 41 131
rect 37 122 41 127
rect 37 120 38 122
rect 40 120 41 122
rect 37 108 41 120
rect 69 131 73 135
rect 84 132 85 134
rect 69 127 81 131
rect 77 122 81 127
rect 77 120 78 122
rect 80 120 81 122
rect 24 105 41 108
rect 24 103 25 105
rect 27 104 41 105
rect 27 103 28 104
rect 13 98 19 99
rect 13 96 15 98
rect 17 96 19 98
rect 13 89 19 96
rect 24 98 28 103
rect 77 108 81 120
rect 64 105 81 108
rect 64 103 65 105
rect 67 104 81 105
rect 67 103 68 104
rect 24 96 25 98
rect 27 96 28 98
rect 24 94 28 96
rect 33 100 39 101
rect 33 98 35 100
rect 37 98 39 100
rect 33 89 39 98
rect 53 98 59 99
rect 53 96 55 98
rect 57 96 59 98
rect 53 89 59 96
rect 64 98 68 103
rect 106 138 110 140
rect 115 139 140 140
rect 115 137 117 139
rect 119 138 140 139
rect 119 137 137 138
rect 115 136 137 137
rect 139 136 140 138
rect 116 131 131 132
rect 116 130 127 131
rect 102 129 127 130
rect 129 129 131 131
rect 102 127 104 129
rect 106 128 131 129
rect 136 131 140 136
rect 145 138 155 139
rect 145 136 147 138
rect 149 136 155 138
rect 145 135 155 136
rect 136 129 137 131
rect 139 129 140 131
rect 106 127 120 128
rect 136 127 140 129
rect 102 126 120 127
rect 109 119 113 121
rect 109 117 110 119
rect 112 117 113 119
rect 109 107 113 117
rect 116 115 120 126
rect 151 131 155 135
rect 151 127 171 131
rect 167 124 171 127
rect 159 122 163 124
rect 159 120 160 122
rect 162 120 163 122
rect 159 115 163 120
rect 167 122 173 124
rect 167 120 170 122
rect 172 120 173 122
rect 167 118 173 120
rect 116 111 123 115
rect 119 110 123 111
rect 119 108 120 110
rect 122 108 123 110
rect 109 103 115 107
rect 119 106 123 108
rect 167 107 171 118
rect 131 106 171 107
rect 131 104 155 106
rect 157 104 171 106
rect 131 103 171 104
rect 64 96 65 98
rect 67 96 68 98
rect 64 94 68 96
rect 73 100 79 101
rect 73 98 75 100
rect 77 98 79 100
rect 73 89 79 98
rect 111 99 135 103
rect 154 99 158 103
rect 195 138 199 140
rect 204 139 229 140
rect 204 137 206 139
rect 208 138 229 139
rect 208 137 226 138
rect 204 136 226 137
rect 228 136 229 138
rect 205 131 220 132
rect 205 130 216 131
rect 191 129 216 130
rect 218 129 220 131
rect 191 127 193 129
rect 195 128 220 129
rect 225 131 229 136
rect 234 138 244 139
rect 234 136 236 138
rect 238 136 244 138
rect 234 135 244 136
rect 225 129 226 131
rect 228 129 229 131
rect 195 127 209 128
rect 225 127 229 129
rect 191 126 209 127
rect 198 119 202 121
rect 198 117 199 119
rect 201 117 202 119
rect 198 107 202 117
rect 205 115 209 126
rect 240 131 244 135
rect 240 127 260 131
rect 256 124 260 127
rect 248 122 252 124
rect 248 120 249 122
rect 251 120 252 122
rect 248 115 252 120
rect 256 122 262 124
rect 256 120 259 122
rect 261 120 262 122
rect 256 118 262 120
rect 205 111 212 115
rect 208 110 212 111
rect 208 108 209 110
rect 211 108 212 110
rect 198 103 204 107
rect 208 106 212 108
rect 256 107 260 118
rect 220 106 260 107
rect 220 104 244 106
rect 246 104 260 106
rect 220 103 260 104
rect 200 99 224 103
rect 243 99 247 103
rect 283 138 289 145
rect 283 136 285 138
rect 287 136 289 138
rect 283 135 289 136
rect 294 136 298 138
rect 294 134 295 136
rect 297 134 298 136
rect 294 132 298 134
rect 303 136 309 145
rect 374 142 378 145
rect 430 143 432 145
rect 434 143 436 145
rect 430 142 436 143
rect 463 142 467 145
rect 519 143 521 145
rect 523 143 525 145
rect 519 142 525 143
rect 374 140 375 142
rect 377 140 378 142
rect 463 140 464 142
rect 466 140 467 142
rect 303 134 305 136
rect 307 134 309 136
rect 321 138 341 139
rect 321 136 323 138
rect 325 136 341 138
rect 321 135 341 136
rect 303 133 309 134
rect 281 128 298 132
rect 281 122 285 128
rect 281 120 282 122
rect 284 120 285 122
rect 281 107 285 120
rect 304 108 305 124
rect 337 131 341 135
rect 352 132 353 134
rect 337 127 349 131
rect 345 122 349 127
rect 345 120 346 122
rect 348 120 349 122
rect 277 100 278 106
rect 281 103 293 107
rect 141 98 147 99
rect 141 96 143 98
rect 145 96 147 98
rect 106 91 112 92
rect 106 89 108 91
rect 110 89 112 91
rect 141 91 147 96
rect 154 97 155 99
rect 157 97 158 99
rect 154 95 158 97
rect 163 98 169 99
rect 163 96 165 98
rect 167 96 169 98
rect 141 89 143 91
rect 145 89 147 91
rect 163 91 169 96
rect 230 98 236 99
rect 230 96 232 98
rect 234 96 236 98
rect 163 89 165 91
rect 167 89 169 91
rect 195 91 201 92
rect 195 89 197 91
rect 199 89 201 91
rect 230 91 236 96
rect 243 97 244 99
rect 246 97 247 99
rect 243 95 247 97
rect 252 98 258 99
rect 252 96 254 98
rect 256 96 258 98
rect 230 89 232 91
rect 234 89 236 91
rect 252 91 258 96
rect 289 98 293 103
rect 345 108 349 120
rect 332 105 349 108
rect 332 103 333 105
rect 335 104 349 105
rect 335 103 336 104
rect 321 98 327 99
rect 289 97 309 98
rect 289 95 305 97
rect 307 95 309 97
rect 289 94 309 95
rect 321 96 323 98
rect 325 96 327 98
rect 252 89 254 91
rect 256 89 258 91
rect 321 89 327 96
rect 332 98 336 103
rect 374 138 378 140
rect 383 139 408 140
rect 383 137 385 139
rect 387 138 408 139
rect 387 137 405 138
rect 383 136 405 137
rect 407 136 408 138
rect 384 131 399 132
rect 384 130 395 131
rect 370 129 395 130
rect 397 129 399 131
rect 370 127 372 129
rect 374 128 399 129
rect 404 131 408 136
rect 413 138 423 139
rect 413 136 415 138
rect 417 136 423 138
rect 413 135 423 136
rect 404 129 405 131
rect 407 129 408 131
rect 374 127 388 128
rect 404 127 408 129
rect 370 126 388 127
rect 377 119 381 121
rect 377 117 378 119
rect 380 117 381 119
rect 377 107 381 117
rect 384 115 388 126
rect 419 131 423 135
rect 419 127 439 131
rect 435 124 439 127
rect 427 122 431 124
rect 427 120 428 122
rect 430 120 431 122
rect 427 115 431 120
rect 435 122 441 124
rect 435 120 438 122
rect 440 120 441 122
rect 435 118 441 120
rect 384 111 391 115
rect 387 110 391 111
rect 387 108 388 110
rect 390 108 391 110
rect 377 103 383 107
rect 387 106 391 108
rect 435 107 439 118
rect 399 106 439 107
rect 399 104 423 106
rect 425 104 439 106
rect 399 103 439 104
rect 332 96 333 98
rect 335 96 336 98
rect 332 94 336 96
rect 341 100 347 101
rect 341 98 343 100
rect 345 98 347 100
rect 341 89 347 98
rect 379 99 403 103
rect 422 99 426 103
rect 463 138 467 140
rect 472 139 497 140
rect 472 137 474 139
rect 476 138 497 139
rect 476 137 494 138
rect 472 136 494 137
rect 496 136 497 138
rect 473 131 488 132
rect 473 130 484 131
rect 459 129 484 130
rect 486 129 488 131
rect 459 127 461 129
rect 463 128 488 129
rect 493 131 497 136
rect 502 138 512 139
rect 502 136 504 138
rect 506 136 512 138
rect 502 135 512 136
rect 493 129 494 131
rect 496 129 497 131
rect 463 127 477 128
rect 493 127 497 129
rect 459 126 477 127
rect 466 119 470 121
rect 466 117 467 119
rect 469 117 470 119
rect 466 107 470 117
rect 473 115 477 126
rect 508 131 512 135
rect 508 127 528 131
rect 524 124 528 127
rect 516 122 520 124
rect 516 120 517 122
rect 519 120 520 122
rect 516 115 520 120
rect 524 122 530 124
rect 524 120 527 122
rect 529 120 530 122
rect 524 118 530 120
rect 473 111 480 115
rect 476 110 480 111
rect 476 108 477 110
rect 479 108 480 110
rect 466 103 472 107
rect 476 106 480 108
rect 524 107 528 118
rect 488 106 528 107
rect 488 104 512 106
rect 514 104 528 106
rect 488 103 528 104
rect 468 99 492 103
rect 511 99 515 103
rect 551 138 557 145
rect 551 136 553 138
rect 555 136 557 138
rect 551 135 557 136
rect 562 136 566 138
rect 562 134 563 136
rect 565 134 566 136
rect 562 132 566 134
rect 571 136 577 145
rect 641 142 645 145
rect 697 143 699 145
rect 701 143 703 145
rect 697 142 703 143
rect 730 142 734 145
rect 786 143 788 145
rect 790 143 792 145
rect 786 142 792 143
rect 641 140 642 142
rect 644 140 645 142
rect 730 140 731 142
rect 733 140 734 142
rect 571 134 573 136
rect 575 134 577 136
rect 589 138 609 139
rect 589 136 591 138
rect 593 136 609 138
rect 589 135 609 136
rect 571 133 577 134
rect 549 128 566 132
rect 549 122 553 128
rect 549 120 550 122
rect 552 120 553 122
rect 549 107 553 120
rect 572 108 573 124
rect 605 131 609 135
rect 620 132 621 134
rect 605 127 617 131
rect 613 122 617 127
rect 613 120 614 122
rect 616 120 617 122
rect 545 100 546 106
rect 549 103 561 107
rect 409 98 415 99
rect 409 96 411 98
rect 413 96 415 98
rect 374 91 380 92
rect 374 89 376 91
rect 378 89 380 91
rect 409 91 415 96
rect 422 97 423 99
rect 425 97 426 99
rect 422 95 426 97
rect 431 98 437 99
rect 431 96 433 98
rect 435 96 437 98
rect 409 89 411 91
rect 413 89 415 91
rect 431 91 437 96
rect 498 98 504 99
rect 498 96 500 98
rect 502 96 504 98
rect 431 89 433 91
rect 435 89 437 91
rect 463 91 469 92
rect 463 89 465 91
rect 467 89 469 91
rect 498 91 504 96
rect 511 97 512 99
rect 514 97 515 99
rect 511 95 515 97
rect 520 98 526 99
rect 520 96 522 98
rect 524 96 526 98
rect 498 89 500 91
rect 502 89 504 91
rect 520 91 526 96
rect 557 98 561 103
rect 613 108 617 120
rect 600 105 617 108
rect 600 103 601 105
rect 603 104 617 105
rect 603 103 604 104
rect 589 98 595 99
rect 557 97 577 98
rect 557 95 573 97
rect 575 95 577 97
rect 557 94 577 95
rect 589 96 591 98
rect 593 96 595 98
rect 520 89 522 91
rect 524 89 526 91
rect 589 89 595 96
rect 600 98 604 103
rect 641 138 645 140
rect 650 139 675 140
rect 650 137 652 139
rect 654 138 675 139
rect 654 137 672 138
rect 650 136 672 137
rect 674 136 675 138
rect 651 131 666 132
rect 651 130 662 131
rect 637 129 662 130
rect 664 129 666 131
rect 637 127 639 129
rect 641 128 666 129
rect 671 131 675 136
rect 680 138 690 139
rect 680 136 682 138
rect 684 136 690 138
rect 680 135 690 136
rect 671 129 672 131
rect 674 129 675 131
rect 641 127 655 128
rect 671 127 675 129
rect 637 126 655 127
rect 644 119 648 121
rect 644 117 645 119
rect 647 117 648 119
rect 644 107 648 117
rect 651 115 655 126
rect 686 131 690 135
rect 686 127 706 131
rect 702 124 706 127
rect 694 122 698 124
rect 694 120 695 122
rect 697 120 698 122
rect 694 115 698 120
rect 702 122 708 124
rect 702 120 705 122
rect 707 120 708 122
rect 702 118 708 120
rect 651 111 658 115
rect 654 110 658 111
rect 654 108 655 110
rect 657 108 658 110
rect 644 103 650 107
rect 654 106 658 108
rect 702 107 706 118
rect 666 106 706 107
rect 666 104 690 106
rect 692 104 706 106
rect 666 103 706 104
rect 600 96 601 98
rect 603 96 604 98
rect 600 94 604 96
rect 609 100 615 101
rect 609 98 611 100
rect 613 98 615 100
rect 609 89 615 98
rect 646 99 670 103
rect 689 99 693 103
rect 730 138 734 140
rect 739 139 764 140
rect 739 137 741 139
rect 743 138 764 139
rect 743 137 761 138
rect 739 136 761 137
rect 763 136 764 138
rect 740 131 755 132
rect 740 130 751 131
rect 726 129 751 130
rect 753 129 755 131
rect 726 127 728 129
rect 730 128 755 129
rect 760 131 764 136
rect 769 138 779 139
rect 769 136 771 138
rect 773 136 779 138
rect 769 135 779 136
rect 760 129 761 131
rect 763 129 764 131
rect 730 127 744 128
rect 760 127 764 129
rect 726 126 744 127
rect 733 119 737 121
rect 733 117 734 119
rect 736 117 737 119
rect 733 107 737 117
rect 740 115 744 126
rect 775 131 779 135
rect 775 127 795 131
rect 791 124 795 127
rect 783 122 787 124
rect 783 120 784 122
rect 786 120 787 122
rect 783 115 787 120
rect 791 122 797 124
rect 791 120 794 122
rect 796 120 797 122
rect 791 118 797 120
rect 740 111 747 115
rect 743 110 747 111
rect 743 108 744 110
rect 746 108 747 110
rect 733 103 739 107
rect 743 106 747 108
rect 791 107 795 118
rect 755 106 795 107
rect 755 104 779 106
rect 781 104 795 106
rect 755 103 795 104
rect 735 99 759 103
rect 778 99 782 103
rect 818 138 824 145
rect 818 136 820 138
rect 822 136 824 138
rect 818 135 824 136
rect 829 136 833 138
rect 829 134 830 136
rect 832 134 833 136
rect 829 132 833 134
rect 838 136 844 145
rect 838 134 840 136
rect 842 134 844 136
rect 838 133 844 134
rect 816 128 833 132
rect 816 122 820 128
rect 816 120 817 122
rect 819 120 820 122
rect 816 107 820 120
rect 839 108 840 124
rect 812 100 813 106
rect 816 103 828 107
rect 676 98 682 99
rect 676 96 678 98
rect 680 96 682 98
rect 641 91 647 92
rect 641 89 643 91
rect 645 89 647 91
rect 676 91 682 96
rect 689 97 690 99
rect 692 97 693 99
rect 689 95 693 97
rect 698 98 704 99
rect 698 96 700 98
rect 702 96 704 98
rect 676 89 678 91
rect 680 89 682 91
rect 698 91 704 96
rect 765 98 771 99
rect 765 96 767 98
rect 769 96 771 98
rect 698 89 700 91
rect 702 89 704 91
rect 730 91 736 92
rect 730 89 732 91
rect 734 89 736 91
rect 765 91 771 96
rect 778 97 779 99
rect 781 97 782 99
rect 778 95 782 97
rect 787 98 793 99
rect 787 96 789 98
rect 791 96 793 98
rect 765 89 767 91
rect 769 89 771 91
rect 787 91 793 96
rect 824 98 828 103
rect 824 97 844 98
rect 824 95 840 97
rect 842 95 844 97
rect 824 94 844 95
rect 787 89 789 91
rect 791 89 793 91
rect 13 66 19 73
rect 13 64 15 66
rect 17 64 19 66
rect 13 63 19 64
rect 24 66 28 68
rect 24 64 25 66
rect 27 64 28 66
rect 24 59 28 64
rect 33 64 39 73
rect 33 62 35 64
rect 37 62 39 64
rect 53 66 59 73
rect 53 64 55 66
rect 57 64 59 66
rect 53 63 59 64
rect 64 66 68 68
rect 64 64 65 66
rect 67 64 68 66
rect 33 61 39 62
rect 24 57 25 59
rect 27 58 28 59
rect 27 57 41 58
rect 24 54 41 57
rect 37 42 41 54
rect 37 40 38 42
rect 40 40 41 42
rect 37 35 41 40
rect 29 31 41 35
rect 64 59 68 64
rect 73 64 79 73
rect 106 71 108 73
rect 110 71 112 73
rect 106 70 112 71
rect 141 71 143 73
rect 145 71 147 73
rect 73 62 75 64
rect 77 62 79 64
rect 73 61 79 62
rect 141 66 147 71
rect 163 71 165 73
rect 167 71 169 73
rect 141 64 143 66
rect 145 64 147 66
rect 141 63 147 64
rect 154 65 158 67
rect 154 63 155 65
rect 157 63 158 65
rect 163 66 169 71
rect 195 71 197 73
rect 199 71 201 73
rect 195 70 201 71
rect 230 71 232 73
rect 234 71 236 73
rect 163 64 165 66
rect 167 64 169 66
rect 163 63 169 64
rect 230 66 236 71
rect 252 71 254 73
rect 256 71 258 73
rect 230 64 232 66
rect 234 64 236 66
rect 230 63 236 64
rect 243 65 247 67
rect 243 63 244 65
rect 246 63 247 65
rect 252 66 258 71
rect 252 64 254 66
rect 256 64 258 66
rect 252 63 258 64
rect 64 57 65 59
rect 67 58 68 59
rect 67 57 81 58
rect 64 54 81 57
rect 29 27 33 31
rect 44 28 45 30
rect 77 42 81 54
rect 77 40 78 42
rect 80 40 81 42
rect 77 35 81 40
rect 69 31 81 35
rect 13 26 33 27
rect 13 24 15 26
rect 17 24 33 26
rect 13 23 33 24
rect 69 27 73 31
rect 84 28 85 30
rect 53 26 73 27
rect 53 24 55 26
rect 57 24 73 26
rect 53 23 73 24
rect 111 59 135 63
rect 154 59 158 63
rect 109 55 115 59
rect 131 58 171 59
rect 131 56 155 58
rect 157 56 171 58
rect 109 45 113 55
rect 119 54 123 56
rect 131 55 171 56
rect 119 52 120 54
rect 122 52 123 54
rect 119 51 123 52
rect 109 43 110 45
rect 112 43 113 45
rect 109 41 113 43
rect 116 47 123 51
rect 116 36 120 47
rect 159 42 163 47
rect 159 40 160 42
rect 162 40 163 42
rect 102 35 120 36
rect 102 33 104 35
rect 106 34 120 35
rect 106 33 131 34
rect 102 32 127 33
rect 116 31 127 32
rect 129 31 131 33
rect 116 30 131 31
rect 136 33 140 35
rect 136 31 137 33
rect 139 31 140 33
rect 136 26 140 31
rect 159 38 163 40
rect 167 44 171 55
rect 167 42 173 44
rect 167 40 170 42
rect 172 40 173 42
rect 167 38 173 40
rect 167 35 171 38
rect 151 31 171 35
rect 151 27 155 31
rect 115 25 137 26
rect 106 22 110 24
rect 115 23 117 25
rect 119 24 137 25
rect 139 24 140 26
rect 119 23 140 24
rect 145 26 155 27
rect 145 24 147 26
rect 149 24 155 26
rect 145 23 155 24
rect 200 59 224 63
rect 243 59 247 63
rect 289 67 309 68
rect 289 65 305 67
rect 307 65 309 67
rect 289 64 309 65
rect 321 66 327 73
rect 321 64 323 66
rect 325 64 327 66
rect 198 55 204 59
rect 220 58 260 59
rect 220 56 244 58
rect 246 56 260 58
rect 198 45 202 55
rect 208 54 212 56
rect 220 55 260 56
rect 208 52 209 54
rect 211 52 212 54
rect 208 51 212 52
rect 198 43 199 45
rect 201 43 202 45
rect 198 41 202 43
rect 205 47 212 51
rect 205 36 209 47
rect 248 42 252 47
rect 248 40 249 42
rect 251 40 252 42
rect 191 35 209 36
rect 191 33 193 35
rect 195 34 209 35
rect 195 33 220 34
rect 191 32 216 33
rect 205 31 216 32
rect 218 31 220 33
rect 205 30 220 31
rect 225 33 229 35
rect 225 31 226 33
rect 228 31 229 33
rect 225 26 229 31
rect 248 38 252 40
rect 256 44 260 55
rect 256 42 262 44
rect 256 40 259 42
rect 261 40 262 42
rect 256 38 262 40
rect 256 35 260 38
rect 240 31 260 35
rect 240 27 244 31
rect 204 25 226 26
rect 115 22 140 23
rect 195 22 199 24
rect 204 23 206 25
rect 208 24 226 25
rect 228 24 229 26
rect 208 23 229 24
rect 234 26 244 27
rect 234 24 236 26
rect 238 24 244 26
rect 234 23 244 24
rect 277 56 278 62
rect 289 59 293 64
rect 321 63 327 64
rect 332 66 336 68
rect 332 64 333 66
rect 335 64 336 66
rect 281 55 293 59
rect 281 42 285 55
rect 281 40 282 42
rect 284 40 285 42
rect 281 34 285 40
rect 304 38 305 54
rect 332 59 336 64
rect 341 64 347 73
rect 374 71 376 73
rect 378 71 380 73
rect 374 70 380 71
rect 409 71 411 73
rect 413 71 415 73
rect 341 62 343 64
rect 345 62 347 64
rect 341 61 347 62
rect 409 66 415 71
rect 431 71 433 73
rect 435 71 437 73
rect 409 64 411 66
rect 413 64 415 66
rect 409 63 415 64
rect 422 65 426 67
rect 422 63 423 65
rect 425 63 426 65
rect 431 66 437 71
rect 463 71 465 73
rect 467 71 469 73
rect 463 70 469 71
rect 498 71 500 73
rect 502 71 504 73
rect 431 64 433 66
rect 435 64 437 66
rect 431 63 437 64
rect 498 66 504 71
rect 520 71 522 73
rect 524 71 526 73
rect 498 64 500 66
rect 502 64 504 66
rect 498 63 504 64
rect 511 65 515 67
rect 511 63 512 65
rect 514 63 515 65
rect 520 66 526 71
rect 520 64 522 66
rect 524 64 526 66
rect 520 63 526 64
rect 332 57 333 59
rect 335 58 336 59
rect 335 57 349 58
rect 332 54 349 57
rect 345 42 349 54
rect 345 40 346 42
rect 348 40 349 42
rect 281 30 298 34
rect 345 35 349 40
rect 337 31 349 35
rect 294 28 298 30
rect 204 22 229 23
rect 283 26 289 27
rect 283 24 285 26
rect 287 24 289 26
rect 294 26 295 28
rect 297 26 298 28
rect 294 24 298 26
rect 303 28 309 29
rect 303 26 305 28
rect 307 26 309 28
rect 337 27 341 31
rect 352 28 353 30
rect 106 20 107 22
rect 109 20 110 22
rect 195 20 196 22
rect 198 20 199 22
rect 106 17 110 20
rect 162 19 168 20
rect 162 17 164 19
rect 166 17 168 19
rect 195 17 199 20
rect 251 19 257 20
rect 251 17 253 19
rect 255 17 257 19
rect 283 17 289 24
rect 303 17 309 26
rect 321 26 341 27
rect 321 24 323 26
rect 325 24 341 26
rect 321 23 341 24
rect 379 59 403 63
rect 422 59 426 63
rect 377 55 383 59
rect 399 58 439 59
rect 399 56 423 58
rect 425 56 439 58
rect 377 45 381 55
rect 387 54 391 56
rect 399 55 439 56
rect 387 52 388 54
rect 390 52 391 54
rect 387 51 391 52
rect 377 43 378 45
rect 380 43 381 45
rect 377 41 381 43
rect 384 47 391 51
rect 384 36 388 47
rect 427 42 431 47
rect 427 40 428 42
rect 430 40 431 42
rect 370 35 388 36
rect 370 33 372 35
rect 374 34 388 35
rect 374 33 399 34
rect 370 32 395 33
rect 384 31 395 32
rect 397 31 399 33
rect 384 30 399 31
rect 404 33 408 35
rect 404 31 405 33
rect 407 31 408 33
rect 404 26 408 31
rect 427 38 431 40
rect 435 44 439 55
rect 435 42 441 44
rect 435 40 438 42
rect 440 40 441 42
rect 435 38 441 40
rect 435 35 439 38
rect 419 31 439 35
rect 419 27 423 31
rect 383 25 405 26
rect 374 22 378 24
rect 383 23 385 25
rect 387 24 405 25
rect 407 24 408 26
rect 387 23 408 24
rect 413 26 423 27
rect 413 24 415 26
rect 417 24 423 26
rect 413 23 423 24
rect 468 59 492 63
rect 511 59 515 63
rect 557 67 577 68
rect 557 65 573 67
rect 575 65 577 67
rect 557 64 577 65
rect 589 66 595 73
rect 589 64 591 66
rect 593 64 595 66
rect 466 55 472 59
rect 488 58 528 59
rect 488 56 512 58
rect 514 56 528 58
rect 466 45 470 55
rect 476 54 480 56
rect 488 55 528 56
rect 476 52 477 54
rect 479 52 480 54
rect 476 51 480 52
rect 466 43 467 45
rect 469 43 470 45
rect 466 41 470 43
rect 473 47 480 51
rect 473 36 477 47
rect 516 42 520 47
rect 516 40 517 42
rect 519 40 520 42
rect 459 35 477 36
rect 459 33 461 35
rect 463 34 477 35
rect 463 33 488 34
rect 459 32 484 33
rect 473 31 484 32
rect 486 31 488 33
rect 473 30 488 31
rect 493 33 497 35
rect 493 31 494 33
rect 496 31 497 33
rect 493 26 497 31
rect 516 38 520 40
rect 524 44 528 55
rect 524 42 530 44
rect 524 40 527 42
rect 529 40 530 42
rect 524 38 530 40
rect 524 35 528 38
rect 508 31 528 35
rect 508 27 512 31
rect 472 25 494 26
rect 383 22 408 23
rect 463 22 467 24
rect 472 23 474 25
rect 476 24 494 25
rect 496 24 497 26
rect 476 23 497 24
rect 502 26 512 27
rect 502 24 504 26
rect 506 24 512 26
rect 502 23 512 24
rect 545 56 546 62
rect 557 59 561 64
rect 589 63 595 64
rect 600 66 604 68
rect 600 64 601 66
rect 603 64 604 66
rect 549 55 561 59
rect 549 42 553 55
rect 549 40 550 42
rect 552 40 553 42
rect 549 34 553 40
rect 572 38 573 54
rect 600 59 604 64
rect 609 64 615 73
rect 641 71 643 73
rect 645 71 647 73
rect 641 70 647 71
rect 676 71 678 73
rect 680 71 682 73
rect 609 62 611 64
rect 613 62 615 64
rect 609 61 615 62
rect 676 66 682 71
rect 698 71 700 73
rect 702 71 704 73
rect 676 64 678 66
rect 680 64 682 66
rect 676 63 682 64
rect 689 65 693 67
rect 689 63 690 65
rect 692 63 693 65
rect 698 66 704 71
rect 730 71 732 73
rect 734 71 736 73
rect 730 70 736 71
rect 765 71 767 73
rect 769 71 771 73
rect 698 64 700 66
rect 702 64 704 66
rect 698 63 704 64
rect 765 66 771 71
rect 787 71 789 73
rect 791 71 793 73
rect 765 64 767 66
rect 769 64 771 66
rect 765 63 771 64
rect 778 65 782 67
rect 778 63 779 65
rect 781 63 782 65
rect 787 66 793 71
rect 787 64 789 66
rect 791 64 793 66
rect 787 63 793 64
rect 600 57 601 59
rect 603 58 604 59
rect 603 57 617 58
rect 600 54 617 57
rect 613 42 617 54
rect 613 40 614 42
rect 616 40 617 42
rect 549 30 566 34
rect 613 35 617 40
rect 605 31 617 35
rect 562 28 566 30
rect 472 22 497 23
rect 551 26 557 27
rect 551 24 553 26
rect 555 24 557 26
rect 562 26 563 28
rect 565 26 566 28
rect 562 24 566 26
rect 571 28 577 29
rect 571 26 573 28
rect 575 26 577 28
rect 605 27 609 31
rect 620 28 621 30
rect 374 20 375 22
rect 377 20 378 22
rect 463 20 464 22
rect 466 20 467 22
rect 374 17 378 20
rect 430 19 436 20
rect 430 17 432 19
rect 434 17 436 19
rect 463 17 467 20
rect 519 19 525 20
rect 519 17 521 19
rect 523 17 525 19
rect 551 17 557 24
rect 571 17 577 26
rect 589 26 609 27
rect 589 24 591 26
rect 593 24 609 26
rect 589 23 609 24
rect 646 59 670 63
rect 689 59 693 63
rect 644 55 650 59
rect 666 58 706 59
rect 666 56 690 58
rect 692 56 706 58
rect 644 45 648 55
rect 654 54 658 56
rect 666 55 706 56
rect 654 52 655 54
rect 657 52 658 54
rect 654 51 658 52
rect 644 43 645 45
rect 647 43 648 45
rect 644 41 648 43
rect 651 47 658 51
rect 651 36 655 47
rect 694 42 698 47
rect 694 40 695 42
rect 697 40 698 42
rect 637 35 655 36
rect 637 33 639 35
rect 641 34 655 35
rect 641 33 666 34
rect 637 32 662 33
rect 651 31 662 32
rect 664 31 666 33
rect 651 30 666 31
rect 671 33 675 35
rect 671 31 672 33
rect 674 31 675 33
rect 671 26 675 31
rect 694 38 698 40
rect 702 44 706 55
rect 702 42 708 44
rect 702 40 705 42
rect 707 40 708 42
rect 702 38 708 40
rect 702 35 706 38
rect 686 31 706 35
rect 686 27 690 31
rect 650 25 672 26
rect 641 22 645 24
rect 650 23 652 25
rect 654 24 672 25
rect 674 24 675 26
rect 654 23 675 24
rect 680 26 690 27
rect 680 24 682 26
rect 684 24 690 26
rect 680 23 690 24
rect 735 59 759 63
rect 778 59 782 63
rect 824 67 844 68
rect 824 65 840 67
rect 842 65 844 67
rect 824 64 844 65
rect 733 55 739 59
rect 755 58 795 59
rect 755 56 779 58
rect 781 56 795 58
rect 733 45 737 55
rect 743 54 747 56
rect 755 55 795 56
rect 743 52 744 54
rect 746 52 747 54
rect 743 51 747 52
rect 733 43 734 45
rect 736 43 737 45
rect 733 41 737 43
rect 740 47 747 51
rect 740 36 744 47
rect 783 42 787 47
rect 783 40 784 42
rect 786 40 787 42
rect 726 35 744 36
rect 726 33 728 35
rect 730 34 744 35
rect 730 33 755 34
rect 726 32 751 33
rect 740 31 751 32
rect 753 31 755 33
rect 740 30 755 31
rect 760 33 764 35
rect 760 31 761 33
rect 763 31 764 33
rect 760 26 764 31
rect 783 38 787 40
rect 791 44 795 55
rect 791 42 797 44
rect 791 40 794 42
rect 796 40 797 42
rect 791 38 797 40
rect 791 35 795 38
rect 775 31 795 35
rect 775 27 779 31
rect 739 25 761 26
rect 650 22 675 23
rect 730 22 734 24
rect 739 23 741 25
rect 743 24 761 25
rect 763 24 764 26
rect 743 23 764 24
rect 769 26 779 27
rect 769 24 771 26
rect 773 24 779 26
rect 769 23 779 24
rect 812 56 813 62
rect 824 59 828 64
rect 816 55 828 59
rect 816 42 820 55
rect 816 40 817 42
rect 819 40 820 42
rect 816 34 820 40
rect 839 38 840 54
rect 816 30 833 34
rect 829 28 833 30
rect 739 22 764 23
rect 818 26 824 27
rect 818 24 820 26
rect 822 24 824 26
rect 829 26 830 28
rect 832 26 833 28
rect 829 24 833 26
rect 838 28 844 29
rect 838 26 840 28
rect 842 26 844 28
rect 641 20 642 22
rect 644 20 645 22
rect 730 20 731 22
rect 733 20 734 22
rect 641 17 645 20
rect 697 19 703 20
rect 697 17 699 19
rect 701 17 703 19
rect 730 17 734 20
rect 786 19 792 20
rect 786 17 788 19
rect 790 17 792 19
rect 818 17 824 24
rect 838 17 844 26
<< via1 >>
rect 25 303 27 305
rect 59 303 61 305
rect 318 303 320 305
rect 595 303 597 305
rect 144 290 146 292
rect 22 273 24 275
rect 46 272 48 274
rect 62 264 64 266
rect 14 247 16 249
rect 54 256 56 258
rect 86 260 88 262
rect 144 272 146 274
rect 96 264 98 266
rect 177 272 179 274
rect 128 256 130 258
rect 216 264 218 266
rect 236 264 238 266
rect 266 258 268 260
rect 330 273 332 275
rect 290 257 292 259
rect 306 259 308 261
rect 186 240 188 242
rect 278 240 280 242
rect 354 272 356 274
rect 322 248 324 250
rect 412 272 414 274
rect 364 264 366 266
rect 445 272 447 274
rect 396 256 398 258
rect 484 264 486 266
rect 504 264 506 266
rect 534 258 536 260
rect 598 273 600 275
rect 558 257 560 259
rect 574 259 576 261
rect 454 240 456 242
rect 546 239 548 241
rect 590 256 592 258
rect 622 272 624 274
rect 679 272 681 274
rect 631 264 633 266
rect 712 272 714 274
rect 663 256 665 258
rect 751 264 753 266
rect 771 264 773 266
rect 801 258 803 260
rect 825 257 827 259
rect 841 259 843 261
rect 721 240 723 242
rect 813 240 815 242
rect 14 201 16 203
rect 22 175 24 177
rect 186 208 188 210
rect 278 208 280 210
rect 54 192 56 194
rect 46 176 48 178
rect 62 184 64 186
rect 86 188 88 190
rect 96 184 98 186
rect 128 192 130 194
rect 144 176 146 178
rect 177 176 179 178
rect 216 184 218 186
rect 236 184 238 186
rect 266 190 268 192
rect 290 191 292 193
rect 322 201 324 203
rect 454 208 456 210
rect 546 208 548 210
rect 306 189 308 191
rect 330 175 332 177
rect 354 176 356 178
rect 364 184 366 186
rect 396 192 398 194
rect 412 176 414 178
rect 445 176 447 178
rect 484 184 486 186
rect 504 184 506 186
rect 534 190 536 192
rect 558 191 560 193
rect 590 201 592 203
rect 721 208 723 210
rect 813 208 815 210
rect 574 189 576 191
rect 598 175 600 177
rect 622 176 624 178
rect 631 184 633 186
rect 663 192 665 194
rect 679 176 681 178
rect 712 176 714 178
rect 751 184 753 186
rect 771 184 773 186
rect 801 190 803 192
rect 825 191 827 193
rect 841 189 843 191
rect 22 129 24 131
rect 21 112 23 114
rect 46 128 48 130
rect 62 120 64 122
rect 54 112 56 114
rect 86 116 88 118
rect 144 128 146 130
rect 96 120 98 122
rect 177 128 179 130
rect 128 112 130 114
rect 216 120 218 122
rect 236 120 238 122
rect 266 114 268 116
rect 329 128 331 130
rect 290 113 292 115
rect 306 115 308 117
rect 186 96 188 98
rect 278 96 280 98
rect 354 128 356 130
rect 322 103 324 105
rect 412 128 414 130
rect 364 120 366 122
rect 445 128 447 130
rect 396 112 398 114
rect 484 120 486 122
rect 504 120 506 122
rect 534 114 536 116
rect 598 129 600 131
rect 558 113 560 115
rect 574 115 576 117
rect 454 96 456 98
rect 546 96 548 98
rect 622 128 624 130
rect 590 103 592 105
rect 679 128 681 130
rect 631 120 633 122
rect 712 128 714 130
rect 663 112 665 114
rect 751 120 753 122
rect 771 120 773 122
rect 801 114 803 116
rect 825 113 827 115
rect 841 115 843 117
rect 721 96 723 98
rect 813 96 815 98
rect 14 57 16 59
rect 22 31 24 33
rect 186 64 188 66
rect 278 64 280 66
rect 54 48 56 50
rect 46 32 48 34
rect 62 40 64 42
rect 86 44 88 46
rect 96 40 98 42
rect 128 48 130 50
rect 144 32 146 34
rect 177 32 179 34
rect 216 40 218 42
rect 236 40 238 42
rect 266 46 268 48
rect 290 47 292 49
rect 322 57 324 59
rect 454 64 456 66
rect 546 64 548 66
rect 306 45 308 47
rect 339 40 341 42
rect 354 32 356 34
rect 364 40 366 42
rect 396 48 398 50
rect 412 32 414 34
rect 445 32 447 34
rect 484 40 486 42
rect 504 40 506 42
rect 534 46 536 48
rect 558 47 560 49
rect 590 57 592 59
rect 721 64 723 66
rect 813 64 815 66
rect 574 45 576 47
rect 607 40 609 42
rect 622 32 624 34
rect 631 40 633 42
rect 663 48 665 50
rect 679 32 681 34
rect 712 32 714 34
rect 751 40 753 42
rect 771 40 773 42
rect 801 46 803 48
rect 825 47 827 49
rect 841 45 843 47
rect 308 13 310 15
rect 576 13 578 15
rect 843 13 845 15
rect 12 1 14 3
rect 57 1 59 3
rect 330 1 332 3
rect 595 1 597 3
<< via2 >>
rect 21 303 23 305
rect 63 303 65 305
rect 322 303 324 305
rect 599 303 601 305
rect 12 298 14 300
rect 306 298 308 300
rect 614 298 616 300
rect 50 264 52 266
rect 63 256 65 258
rect 21 183 23 185
rect 15 112 17 114
rect 590 272 592 274
rect 331 264 333 266
rect 322 252 324 254
rect 236 242 238 244
rect 599 256 601 258
rect 504 242 506 244
rect 771 242 773 244
rect 50 192 52 194
rect 312 208 314 210
rect 50 120 52 122
rect 61 112 63 114
rect 331 192 333 194
rect 322 176 324 178
rect 331 120 333 122
rect 580 208 582 210
rect 322 109 324 111
rect 590 193 592 195
rect 598 184 600 186
rect 590 129 592 131
rect 847 208 849 210
rect 599 112 601 114
rect 236 97 238 99
rect 504 97 506 99
rect 771 97 773 99
rect 310 64 312 66
rect 50 48 52 50
rect 17 31 19 33
rect 578 64 580 66
rect 331 48 333 50
rect 590 48 592 50
rect 845 64 847 66
rect 17 1 19 3
rect 61 1 63 3
rect 326 1 328 3
rect 599 1 601 3
<< labels >>
rlabel alu0 127 24 127 24 6 ad1n2
rlabel alu0 138 28 138 28 6 ad1n2
rlabel alu1 141 13 141 13 6 vss
rlabel alu1 141 77 141 77 6 vdd
rlabel alu1 97 39 97 39 1 ad1fa1ha1s
rlabel alu0 118 40 118 40 1 ad1fa1ha1sn
rlabel pmos 161 49 161 49 1 ad1fa1ha1b
rlabel alu1 147 41 147 41 1 ad1fa1ha1a
rlabel via1 178 33 178 33 1 ad1fa1ha1c
rlabel alu0 112 52 112 52 1 ad1fa1ha1cn
rlabel alu1 186 47 186 47 1 ad1fa1ha2s
rlabel alu1 253 25 253 25 1 ad1fa1ha2co
rlabel alu1 236 41 236 41 1 ad1fa1ha2a
rlabel alu1 218 45 218 45 1 ad1fa1ha2b
rlabel alu0 202 56 202 56 1 ad1fa1ha2cn
rlabel polyct0 283 41 283 41 1 ad1fa1ozn
rlabel polyct1 294 41 294 41 1 ad1fa1oa
rlabel polyct1 306 41 306 41 1 ad1fa1ob
rlabel via1 279 65 279 65 1 ad1fa1oz
rlabel alu2 315 77 315 77 1 ad1s0
rlabel nwell 85 48 85 48 3 ad1b0
rlabel alu2 237 66 237 66 1 ad1cin1
rlabel alu2 84 33 84 33 3 ad1a0
rlabel alu0 127 138 127 138 8 ad1n3
rlabel alu0 138 134 138 134 8 ad1n3
rlabel alu1 141 149 141 149 8 vss
rlabel alu1 141 85 141 85 8 vdd
rlabel alu1 97 123 97 123 5 ad1fa2ha2s
rlabel alu0 118 122 118 122 5 ad1fa2ha2sn
rlabel pmos 161 113 161 113 5 ad1fa2ha2b
rlabel alu1 147 121 147 121 5 ad1fa2ha2a
rlabel via1 178 129 178 129 5 ad1fa2ha2c
rlabel alu0 112 110 112 110 5 ad1fa2ha2cn
rlabel alu1 186 115 186 115 5 ad1fa2ha3s
rlabel alu1 253 137 253 137 5 ad1fa2ha3co
rlabel alu1 236 121 236 121 5 ad1fa2ha3a
rlabel alu1 218 117 218 117 5 ad1fa2ha3b
rlabel alu0 202 106 202 106 5 ad1fa2ha3cn
rlabel polyct0 283 121 283 121 5 ad1fa2ozn
rlabel polyct1 294 121 294 121 5 ad1fa2oa
rlabel polyct1 306 121 306 121 5 ad1fa2ob
rlabel via1 279 97 279 97 5 ad1fa2oz
rlabel alu2 315 85 315 85 5 ad1s1
rlabel nwell 85 114 85 114 3 ad1b1
rlabel alu2 237 94 237 94 1 ad1cin2
rlabel alu2 85 129 85 129 3 ad1a1
rlabel alu0 127 168 127 168 6 ad1n4
rlabel alu0 138 172 138 172 6 ad1n4
rlabel alu1 141 157 141 157 6 vss
rlabel alu1 141 221 141 221 6 vdd
rlabel alu1 97 183 97 183 1 ad1fa3ha3s
rlabel alu0 118 184 118 184 1 ad1fa3ha3sn
rlabel pmos 161 193 161 193 1 ad1fa3ha3b
rlabel alu1 147 185 147 185 1 ad1fa3ha3a
rlabel via1 178 177 178 177 1 ad1fa3ha3c
rlabel alu0 112 196 112 196 1 ad1fa3ha3cn
rlabel alu1 186 191 186 191 1 ad1fa3ha4s
rlabel alu1 253 169 253 169 1 ad1fa3ha4co
rlabel alu1 236 185 236 185 1 ad1fa3ha4a
rlabel alu1 218 189 218 189 1 ad1fa3ha4b
rlabel alu0 202 200 202 200 1 ad1fa3ha4cn
rlabel polyct0 283 185 283 185 1 ad1fa3ozn
rlabel polyct1 294 185 294 185 1 ad1fa3oa
rlabel polyct1 306 185 306 185 1 ad1fa3ob
rlabel via1 279 209 279 209 1 ad1fa3oz
rlabel alu2 315 221 315 221 1 ad1s2
rlabel nwell 85 192 85 192 3 ad1b2
rlabel alu2 237 212 237 212 1 ad1cin3
rlabel alu2 86 177 86 177 3 ad1a2
rlabel alu0 127 282 127 282 8 ad1n5
rlabel alu0 138 278 138 278 8 ad1n5
rlabel alu1 141 229 141 229 8 vdd
rlabel alu1 97 267 97 267 5 ad1fa4ha4s
rlabel alu0 118 266 118 266 5 ad1fa4ha4sn
rlabel alu1 147 265 147 265 5 ad1fa4ha4a
rlabel via1 178 273 178 273 5 ad1fa4ha4c
rlabel alu0 112 254 112 254 5 ad1fa4ha4cn
rlabel alu1 186 259 186 259 5 ad1fa4ha5s
rlabel alu1 253 281 253 281 5 ad1fa4ha5co
rlabel alu1 236 265 236 265 5 ad1fa4ha5a
rlabel alu1 218 261 218 261 5 ad1fa4ha5b
rlabel alu0 202 250 202 250 5 ad1fa4ha5cn
rlabel polyct0 283 265 283 265 5 ad1fa4ozn
rlabel polyct1 294 265 294 265 5 ad1fa4oa
rlabel polyct1 306 265 306 265 5 ad1fa4ob
rlabel via1 279 241 279 241 5 ad1fa4oz
rlabel alu2 315 229 315 229 5 ad1s3
rlabel nwell 85 258 85 258 3 ad1b3
rlabel alu2 237 239 237 239 1 ad1cin4
rlabel pmos 161 257 161 257 5 ad1fa4ha4b
rlabel alu1 141 293 141 293 8 vss
rlabel alu2 145 287 145 287 1 ad1a3
rlabel alu1 87 268 87 268 1 a8z
rlabel alu1 47 269 47 269 1 a7z
rlabel alu1 55 253 55 253 1 a8b
rlabel alu1 63 269 63 269 1 a8a
rlabel alu1 15 253 15 253 1 a7b
rlabel alu1 23 269 23 269 1 a7a
rlabel alu1 71 293 71 293 2 vss
rlabel alu2 93 177 93 177 7 X4
rlabel alu1 63 181 63 181 1 a6a
rlabel alu1 55 198 55 198 1 a6b
rlabel alu1 86 183 86 183 1 a6z
rlabel alu1 47 189 47 189 1 a5z
rlabel alu1 23 181 23 181 1 a5a
rlabel alu1 15 197 15 197 1 a5b
rlabel alu1 71 221 71 221 4 vdd
rlabel alu1 71 149 71 149 2 vss
rlabel alu2 94 129 94 129 7 X2
rlabel alu1 22 125 22 125 1 a3b
rlabel alu1 15 109 15 109 1 a3a
rlabel alu1 47 125 47 125 1 a3z
rlabel alu1 63 125 63 125 1 a4b
rlabel alu1 55 109 55 109 1 a4a
rlabel alu1 87 125 87 125 1 a4z
rlabel alu1 71 13 71 13 4 vss
rlabel alu1 71 77 71 77 4 vdd
rlabel alu1 87 39 87 39 1 a2z
rlabel alu1 63 37 63 37 1 a2a
rlabel alu1 55 54 55 54 1 a2b
rlabel alu1 15 53 15 53 1 a1b
rlabel alu1 47 39 47 39 1 a1z
rlabel alu1 23 37 23 37 1 a1a
rlabel alu2 8 58 8 58 3 B0
rlabel alu2 93 33 93 33 7 X0
rlabel alu2 8 130 8 130 3 B0
rlabel alu2 8 202 8 202 3 B0
rlabel alu2 8 273 8 273 3 B0
rlabel alu2 90 49 90 49 1 X1
rlabel alu2 90 112 90 112 1 X3
rlabel alu2 90 194 90 194 1 X5
rlabel alu2 90 256 90 256 1 X7
rlabel alu2 311 77 311 77 1 P1
rlabel alu3 310 67 310 67 1 ad1cout1
rlabel via1 323 104 323 104 1 A1
rlabel via2 323 177 323 177 1 A2
rlabel alu2 313 240 313 240 1 ad1cout4
rlabel alu1 323 248 323 248 1 A3
rlabel alu2 358 33 358 33 1 X8
rlabel alu2 358 177 358 177 1 X10
rlabel alu2 358 273 358 273 1 X11
rlabel alu0 395 24 395 24 6 ad2n2
rlabel alu0 406 28 406 28 6 ad2n2
rlabel alu1 409 13 409 13 6 vss
rlabel alu1 409 77 409 77 6 vdd
rlabel alu1 365 39 365 39 1 ad2fa1ha1s
rlabel alu0 386 40 386 40 1 ad2fa1ha1sn
rlabel pmos 429 49 429 49 1 ad2fa1ha1b
rlabel alu1 415 41 415 41 1 ad2fa1ha1a
rlabel via1 446 33 446 33 1 ad2fa1ha1c
rlabel alu0 380 52 380 52 1 ad2fa1ha1cn
rlabel alu1 454 47 454 47 1 ad2fa1ha2s
rlabel alu1 521 25 521 25 1 ad2fa1ha2co
rlabel alu1 504 41 504 41 1 ad2fa1ha2a
rlabel alu1 486 45 486 45 1 ad2fa1ha2b
rlabel alu0 470 56 470 56 1 ad2fa1ha2cn
rlabel polyct0 551 41 551 41 1 ad2fa1ozn
rlabel polyct1 562 41 562 41 1 ad2fa1oa
rlabel polyct1 574 41 574 41 1 ad2fa1ob
rlabel via1 547 65 547 65 1 ad2fa1oz
rlabel alu2 505 66 505 66 1 ad2cin1
rlabel alu0 395 138 395 138 8 ad2n3
rlabel alu0 406 134 406 134 8 ad2n3
rlabel alu1 409 149 409 149 8 vss
rlabel alu1 409 85 409 85 8 vdd
rlabel alu1 365 123 365 123 5 ad2fa2ha2s
rlabel alu0 386 122 386 122 5 ad2fa2ha2sn
rlabel pmos 429 113 429 113 5 ad2fa2ha2b
rlabel alu1 415 121 415 121 5 ad2fa2ha2a
rlabel via1 446 129 446 129 5 ad2fa2ha2c
rlabel alu0 380 110 380 110 5 ad2fa2ha2cn
rlabel alu1 454 115 454 115 5 ad2fa2ha3s
rlabel alu1 521 137 521 137 5 ad2fa2ha3co
rlabel alu1 504 121 504 121 5 ad2fa2ha3a
rlabel alu1 486 117 486 117 5 ad2fa2ha3b
rlabel alu0 470 106 470 106 5 ad2fa2ha3cn
rlabel polyct0 551 121 551 121 5 ad2fa2ozn
rlabel polyct1 562 121 562 121 5 ad2fa2oa
rlabel polyct1 574 121 574 121 5 ad2fa2ob
rlabel via1 547 97 547 97 5 ad2fa2oz
rlabel alu2 583 85 583 85 5 ad2s1
rlabel alu2 353 114 353 114 3 ad2b1
rlabel alu2 505 94 505 94 1 ad2cin2
rlabel alu0 395 168 395 168 6 ad2n4
rlabel alu0 406 172 406 172 6 ad2n4
rlabel alu1 409 157 409 157 6 vss
rlabel alu1 409 221 409 221 6 vdd
rlabel alu1 365 183 365 183 1 ad2fa3ha3s
rlabel alu0 386 184 386 184 1 ad2fa3ha3sn
rlabel pmos 429 193 429 193 1 ad2fa3ha3b
rlabel alu1 415 185 415 185 1 ad2fa3ha3a
rlabel via1 446 177 446 177 1 ad2fa3ha3c
rlabel alu0 380 196 380 196 1 ad2fa3ha3cn
rlabel alu1 454 191 454 191 1 ad2fa3ha4s
rlabel alu1 521 169 521 169 1 ad2fa3ha4co
rlabel alu1 504 185 504 185 1 ad2fa3ha4a
rlabel alu1 486 189 486 189 1 ad2fa3ha4b
rlabel alu0 470 200 470 200 1 ad2fa3ha4cn
rlabel polyct0 551 185 551 185 1 ad2fa3ozn
rlabel polyct1 562 185 562 185 1 ad2fa3oa
rlabel polyct1 574 185 574 185 1 ad2fa3ob
rlabel via1 547 209 547 209 1 ad2fa3oz
rlabel alu2 583 221 583 221 1 ad2s2
rlabel alu2 353 192 353 192 3 ad2b2
rlabel alu2 505 212 505 212 1 ad2cin3
rlabel alu2 354 177 354 177 3 ad2a2
rlabel alu0 395 282 395 282 8 ad2n5
rlabel alu0 406 278 406 278 8 ad2n5
rlabel alu1 409 229 409 229 8 vdd
rlabel alu1 365 267 365 267 5 ad2fa4ha4s
rlabel alu0 386 266 386 266 5 ad2fa4ha4sn
rlabel alu1 415 265 415 265 5 ad2fa4ha4a
rlabel via1 446 273 446 273 5 ad2fa4ha4c
rlabel alu0 380 254 380 254 5 ad2fa4ha4cn
rlabel alu1 454 259 454 259 5 ad2fa4ha5s
rlabel alu1 521 281 521 281 5 ad2fa4ha5co
rlabel alu1 504 265 504 265 5 ad2fa4ha5a
rlabel alu1 486 261 486 261 5 ad2fa4ha5b
rlabel alu0 470 250 470 250 5 ad2fa4ha5cn
rlabel polyct0 551 265 551 265 5 ad2fa4ozn
rlabel polyct1 562 265 562 265 5 ad2fa4oa
rlabel polyct1 574 265 574 265 5 ad2fa4ob
rlabel alu2 583 229 583 229 5 ad2s3
rlabel alu2 353 258 353 258 3 ad2b3
rlabel alu2 505 239 505 239 1 ad2cin4
rlabel alu2 354 273 354 273 3 ad2a3
rlabel alu2 586 240 586 240 7 ad2cout4
rlabel pmos 429 257 429 257 5 ad2fa4ha4b
rlabel alu1 409 293 409 293 8 vss
rlabel alu2 358 49 358 49 1 ad2b0
rlabel alu2 361 129 361 129 1 X9
rlabel alu1 591 248 591 248 1 A3
rlabel alu2 593 178 593 178 1 A2
rlabel via1 591 104 591 104 1 A1
rlabel alu1 599 32 599 32 1 A0
rlabel via1 623 273 623 273 1 X15
rlabel via1 623 177 623 177 1 X14
rlabel via1 623 129 623 129 1 X13
rlabel via1 623 33 623 33 1 X12
rlabel via2 581 209 581 209 1 ad2cout3
rlabel alu2 582 96 582 96 1 ad2cout2
rlabel via2 579 65 579 65 1 ad2cout1
rlabel alu2 644 177 644 177 3 ad3a2
rlabel alu2 580 77 580 77 1 P2
rlabel via1 547 240 547 240 5 ad2fa4oz
rlabel alu1 676 293 676 293 8 vss
rlabel pmos 696 257 696 257 5 ad3fa4ha4b
rlabel alu2 772 239 772 239 1 ad3cin4
rlabel via1 814 241 814 241 5 ad3fa4oz
rlabel polyct1 841 265 841 265 5 ad3fa4ob
rlabel polyct1 829 265 829 265 5 ad3fa4oa
rlabel polyct0 818 265 818 265 5 ad3fa4ozn
rlabel alu0 737 250 737 250 5 ad3fa4ha5cn
rlabel alu1 753 261 753 261 5 ad3fa4ha5b
rlabel alu1 771 265 771 265 5 ad3fa4ha5a
rlabel alu1 788 281 788 281 5 ad3fa4ha5co
rlabel alu1 721 259 721 259 5 ad3fa4ha5s
rlabel alu0 647 254 647 254 5 ad3fa4ha4cn
rlabel via1 713 273 713 273 5 ad3fa4ha4c
rlabel alu1 682 265 682 265 5 ad3fa4ha4a
rlabel alu0 653 266 653 266 5 ad3fa4ha4sn
rlabel alu1 632 267 632 267 5 ad3fa4ha4s
rlabel alu1 676 229 676 229 8 vdd
rlabel alu0 673 278 673 278 8 ad3n5
rlabel alu0 662 282 662 282 8 ad3n5
rlabel alu2 772 212 772 212 1 ad3cin3
rlabel alu2 853 210 853 210 7 ad3cout3
rlabel via1 814 209 814 209 1 ad3fa3oz
rlabel polyct1 841 185 841 185 1 ad3fa3ob
rlabel polyct1 829 185 829 185 1 ad3fa3oa
rlabel polyct0 818 185 818 185 1 ad3fa3ozn
rlabel alu0 737 200 737 200 1 ad3fa3ha4cn
rlabel alu1 753 189 753 189 1 ad3fa3ha4b
rlabel alu1 771 185 771 185 1 ad3fa3ha4a
rlabel alu1 788 169 788 169 1 ad3fa3ha4co
rlabel alu1 721 191 721 191 1 ad3fa3ha4s
rlabel alu0 647 196 647 196 1 ad3fa3ha3cn
rlabel via1 713 177 713 177 1 ad3fa3ha3c
rlabel alu1 682 185 682 185 1 ad3fa3ha3a
rlabel pmos 696 193 696 193 1 ad3fa3ha3b
rlabel alu0 653 184 653 184 1 ad3fa3ha3sn
rlabel alu1 632 183 632 183 1 ad3fa3ha3s
rlabel alu1 676 221 676 221 6 vdd
rlabel alu1 676 157 676 157 6 vss
rlabel alu0 673 172 673 172 6 ad3n4
rlabel alu0 662 168 662 168 6 ad3n4
rlabel alu2 772 94 772 94 1 ad3cin2
rlabel via1 814 97 814 97 5 ad3fa2oz
rlabel polyct1 841 121 841 121 5 ad3fa2ob
rlabel polyct1 829 121 829 121 5 ad3fa2oa
rlabel polyct0 818 121 818 121 5 ad3fa2ozn
rlabel alu0 737 106 737 106 5 ad3fa2ha3cn
rlabel alu1 753 117 753 117 5 ad3fa2ha3b
rlabel alu1 771 121 771 121 5 ad3fa2ha3a
rlabel alu1 788 137 788 137 5 ad3fa2ha3co
rlabel alu1 721 115 721 115 5 ad3fa2ha3s
rlabel alu0 647 110 647 110 5 ad3fa2ha2cn
rlabel via1 713 129 713 129 5 ad3fa2ha2c
rlabel alu1 682 121 682 121 5 ad3fa2ha2a
rlabel pmos 696 113 696 113 5 ad3fa2ha2b
rlabel alu0 653 122 653 122 5 ad3fa2ha2sn
rlabel alu1 632 123 632 123 5 ad3fa2ha2s
rlabel alu1 676 85 676 85 8 vdd
rlabel alu1 676 149 676 149 8 vss
rlabel alu0 673 134 673 134 8 ad3n3
rlabel alu0 662 138 662 138 8 ad3n3
rlabel alu2 772 66 772 66 1 ad3cin1
rlabel alu2 853 66 853 66 7 ad3cout1
rlabel via1 814 65 814 65 1 ad3fa1oz
rlabel polyct1 841 41 841 41 1 ad3fa1ob
rlabel polyct1 829 41 829 41 1 ad3fa1oa
rlabel polyct0 818 41 818 41 1 ad3fa1ozn
rlabel alu0 737 56 737 56 1 ad3fa1ha2cn
rlabel alu1 753 45 753 45 1 ad3fa1ha2b
rlabel alu1 771 41 771 41 1 ad3fa1ha2a
rlabel alu1 788 25 788 25 1 ad3fa1ha2co
rlabel alu1 721 47 721 47 1 ad3fa1ha2s
rlabel alu0 647 52 647 52 1 ad3fa1ha1cn
rlabel via1 713 33 713 33 1 ad3fa1ha1c
rlabel alu1 682 41 682 41 1 ad3fa1ha1a
rlabel pmos 696 49 696 49 1 ad3fa1ha1b
rlabel alu0 653 40 653 40 1 ad3fa1ha1sn
rlabel alu1 632 39 632 39 1 ad3fa1ha1s
rlabel alu1 676 77 676 77 6 vdd
rlabel alu1 676 13 676 13 6 vss
rlabel alu0 673 28 673 28 6 ad3n2
rlabel alu0 662 24 662 24 6 ad3n2
rlabel alu2 839 77 839 77 1 P3
rlabel alu2 834 85 834 85 1 P4
rlabel alu2 834 220 834 220 1 P5
rlabel alu2 833 230 833 230 1 P6
rlabel alu2 848 96 848 96 1 ad3cout2
rlabel alu3 51 287 51 287 1 B1
rlabel alu2 315 96 315 96 1 ad1cout2
rlabel via2 313 209 313 209 1 ad1cout3
rlabel alu3 332 286 332 286 1 B2
rlabel alu3 591 287 591 287 1 B3
rlabel alu2 87 286 87 286 1 P0
rlabel alu2 5 6 5 6 3 A0
rlabel alu1 5 2 5 2 2 A1
rlabel alu2 14 299 14 299 1 A2
rlabel alu1 14 304 14 304 5 A3
rlabel via1 340 41 340 41 1 A0
rlabel via1 15 248 15 248 1 A0
rlabel via1 55 257 55 257 1 A3
rlabel alu2 852 240 852 240 7 P7
<< end >>
