magic
tech scmos
timestamp 1199973072
<< ab >>
rect 0 0 32 88
<< nwell >>
rect -5 40 37 97
<< pwell >>
rect -5 -9 37 40
<< poly >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 41 14 43
rect 2 39 7 41
rect 9 39 14 41
rect 2 37 14 39
rect 18 41 30 43
rect 18 39 23 41
rect 25 39 30 41
rect 18 37 30 39
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndif >>
rect 2 25 9 34
rect 2 23 4 25
rect 6 23 9 25
rect 2 18 9 23
rect 2 16 4 18
rect 6 16 9 18
rect 2 14 9 16
rect 11 32 21 34
rect 11 30 15 32
rect 17 30 21 32
rect 11 25 21 30
rect 11 23 15 25
rect 17 23 21 25
rect 11 14 21 23
rect 23 18 30 34
rect 23 16 26 18
rect 28 16 30 18
rect 23 14 30 16
rect 13 2 19 14
<< pdif >>
rect 13 74 19 86
rect 2 72 9 74
rect 2 70 4 72
rect 6 70 9 72
rect 2 65 9 70
rect 2 63 4 65
rect 6 63 9 65
rect 2 46 9 63
rect 11 46 21 74
rect 23 62 30 74
rect 23 60 26 62
rect 28 60 30 62
rect 23 55 30 60
rect 23 53 26 55
rect 28 53 30 55
rect 23 46 30 53
<< alu1 >>
rect -2 89 34 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 34 89
rect -2 86 34 87
rect 3 81 7 86
rect 3 79 4 81
rect 6 79 7 81
rect 3 72 7 79
rect 3 70 4 72
rect 6 70 7 72
rect 3 65 7 70
rect 3 63 4 65
rect 6 63 7 65
rect 3 61 7 63
rect 22 62 29 64
rect 22 60 26 62
rect 28 60 29 62
rect 22 55 29 60
rect 6 41 10 55
rect 6 39 7 41
rect 9 39 10 41
rect 6 33 10 39
rect 14 53 26 55
rect 28 53 29 55
rect 14 51 29 53
rect 14 32 18 51
rect 14 30 15 32
rect 17 30 18 32
rect 3 25 7 27
rect 3 23 4 25
rect 6 23 7 25
rect 3 18 7 23
rect 3 16 4 18
rect 6 16 7 18
rect 14 25 18 30
rect 22 41 26 47
rect 22 39 23 41
rect 25 39 26 41
rect 22 25 26 39
rect 14 23 15 25
rect 17 23 18 25
rect 14 17 18 23
rect 25 18 29 20
rect 3 9 7 16
rect 3 7 4 9
rect 6 7 7 9
rect 3 2 7 7
rect 25 16 26 18
rect 28 16 29 18
rect 25 9 29 16
rect 25 7 26 9
rect 28 7 29 9
rect 25 2 29 7
rect -2 1 34 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< alu2 >>
rect -2 89 34 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 34 89
rect -2 81 34 87
rect -2 79 4 81
rect 6 79 34 81
rect -2 76 34 79
rect -2 9 34 12
rect -2 7 4 9
rect 6 7 26 9
rect 28 7 34 9
rect -2 1 34 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 32 3
rect 25 -1 27 1
rect 29 -1 32 1
rect 25 -3 32 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 32 91
rect 25 87 27 89
rect 29 87 32 89
rect 25 85 32 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
<< polyct1 >>
rect 7 39 9 41
rect 23 39 25 41
<< ndifct1 >>
rect 4 23 6 25
rect 4 16 6 18
rect 15 30 17 32
rect 15 23 17 25
rect 26 16 28 18
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
<< pdifct1 >>
rect 4 70 6 72
rect 4 63 6 65
rect 26 60 28 62
rect 26 53 28 55
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 4 79 6 81
rect 4 7 6 9
rect 26 7 28 9
rect 7 -1 9 1
rect 23 -1 25 1
<< labels >>
rlabel alu1 8 44 8 44 6 a
rlabel alu1 16 36 16 36 6 z
rlabel alu1 24 36 24 36 6 b
rlabel alu1 24 60 24 60 6 z
rlabel alu2 16 6 16 6 6 vss
rlabel alu2 16 82 16 82 6 vdd
<< end >>
