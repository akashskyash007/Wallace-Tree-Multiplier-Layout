magic
tech scmos
timestamp 1199203601
<< ab >>
rect 0 0 160 80
<< nwell >>
rect -5 36 165 88
<< pwell >>
rect -5 -8 165 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 71 72
rect 49 67 51 70
rect 59 67 61 70
rect 69 67 71 70
rect 79 67 81 72
rect 89 67 91 72
rect 119 67 121 72
rect 129 67 131 72
rect 139 67 141 72
rect 149 67 151 72
rect 99 61 101 65
rect 109 61 111 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 41 39
rect 49 38 51 42
rect 59 38 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 99 39 101 42
rect 109 39 111 42
rect 119 39 121 42
rect 129 39 131 42
rect 139 39 141 42
rect 149 39 151 42
rect 66 37 72 39
rect 9 35 11 37
rect 13 35 32 37
rect 9 33 32 35
rect 66 35 68 37
rect 70 35 72 37
rect 20 30 22 33
rect 30 30 32 33
rect 50 30 52 34
rect 60 30 62 34
rect 66 33 72 35
rect 70 30 72 33
rect 77 37 94 39
rect 77 35 79 37
rect 81 35 86 37
rect 88 35 94 37
rect 77 33 94 35
rect 77 30 79 33
rect 92 30 94 33
rect 99 37 111 39
rect 99 35 101 37
rect 103 35 111 37
rect 99 33 111 35
rect 115 37 121 39
rect 115 35 117 37
rect 119 35 121 37
rect 115 33 121 35
rect 128 37 151 39
rect 128 35 147 37
rect 149 35 151 37
rect 128 33 151 35
rect 99 30 101 33
rect 109 30 111 33
rect 116 30 118 33
rect 128 30 130 33
rect 138 30 140 33
rect 20 6 22 11
rect 30 8 32 11
rect 50 8 52 11
rect 60 8 62 11
rect 30 6 62 8
rect 70 6 72 10
rect 77 6 79 10
rect 92 8 94 16
rect 99 12 101 16
rect 109 12 111 16
rect 116 8 118 16
rect 92 6 118 8
rect 128 6 130 11
rect 138 6 140 11
<< ndif >>
rect 13 23 20 30
rect 13 21 15 23
rect 17 21 20 23
rect 13 15 20 21
rect 13 13 15 15
rect 17 13 20 15
rect 13 11 20 13
rect 22 28 30 30
rect 22 26 25 28
rect 27 26 30 28
rect 22 21 30 26
rect 22 19 25 21
rect 27 19 30 21
rect 22 11 30 19
rect 32 23 39 30
rect 45 23 50 30
rect 32 21 35 23
rect 37 21 39 23
rect 32 15 39 21
rect 43 21 50 23
rect 43 19 45 21
rect 47 19 50 21
rect 43 17 50 19
rect 32 13 35 15
rect 37 13 39 15
rect 32 11 39 13
rect 45 11 50 17
rect 52 28 60 30
rect 52 26 55 28
rect 57 26 60 28
rect 52 11 60 26
rect 62 21 70 30
rect 62 19 65 21
rect 67 19 70 21
rect 62 11 70 19
rect 65 10 70 11
rect 72 10 77 30
rect 79 16 92 30
rect 94 16 99 30
rect 101 21 109 30
rect 101 19 104 21
rect 106 19 109 21
rect 101 16 109 19
rect 111 16 116 30
rect 118 20 128 30
rect 118 18 121 20
rect 123 18 128 20
rect 118 16 128 18
rect 79 11 90 16
rect 79 10 84 11
rect 81 9 84 10
rect 86 9 90 11
rect 81 7 90 9
rect 120 11 128 16
rect 130 28 138 30
rect 130 26 133 28
rect 135 26 138 28
rect 130 21 138 26
rect 130 19 133 21
rect 135 19 138 21
rect 130 11 138 19
rect 140 23 147 30
rect 140 21 143 23
rect 145 21 147 23
rect 140 15 147 21
rect 140 13 143 15
rect 145 13 147 15
rect 140 11 147 13
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 42 19 59
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 42 39 59
rect 41 67 46 70
rect 41 60 49 67
rect 41 58 44 60
rect 46 58 49 60
rect 41 53 49 58
rect 41 51 44 53
rect 46 51 49 53
rect 41 42 49 51
rect 51 62 59 67
rect 51 60 54 62
rect 56 60 59 62
rect 51 46 59 60
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 53 69 67
rect 61 51 64 53
rect 66 51 69 53
rect 61 46 69 51
rect 61 44 64 46
rect 66 44 69 46
rect 61 42 69 44
rect 71 62 79 67
rect 71 60 74 62
rect 76 60 79 62
rect 71 55 79 60
rect 71 53 74 55
rect 76 53 79 55
rect 71 42 79 53
rect 81 53 89 67
rect 81 51 84 53
rect 86 51 89 53
rect 81 46 89 51
rect 81 44 84 46
rect 86 44 89 46
rect 81 42 89 44
rect 91 61 96 67
rect 114 61 119 67
rect 91 55 99 61
rect 91 53 94 55
rect 96 53 99 55
rect 91 42 99 53
rect 101 46 109 61
rect 101 44 104 46
rect 106 44 109 46
rect 101 42 109 44
rect 111 54 119 61
rect 111 52 114 54
rect 116 52 119 54
rect 111 42 119 52
rect 121 53 129 67
rect 121 51 124 53
rect 126 51 129 53
rect 121 46 129 51
rect 121 44 124 46
rect 126 44 129 46
rect 121 42 129 44
rect 131 65 139 67
rect 131 63 134 65
rect 136 63 139 65
rect 131 57 139 63
rect 131 55 134 57
rect 136 55 139 57
rect 131 42 139 55
rect 141 53 149 67
rect 141 51 144 53
rect 146 51 149 53
rect 141 46 149 51
rect 141 44 144 46
rect 146 44 149 46
rect 141 42 149 44
rect 151 65 158 67
rect 151 63 154 65
rect 156 63 158 65
rect 151 57 158 63
rect 151 55 154 57
rect 156 55 158 57
rect 151 42 158 55
<< alu1 >>
rect -2 81 162 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 162 81
rect -2 68 162 79
rect 52 46 58 47
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 2 25 6 33
rect 42 44 54 46
rect 56 44 58 46
rect 42 42 58 44
rect 42 22 46 42
rect 154 38 158 47
rect 145 37 158 38
rect 145 35 147 37
rect 149 35 158 37
rect 145 33 158 35
rect 42 21 108 22
rect 42 19 45 21
rect 47 19 65 21
rect 67 19 104 21
rect 106 19 108 21
rect 42 18 108 19
rect -2 11 162 12
rect -2 9 84 11
rect 86 9 162 11
rect -2 1 162 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 162 1
rect -2 -2 162 -1
<< ptie >>
rect 0 1 160 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 160 1
rect 0 -3 160 -1
<< ntie >>
rect 0 81 160 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 160 81
rect 0 77 160 79
<< nmos >>
rect 20 11 22 30
rect 30 11 32 30
rect 50 11 52 30
rect 60 11 62 30
rect 70 10 72 30
rect 77 10 79 30
rect 92 16 94 30
rect 99 16 101 30
rect 109 16 111 30
rect 116 16 118 30
rect 128 11 130 30
rect 138 11 140 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 67
rect 59 42 61 67
rect 69 42 71 67
rect 79 42 81 67
rect 89 42 91 67
rect 99 42 101 61
rect 109 42 111 61
rect 119 42 121 67
rect 129 42 131 67
rect 139 42 141 67
rect 149 42 151 67
<< polyct0 >>
rect 68 35 70 37
rect 79 35 81 37
rect 86 35 88 37
rect 101 35 103 37
rect 117 35 119 37
<< polyct1 >>
rect 11 35 13 37
rect 147 35 149 37
<< ndifct0 >>
rect 15 21 17 23
rect 15 13 17 15
rect 25 26 27 28
rect 25 19 27 21
rect 35 21 37 23
rect 35 13 37 15
rect 55 26 57 28
rect 121 18 123 20
rect 133 26 135 28
rect 133 19 135 21
rect 143 21 145 23
rect 143 13 145 15
<< ndifct1 >>
rect 45 19 47 21
rect 65 19 67 21
rect 104 19 106 21
rect 84 9 86 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
<< pdifct0 >>
rect 4 51 6 53
rect 4 44 6 46
rect 14 66 16 68
rect 14 59 16 61
rect 24 51 26 53
rect 24 44 26 46
rect 34 66 36 68
rect 34 59 36 61
rect 44 58 46 60
rect 44 51 46 53
rect 54 60 56 62
rect 64 51 66 53
rect 64 44 66 46
rect 74 60 76 62
rect 74 53 76 55
rect 84 51 86 53
rect 84 44 86 46
rect 94 53 96 55
rect 104 44 106 46
rect 114 52 116 54
rect 124 51 126 53
rect 124 44 126 46
rect 134 63 136 65
rect 134 55 136 57
rect 144 51 146 53
rect 144 44 146 46
rect 154 63 156 65
rect 154 55 156 57
<< pdifct1 >>
rect 54 44 56 46
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 61 18 66
rect 12 59 14 61
rect 16 59 18 61
rect 12 58 18 59
rect 32 66 34 68
rect 36 66 38 68
rect 32 61 38 66
rect 133 65 137 68
rect 133 63 134 65
rect 136 63 137 65
rect 52 62 97 63
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 43 60 47 62
rect 43 58 44 60
rect 46 58 47 60
rect 52 60 54 62
rect 56 60 74 62
rect 76 60 97 62
rect 52 59 97 60
rect 43 54 47 58
rect 73 55 77 59
rect 93 55 97 59
rect 133 57 137 63
rect 133 55 134 57
rect 136 55 137 57
rect 153 65 157 68
rect 153 63 154 65
rect 156 63 157 65
rect 153 57 157 63
rect 153 55 154 57
rect 156 55 157 57
rect 2 53 68 54
rect 2 51 4 53
rect 6 51 24 53
rect 26 51 44 53
rect 46 51 64 53
rect 66 51 68 53
rect 73 53 74 55
rect 76 53 77 55
rect 73 51 77 53
rect 82 53 87 55
rect 82 51 84 53
rect 86 51 87 53
rect 93 53 94 55
rect 96 54 118 55
rect 96 53 114 54
rect 93 52 114 53
rect 116 52 118 54
rect 93 51 118 52
rect 123 53 127 55
rect 133 53 137 55
rect 143 53 147 55
rect 153 53 157 55
rect 123 51 124 53
rect 126 51 127 53
rect 2 50 68 51
rect 2 46 7 50
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 23 46 28 50
rect 62 47 68 50
rect 82 47 87 51
rect 23 44 24 46
rect 26 44 28 46
rect 23 42 28 44
rect 24 28 28 42
rect 24 26 25 28
rect 27 26 28 28
rect 14 23 18 25
rect 14 21 15 23
rect 17 21 18 23
rect 14 15 18 21
rect 24 21 28 26
rect 62 46 78 47
rect 62 44 64 46
rect 66 44 78 46
rect 62 43 78 44
rect 82 46 98 47
rect 82 44 84 46
rect 86 44 98 46
rect 82 43 98 44
rect 102 46 117 47
rect 102 44 104 46
rect 106 44 117 46
rect 102 43 117 44
rect 24 19 25 21
rect 27 19 28 21
rect 24 17 28 19
rect 34 23 38 25
rect 34 21 35 23
rect 37 21 38 23
rect 14 13 15 15
rect 17 13 18 15
rect 14 12 18 13
rect 34 15 38 21
rect 67 37 71 39
rect 67 35 68 37
rect 70 35 71 37
rect 67 30 71 35
rect 74 38 78 43
rect 94 38 98 43
rect 113 38 117 43
rect 123 46 127 51
rect 143 51 144 53
rect 146 51 147 53
rect 143 46 147 51
rect 123 44 124 46
rect 126 44 144 46
rect 146 44 147 46
rect 123 42 147 44
rect 74 37 90 38
rect 74 35 79 37
rect 81 35 86 37
rect 88 35 90 37
rect 74 34 90 35
rect 94 37 105 38
rect 94 35 101 37
rect 103 35 105 37
rect 94 34 105 35
rect 113 37 121 38
rect 113 35 117 37
rect 119 35 121 37
rect 113 34 121 35
rect 94 30 98 34
rect 132 30 136 42
rect 53 28 136 30
rect 53 26 55 28
rect 57 26 133 28
rect 135 26 136 28
rect 53 25 59 26
rect 120 20 124 22
rect 120 18 121 20
rect 123 18 124 20
rect 34 13 35 15
rect 37 13 38 15
rect 34 12 38 13
rect 120 12 124 18
rect 132 21 136 26
rect 132 19 133 21
rect 135 19 136 21
rect 132 17 136 19
rect 142 23 146 25
rect 142 21 143 23
rect 145 21 146 23
rect 142 15 146 21
rect 142 13 143 15
rect 145 13 146 15
rect 142 12 146 13
<< labels >>
rlabel alu0 4 48 4 48 6 bn
rlabel alu0 26 35 26 35 6 bn
rlabel alu0 45 56 45 56 6 bn
rlabel alu0 69 32 69 32 6 an
rlabel alu0 70 45 70 45 6 bn
rlabel alu0 82 36 82 36 6 bn
rlabel alu0 84 49 84 49 6 an
rlabel alu0 35 52 35 52 6 bn
rlabel alu0 90 45 90 45 6 an
rlabel alu0 99 36 99 36 6 an
rlabel alu0 115 40 115 40 6 bn
rlabel alu0 109 45 109 45 6 bn
rlabel alu0 94 28 94 28 6 an
rlabel alu0 134 31 134 31 6 an
rlabel alu0 145 48 145 48 6 an
rlabel alu0 125 48 125 48 6 an
rlabel alu1 4 32 4 32 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 76 20 76 20 6 z
rlabel alu1 44 32 44 32 6 z
rlabel alu1 52 44 52 44 6 z
rlabel alu1 80 6 80 6 6 vss
rlabel alu1 100 20 100 20 6 z
rlabel alu1 92 20 92 20 6 z
rlabel alu1 84 20 84 20 6 z
rlabel alu1 80 74 80 74 6 vdd
rlabel polyct1 148 36 148 36 6 a
rlabel alu1 156 40 156 40 6 a
<< end >>
