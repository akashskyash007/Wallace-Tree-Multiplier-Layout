magic
tech scmos
timestamp 1199203158
<< ab >>
rect 0 0 96 72
<< nwell >>
rect -5 32 101 77
<< pwell >>
rect -5 -5 101 32
<< poly >>
rect 12 66 14 70
rect 19 66 21 70
rect 29 66 31 70
rect 36 66 38 70
rect 52 66 54 70
rect 59 66 61 70
rect 69 66 71 70
rect 76 66 78 70
rect 12 35 14 38
rect 19 35 21 38
rect 29 35 31 38
rect 36 35 38 38
rect 52 35 54 38
rect 59 35 61 38
rect 69 35 71 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 31 35
rect 19 31 24 33
rect 26 31 31 33
rect 19 29 31 31
rect 35 33 41 35
rect 35 31 37 33
rect 39 31 41 33
rect 35 29 41 31
rect 9 26 11 29
rect 19 26 21 29
rect 29 26 31 29
rect 39 26 41 29
rect 49 33 55 35
rect 49 31 51 33
rect 53 31 55 33
rect 49 29 55 31
rect 59 33 71 35
rect 76 35 78 38
rect 76 33 87 35
rect 59 31 67 33
rect 69 31 71 33
rect 59 29 71 31
rect 49 26 51 29
rect 59 26 61 29
rect 69 26 71 29
rect 81 31 83 33
rect 85 31 87 33
rect 81 29 87 31
rect 81 26 83 29
rect 69 12 71 17
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 39 7 41 12
rect 49 7 51 12
rect 59 7 61 12
rect 81 12 83 17
<< ndif >>
rect 4 18 9 26
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 12 19 22
rect 21 16 29 26
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 31 24 39 26
rect 31 22 34 24
rect 36 22 39 24
rect 31 12 39 22
rect 41 23 49 26
rect 41 21 44 23
rect 46 21 49 23
rect 41 16 49 21
rect 41 14 44 16
rect 46 14 49 16
rect 41 12 49 14
rect 51 16 59 26
rect 51 14 54 16
rect 56 14 59 16
rect 51 12 59 14
rect 61 24 69 26
rect 61 22 64 24
rect 66 22 69 24
rect 61 17 69 22
rect 71 17 81 26
rect 83 23 88 26
rect 83 21 90 23
rect 83 19 86 21
rect 88 19 90 21
rect 83 17 90 19
rect 61 12 66 17
rect 73 7 79 17
rect 73 5 75 7
rect 77 5 79 7
rect 73 3 79 5
<< pdif >>
rect 4 64 12 66
rect 4 62 7 64
rect 9 62 12 64
rect 4 57 12 62
rect 4 55 7 57
rect 9 55 12 57
rect 4 38 12 55
rect 14 38 19 66
rect 21 57 29 66
rect 21 55 24 57
rect 26 55 29 57
rect 21 50 29 55
rect 21 48 24 50
rect 26 48 29 50
rect 21 38 29 48
rect 31 38 36 66
rect 38 64 52 66
rect 38 62 45 64
rect 47 62 52 64
rect 38 57 52 62
rect 38 55 45 57
rect 47 55 52 57
rect 38 38 52 55
rect 54 38 59 66
rect 61 57 69 66
rect 61 55 64 57
rect 66 55 69 57
rect 61 50 69 55
rect 61 48 64 50
rect 66 48 69 50
rect 61 38 69 48
rect 71 38 76 66
rect 78 59 83 66
rect 78 57 88 59
rect 78 55 83 57
rect 85 55 88 57
rect 78 50 88 55
rect 78 48 83 50
rect 85 48 88 50
rect 78 38 88 48
<< alu1 >>
rect -2 67 98 72
rect -2 65 89 67
rect 91 65 98 67
rect -2 64 98 65
rect 63 57 70 59
rect 63 55 64 57
rect 66 55 70 57
rect 63 53 70 55
rect 63 50 67 53
rect 2 48 24 50
rect 26 48 64 50
rect 66 48 67 50
rect 2 46 67 48
rect 2 25 6 46
rect 74 42 78 51
rect 12 38 40 42
rect 36 35 40 38
rect 50 38 86 42
rect 17 33 31 34
rect 17 31 24 33
rect 26 31 31 33
rect 17 30 31 31
rect 36 33 46 35
rect 36 31 37 33
rect 39 31 46 33
rect 36 29 46 31
rect 50 33 54 38
rect 50 31 51 33
rect 53 31 54 33
rect 50 29 54 31
rect 65 33 78 34
rect 65 31 67 33
rect 69 31 78 33
rect 65 30 78 31
rect 2 24 38 25
rect 2 22 14 24
rect 16 22 34 24
rect 36 22 38 24
rect 2 21 38 22
rect 74 21 78 30
rect 82 33 86 38
rect 82 31 83 33
rect 85 31 86 33
rect 82 29 86 31
rect -2 7 98 8
rect -2 5 75 7
rect 77 5 85 7
rect 87 5 98 7
rect -2 0 98 5
<< ptie >>
rect 83 7 89 9
rect 83 5 85 7
rect 87 5 89 7
rect 83 3 89 5
<< ntie >>
rect 87 67 93 69
rect 87 65 89 67
rect 91 65 93 67
rect 87 63 93 65
<< nmos >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 12 31 26
rect 39 12 41 26
rect 49 12 51 26
rect 59 12 61 26
rect 69 17 71 26
rect 81 17 83 26
<< pmos >>
rect 12 38 14 66
rect 19 38 21 66
rect 29 38 31 66
rect 36 38 38 66
rect 52 38 54 66
rect 59 38 61 66
rect 69 38 71 66
rect 76 38 78 66
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 24 31 26 33
rect 37 31 39 33
rect 51 31 53 33
rect 67 31 69 33
rect 83 31 85 33
<< ndifct0 >>
rect 4 14 6 16
rect 24 14 26 16
rect 44 21 46 23
rect 44 14 46 16
rect 54 14 56 16
rect 64 22 66 24
rect 86 19 88 21
<< ndifct1 >>
rect 14 22 16 24
rect 34 22 36 24
rect 75 5 77 7
<< ntiect1 >>
rect 89 65 91 67
<< ptiect1 >>
rect 85 5 87 7
<< pdifct0 >>
rect 7 62 9 64
rect 7 55 9 57
rect 24 55 26 57
rect 45 62 47 64
rect 45 55 47 57
rect 83 55 85 57
rect 83 48 85 50
<< pdifct1 >>
rect 24 48 26 50
rect 64 55 66 57
rect 64 48 66 50
<< alu0 >>
rect 5 62 7 64
rect 9 62 11 64
rect 5 57 11 62
rect 43 62 45 64
rect 47 62 49 64
rect 5 55 7 57
rect 9 55 11 57
rect 5 54 11 55
rect 23 57 27 59
rect 23 55 24 57
rect 26 55 27 57
rect 23 50 27 55
rect 43 57 49 62
rect 43 55 45 57
rect 47 55 49 57
rect 43 54 49 55
rect 82 57 86 64
rect 82 55 83 57
rect 85 55 86 57
rect 82 50 86 55
rect 82 48 83 50
rect 85 48 86 50
rect 82 46 86 48
rect 10 38 12 42
rect 10 33 14 38
rect 10 31 11 33
rect 13 31 14 33
rect 10 29 14 31
rect 43 24 68 25
rect 43 23 64 24
rect 43 21 44 23
rect 46 22 64 23
rect 66 22 68 24
rect 46 21 68 22
rect 85 21 89 23
rect 43 17 48 21
rect 64 17 68 21
rect 85 19 86 21
rect 88 19 89 21
rect 85 17 89 19
rect 2 16 48 17
rect 2 14 4 16
rect 6 14 24 16
rect 26 14 44 16
rect 46 14 48 16
rect 2 13 48 14
rect 52 16 58 17
rect 52 14 54 16
rect 56 14 58 16
rect 52 8 58 14
rect 64 13 89 17
<< labels >>
rlabel ndifct0 25 15 25 15 6 n3
rlabel alu0 45 19 45 19 6 n3
rlabel alu0 55 23 55 23 6 n3
rlabel alu0 87 18 87 18 6 n3
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 32 28 32 6 b2
rlabel alu1 20 32 20 32 6 b2
rlabel alu1 20 40 20 40 6 b1
rlabel alu1 28 40 28 40 6 b1
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 48 4 48 4 6 vss
rlabel alu1 44 32 44 32 6 b1
rlabel polyct1 52 32 52 32 6 a1
rlabel alu1 36 40 36 40 6 b1
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 48 68 48 68 6 vdd
rlabel alu1 76 24 76 24 6 a2
rlabel polyct1 68 32 68 32 6 a2
rlabel alu1 60 40 60 40 6 a1
rlabel alu1 68 40 68 40 6 a1
rlabel alu1 76 44 76 44 6 a1
rlabel alu1 60 48 60 48 6 z
rlabel alu1 68 56 68 56 6 z
rlabel polyct1 84 32 84 32 6 a1
<< end >>
