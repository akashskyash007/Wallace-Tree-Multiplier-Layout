magic
tech scmos
timestamp 1199202857
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 31 70 33 74
rect 41 70 43 74
rect 53 70 55 74
rect 63 70 65 74
rect 75 70 77 74
rect 85 70 87 74
rect 9 39 11 52
rect 19 49 21 52
rect 19 47 27 49
rect 19 45 22 47
rect 24 45 27 47
rect 19 43 27 45
rect 9 37 21 39
rect 15 35 17 37
rect 19 35 21 37
rect 15 33 21 35
rect 25 36 27 43
rect 31 47 33 54
rect 41 51 43 54
rect 53 51 55 54
rect 63 51 65 54
rect 41 49 55 51
rect 59 49 65 51
rect 75 49 77 56
rect 85 53 87 56
rect 83 50 87 53
rect 31 45 37 47
rect 31 43 33 45
rect 35 43 37 45
rect 31 41 37 43
rect 25 33 28 36
rect 19 30 21 33
rect 26 30 28 33
rect 33 30 35 41
rect 41 39 43 49
rect 59 45 61 49
rect 54 43 61 45
rect 54 41 56 43
rect 58 42 61 43
rect 73 47 79 49
rect 73 45 75 47
rect 77 45 79 47
rect 73 43 79 45
rect 58 41 60 42
rect 73 41 75 43
rect 54 39 60 41
rect 65 39 75 41
rect 83 39 85 50
rect 41 37 47 39
rect 41 36 43 37
rect 40 35 43 36
rect 45 35 47 37
rect 40 33 52 35
rect 40 30 42 33
rect 50 30 52 33
rect 57 30 59 39
rect 65 36 67 39
rect 64 33 67 36
rect 81 37 87 39
rect 81 35 83 37
rect 85 35 87 37
rect 71 33 87 35
rect 64 30 66 33
rect 71 30 73 33
rect 19 6 21 11
rect 26 6 28 11
rect 33 6 35 11
rect 40 6 42 11
rect 50 6 52 11
rect 57 6 59 11
rect 64 6 66 11
rect 71 6 73 11
<< ndif >>
rect 10 14 19 30
rect 10 12 13 14
rect 15 12 19 14
rect 10 11 19 12
rect 21 11 26 30
rect 28 11 33 30
rect 35 11 40 30
rect 42 21 50 30
rect 42 19 45 21
rect 47 19 50 21
rect 42 11 50 19
rect 52 11 57 30
rect 59 11 64 30
rect 66 11 71 30
rect 73 15 81 30
rect 73 13 76 15
rect 78 13 81 15
rect 73 11 81 13
rect 10 9 17 11
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 52 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 52 19 59
rect 21 68 31 70
rect 21 66 25 68
rect 27 66 31 68
rect 21 54 31 66
rect 33 61 41 70
rect 33 59 36 61
rect 38 59 41 61
rect 33 54 41 59
rect 43 68 53 70
rect 43 66 47 68
rect 49 66 53 68
rect 43 54 53 66
rect 55 61 63 70
rect 55 59 58 61
rect 60 59 63 61
rect 55 54 63 59
rect 65 68 75 70
rect 65 66 69 68
rect 71 66 75 68
rect 65 56 75 66
rect 77 61 85 70
rect 77 59 80 61
rect 82 59 85 61
rect 77 56 85 59
rect 87 68 94 70
rect 87 66 90 68
rect 92 66 94 68
rect 87 60 94 66
rect 87 58 90 60
rect 92 58 94 60
rect 87 56 94 58
rect 65 54 73 56
rect 21 52 29 54
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 12 61 84 62
rect 12 59 14 61
rect 16 59 36 61
rect 38 59 58 61
rect 60 59 80 61
rect 82 59 84 61
rect 12 58 84 59
rect 12 55 16 58
rect 2 50 16 55
rect 21 50 78 54
rect 2 22 6 50
rect 21 47 25 50
rect 21 46 22 47
rect 17 45 22 46
rect 24 45 25 47
rect 74 47 78 50
rect 17 42 25 45
rect 31 45 63 46
rect 31 43 33 45
rect 35 43 63 45
rect 31 42 56 43
rect 58 41 63 43
rect 15 37 27 38
rect 15 35 17 37
rect 19 35 27 37
rect 15 34 27 35
rect 33 37 47 38
rect 33 35 43 37
rect 45 35 47 37
rect 33 34 47 35
rect 57 34 63 41
rect 74 45 75 47
rect 77 45 78 47
rect 23 30 27 34
rect 74 33 78 45
rect 82 37 86 39
rect 82 35 83 37
rect 85 35 86 37
rect 23 26 63 30
rect 2 21 49 22
rect 2 19 45 21
rect 47 19 49 21
rect 2 18 49 19
rect 82 17 86 35
rect -2 1 98 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 19 11 21 30
rect 26 11 28 30
rect 33 11 35 30
rect 40 11 42 30
rect 50 11 52 30
rect 57 11 59 30
rect 64 11 66 30
rect 71 11 73 30
<< pmos >>
rect 9 52 11 70
rect 19 52 21 70
rect 31 54 33 70
rect 41 54 43 70
rect 53 54 55 70
rect 63 54 65 70
rect 75 56 77 70
rect 85 56 87 70
<< polyct0 >>
rect 56 41 57 42
<< polyct1 >>
rect 22 45 24 47
rect 17 35 19 37
rect 33 43 35 45
rect 56 42 58 43
rect 75 45 77 47
rect 57 41 58 42
rect 43 35 45 37
rect 83 35 85 37
<< ndifct0 >>
rect 13 12 15 14
rect 76 13 78 15
<< ndifct1 >>
rect 45 19 47 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 25 66 27 68
rect 47 66 49 68
rect 69 66 71 68
rect 90 66 92 68
rect 90 58 92 60
<< pdifct1 >>
rect 14 59 16 61
rect 36 59 38 61
rect 58 59 60 61
rect 80 59 82 61
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 23 66 25 68
rect 27 66 29 68
rect 23 65 29 66
rect 45 66 47 68
rect 49 66 51 68
rect 45 65 51 66
rect 67 66 69 68
rect 71 66 73 68
rect 67 65 73 66
rect 88 66 90 68
rect 92 66 93 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 88 60 93 66
rect 88 58 90 60
rect 92 58 93 60
rect 55 41 56 42
rect 55 39 57 41
rect 88 42 93 58
rect 63 26 82 29
rect 57 25 82 26
rect 75 15 79 17
rect 11 14 17 15
rect 11 12 13 14
rect 15 12 17 14
rect 75 13 76 15
rect 78 13 79 15
rect 75 12 79 13
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 20 36 20 36 6 a
rlabel alu1 20 44 20 44 6 b
rlabel alu1 28 52 28 52 6 b
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 20 44 20 6 z
rlabel alu1 44 28 44 28 6 a
rlabel alu1 52 28 52 28 6 a
rlabel alu1 36 36 36 36 6 d
rlabel alu1 36 44 36 44 6 c
rlabel polyct1 44 36 44 36 6 d
rlabel alu1 44 44 44 44 6 c
rlabel alu1 52 44 52 44 6 c
rlabel alu1 44 52 44 52 6 b
rlabel alu1 52 52 52 52 6 b
rlabel alu1 36 52 36 52 6 b
rlabel alu1 36 60 36 60 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 52 60 52 60 6 z
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 60 28 60 28 6 a
rlabel alu1 60 40 60 40 6 c
rlabel alu1 76 40 76 40 6 b
rlabel alu1 68 52 68 52 6 b
rlabel alu1 60 52 60 52 6 b
rlabel alu1 60 60 60 60 6 z
rlabel alu1 68 60 68 60 6 z
rlabel alu1 76 60 76 60 6 z
rlabel alu1 84 28 84 28 6 a
<< end >>
