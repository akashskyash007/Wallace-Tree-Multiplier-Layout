magic
tech scmos
timestamp 1199202746
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 63 11 69
rect 19 63 21 69
rect 31 61 33 65
rect 41 61 43 65
rect 9 39 11 44
rect 19 41 21 44
rect 31 41 33 44
rect 19 39 33 41
rect 41 39 43 44
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 27 39
rect 29 37 31 39
rect 19 35 31 37
rect 41 37 47 39
rect 41 35 43 37
rect 45 35 47 37
rect 12 30 14 33
rect 19 30 21 35
rect 29 30 31 35
rect 36 33 47 35
rect 36 30 38 33
rect 12 8 14 13
rect 19 8 21 13
rect 29 12 31 17
rect 36 12 38 17
<< ndif >>
rect 3 13 12 30
rect 14 13 19 30
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 17 29 19
rect 31 17 36 30
rect 38 21 46 30
rect 38 19 41 21
rect 43 19 46 21
rect 38 17 46 19
rect 21 13 26 17
rect 3 11 10 13
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
<< pdif >>
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 44 9 52
rect 11 55 19 63
rect 11 53 14 55
rect 16 53 19 55
rect 11 48 19 53
rect 11 46 14 48
rect 16 46 19 48
rect 11 44 19 46
rect 21 61 29 63
rect 21 59 25 61
rect 27 59 31 61
rect 21 44 31 59
rect 33 59 41 61
rect 33 57 36 59
rect 38 57 41 59
rect 33 52 41 57
rect 33 50 36 52
rect 38 50 41 52
rect 33 44 41 50
rect 43 59 50 61
rect 43 57 46 59
rect 48 57 50 59
rect 43 52 50 57
rect 43 50 46 52
rect 48 50 50 52
rect 43 44 50 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 34 59 40 63
rect 13 55 17 58
rect 13 53 14 55
rect 16 54 17 55
rect 34 57 36 59
rect 38 57 40 59
rect 34 54 40 57
rect 16 53 40 54
rect 13 52 40 53
rect 13 50 36 52
rect 38 50 40 52
rect 13 48 17 50
rect 13 47 14 48
rect 2 46 14 47
rect 16 46 17 48
rect 2 43 17 46
rect 2 22 6 43
rect 25 42 39 46
rect 25 39 31 42
rect 10 37 18 39
rect 10 35 11 37
rect 13 35 18 37
rect 10 33 18 35
rect 25 37 27 39
rect 29 37 31 39
rect 25 34 31 37
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 14 30 18 33
rect 41 30 47 35
rect 14 26 47 30
rect 2 21 31 22
rect 2 19 24 21
rect 26 19 31 21
rect 2 18 31 19
rect -2 11 58 12
rect -2 9 6 11
rect 8 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 12 13 14 30
rect 19 13 21 30
rect 29 17 31 30
rect 36 17 38 30
<< pmos >>
rect 9 44 11 63
rect 19 44 21 63
rect 31 44 33 61
rect 41 44 43 61
<< polyct1 >>
rect 11 35 13 37
rect 27 37 29 39
rect 43 35 45 37
<< ndifct0 >>
rect 41 19 43 21
<< ndifct1 >>
rect 24 19 26 21
rect 6 9 8 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 59 6 61
rect 4 52 6 54
rect 25 59 27 61
rect 46 57 48 59
rect 46 50 48 52
<< pdifct1 >>
rect 14 53 16 55
rect 14 46 16 48
rect 36 57 38 59
rect 36 50 38 52
<< alu0 >>
rect 2 61 8 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 54 8 59
rect 23 61 29 68
rect 23 59 25 61
rect 27 59 29 61
rect 23 58 29 59
rect 2 52 4 54
rect 6 52 8 54
rect 2 51 8 52
rect 34 49 40 50
rect 44 59 50 68
rect 44 57 46 59
rect 48 57 50 59
rect 44 52 50 57
rect 44 50 46 52
rect 48 50 50 52
rect 44 49 50 50
rect 39 21 45 22
rect 39 19 41 21
rect 43 19 45 21
rect 39 12 45 19
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 a
<< end >>
