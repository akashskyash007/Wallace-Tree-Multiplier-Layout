magic
tech scmos
timestamp 1199470235
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 17 85 19 90
rect 25 85 27 90
rect 37 85 39 89
rect 45 85 47 89
rect 17 53 19 65
rect 25 62 27 65
rect 25 59 29 62
rect 27 53 29 59
rect 37 53 39 65
rect 45 62 47 65
rect 45 60 53 62
rect 45 59 49 60
rect 47 58 49 59
rect 51 58 53 60
rect 47 56 53 58
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 11 47 23 49
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 37 51 43 53
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 11 36 13 47
rect 27 41 29 47
rect 37 42 39 47
rect 23 39 29 41
rect 35 39 39 42
rect 23 36 25 39
rect 35 36 37 39
rect 47 36 49 56
rect 11 22 13 27
rect 23 22 25 27
rect 35 22 37 27
rect 47 22 49 27
<< ndif >>
rect 6 33 11 36
rect 3 31 11 33
rect 3 29 5 31
rect 7 29 11 31
rect 3 27 11 29
rect 13 31 23 36
rect 13 29 17 31
rect 19 29 23 31
rect 13 27 23 29
rect 25 31 35 36
rect 25 29 29 31
rect 31 29 35 31
rect 25 27 35 29
rect 37 27 47 36
rect 49 33 54 36
rect 49 31 57 33
rect 49 29 53 31
rect 55 29 57 31
rect 49 27 57 29
rect 39 21 45 27
rect 39 19 41 21
rect 43 19 45 21
rect 39 16 45 19
<< pdif >>
rect 8 91 15 93
rect 8 89 11 91
rect 13 89 15 91
rect 8 85 15 89
rect 8 65 17 85
rect 19 65 25 85
rect 27 81 37 85
rect 27 79 31 81
rect 33 79 37 81
rect 27 65 37 79
rect 39 65 45 85
rect 47 81 56 85
rect 47 79 51 81
rect 53 79 56 81
rect 47 65 56 79
<< alu1 >>
rect -2 95 62 100
rect -2 93 39 95
rect 41 93 49 95
rect 51 93 62 95
rect -2 91 62 93
rect -2 89 11 91
rect 13 89 62 91
rect -2 88 62 89
rect 8 81 34 83
rect 8 79 31 81
rect 33 79 34 81
rect 8 77 34 79
rect 8 43 12 77
rect 38 73 42 83
rect 50 81 54 88
rect 50 79 51 81
rect 53 79 54 81
rect 50 77 54 79
rect 18 67 32 73
rect 38 67 52 73
rect 18 51 22 67
rect 18 49 19 51
rect 21 49 22 51
rect 18 47 22 49
rect 28 51 32 63
rect 28 49 29 51
rect 31 49 32 51
rect 28 43 32 49
rect 38 52 42 63
rect 48 60 52 67
rect 48 58 49 60
rect 51 58 52 60
rect 48 56 52 58
rect 38 51 53 52
rect 38 49 39 51
rect 41 49 53 51
rect 38 47 53 49
rect 8 37 22 43
rect 28 37 42 43
rect 48 37 53 47
rect 4 31 8 33
rect 4 29 5 31
rect 7 29 8 31
rect 4 22 8 29
rect 16 31 22 37
rect 16 29 17 31
rect 19 29 22 31
rect 16 27 22 29
rect 27 31 57 32
rect 27 29 29 31
rect 31 29 53 31
rect 55 29 57 31
rect 27 28 57 29
rect 27 22 31 28
rect 4 18 31 22
rect 40 21 44 23
rect 40 19 41 21
rect 43 19 44 21
rect 40 12 44 19
rect -2 7 62 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 62 7
rect -2 0 62 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 37 95 53 97
rect 37 93 39 95
rect 41 93 49 95
rect 51 93 53 95
rect 37 91 53 93
<< nmos >>
rect 11 27 13 36
rect 23 27 25 36
rect 35 27 37 36
rect 47 27 49 36
<< pmos >>
rect 17 65 19 85
rect 25 65 27 85
rect 37 65 39 85
rect 45 65 47 85
<< polyct1 >>
rect 49 58 51 60
rect 19 49 21 51
rect 29 49 31 51
rect 39 49 41 51
<< ndifct1 >>
rect 5 29 7 31
rect 17 29 19 31
rect 29 29 31 31
rect 53 29 55 31
rect 41 19 43 21
<< ntiect1 >>
rect 39 93 41 95
rect 49 93 51 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 11 89 13 91
rect 31 79 33 81
rect 51 79 53 81
<< labels >>
rlabel ndifct1 6 30 6 30 6 n3
rlabel ndifct1 30 30 30 30 6 n3
rlabel ndifct1 54 30 54 30 6 n3
rlabel alu1 10 60 10 60 6 z
rlabel alu1 20 35 20 35 6 z
rlabel alu1 20 60 20 60 6 b1
rlabel alu1 20 80 20 80 6 z
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 40 40 40 40 6 b2
rlabel polyct1 30 50 30 50 6 b2
rlabel alu1 30 70 30 70 6 b1
rlabel alu1 40 55 40 55 6 a2
rlabel alu1 40 75 40 75 6 a1
rlabel alu1 30 80 30 80 6 z
rlabel alu1 30 94 30 94 6 vdd
rlabel alu1 50 45 50 45 6 a2
rlabel alu1 50 65 50 65 6 a1
<< end >>
