magic
tech scmos
timestamp 1199973087
<< ab >>
rect 0 0 32 88
<< nwell >>
rect -5 40 37 97
<< pwell >>
rect -5 -9 37 40
<< poly >>
rect 2 81 11 83
rect 2 79 7 81
rect 9 79 11 81
rect 2 77 11 79
rect 9 74 11 77
rect 21 81 30 83
rect 21 79 23 81
rect 25 79 30 81
rect 21 77 30 79
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 37 14 43
rect 18 37 30 43
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndif >>
rect 2 14 9 34
rect 11 14 21 34
rect 23 14 30 34
rect 13 9 19 14
rect 13 7 15 9
rect 17 7 19 9
rect 13 2 19 7
<< pdif >>
rect 13 81 19 86
rect 13 79 15 81
rect 17 79 19 81
rect 13 74 19 79
rect 2 46 9 74
rect 11 46 21 74
rect 23 46 30 74
<< alu1 >>
rect -2 89 34 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 34 89
rect -2 86 34 87
rect 5 81 27 82
rect 5 79 7 81
rect 9 79 15 81
rect 17 79 23 81
rect 25 79 27 81
rect 5 78 27 79
rect 13 9 19 10
rect 13 7 15 9
rect 17 7 19 9
rect 13 2 19 7
rect -2 1 34 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< alu2 >>
rect -2 89 34 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 34 89
rect -2 81 34 87
rect -2 79 7 81
rect 9 79 15 81
rect 17 79 23 81
rect 25 79 34 81
rect -2 76 34 79
rect -2 9 34 12
rect -2 7 15 9
rect 17 7 34 9
rect -2 1 34 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 32 3
rect 25 -1 27 1
rect 29 -1 32 1
rect 25 -3 32 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 32 91
rect 25 87 27 89
rect 29 87 32 89
rect 25 85 32 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
<< polyct1 >>
rect 7 79 9 81
rect 23 79 25 81
<< ndifct1 >>
rect 15 7 17 9
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
<< pdifct1 >>
rect 15 79 17 81
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 7 79 9 81
rect 15 79 17 81
rect 23 79 25 81
rect 15 7 17 9
rect 7 -1 9 1
rect 23 -1 25 1
<< labels >>
rlabel alu2 16 6 16 6 6 vss
rlabel alu2 16 82 16 82 6 vdd
<< end >>
