magic
tech scmos
timestamp 1199201633
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 19 61 25 63
rect 19 59 21 61
rect 23 59 25 61
rect 9 54 11 59
rect 19 57 25 59
rect 19 52 21 57
rect 29 52 31 57
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 19 36 23 39
rect 9 33 15 35
rect 9 25 11 33
rect 21 22 23 36
rect 29 31 31 42
rect 28 29 34 31
rect 28 27 30 29
rect 32 27 34 29
rect 28 25 34 27
rect 28 22 30 25
rect 9 15 11 19
rect 21 8 23 13
rect 28 8 30 13
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 22 19 25
rect 11 19 21 22
rect 13 13 21 19
rect 23 13 28 22
rect 30 20 37 22
rect 30 18 33 20
rect 35 18 37 20
rect 30 16 37 18
rect 30 13 35 16
rect 13 11 19 13
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 4 48 9 54
rect 2 46 9 48
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 52 17 54
rect 11 46 19 52
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 46 29 52
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 50 38 52
rect 31 48 34 50
rect 36 48 38 50
rect 31 42 38 48
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 46 6 55
rect 2 44 4 46
rect 2 23 6 44
rect 17 61 30 63
rect 17 59 21 61
rect 23 59 30 61
rect 17 57 30 59
rect 17 50 23 57
rect 2 21 4 23
rect 6 21 14 23
rect 2 17 14 21
rect 34 30 38 39
rect 25 29 38 30
rect 25 27 30 29
rect 32 27 38 29
rect 25 25 38 27
rect -2 11 42 12
rect -2 9 15 11
rect 17 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 19 11 25
rect 21 13 23 22
rect 28 13 30 22
<< pmos >>
rect 9 42 11 54
rect 19 42 21 52
rect 29 42 31 52
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 21 59 23 61
rect 30 27 32 29
<< ndifct0 >>
rect 33 18 35 20
<< ndifct1 >>
rect 4 21 6 23
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 44 16 46
rect 24 44 26 46
rect 34 48 36 50
<< pdifct1 >>
rect 4 44 6 46
<< alu0 >>
rect 6 42 7 48
rect 10 47 14 68
rect 33 50 37 68
rect 33 48 34 50
rect 36 48 37 50
rect 10 46 18 47
rect 10 44 14 46
rect 16 44 18 46
rect 10 43 18 44
rect 22 46 28 47
rect 33 46 37 48
rect 22 44 24 46
rect 26 44 28 46
rect 22 38 28 44
rect 9 37 28 38
rect 9 35 11 37
rect 13 35 28 37
rect 9 34 28 35
rect 6 23 7 25
rect 18 21 22 34
rect 18 20 37 21
rect 18 18 33 20
rect 35 18 37 20
rect 18 17 37 18
<< labels >>
rlabel alu0 18 36 18 36 6 zn
rlabel alu0 25 40 25 40 6 zn
rlabel alu0 27 19 27 19 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 28 28 28 6 b
rlabel alu1 20 56 20 56 6 a
rlabel alu1 28 60 28 60 6 a
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 32 36 32 6 b
<< end >>
