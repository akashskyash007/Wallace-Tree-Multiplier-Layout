magic
tech scmos
timestamp 1199201705
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 58 11 63
rect 19 57 21 61
rect 29 57 31 61
rect 41 58 43 62
rect 9 36 11 46
rect 9 34 15 36
rect 9 32 11 34
rect 13 32 15 34
rect 9 30 15 32
rect 19 35 21 46
rect 29 43 31 46
rect 29 41 37 43
rect 29 40 33 41
rect 31 39 33 40
rect 35 39 37 41
rect 31 37 37 39
rect 19 33 26 35
rect 19 31 21 33
rect 23 31 26 33
rect 9 26 11 30
rect 19 29 26 31
rect 24 26 26 29
rect 31 26 33 37
rect 41 35 43 47
rect 41 33 47 35
rect 41 31 43 33
rect 45 31 47 33
rect 38 29 47 31
rect 38 26 40 29
rect 9 15 11 20
rect 24 10 26 15
rect 31 10 33 15
rect 38 11 40 15
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 11 20 24 26
rect 13 15 24 20
rect 26 15 31 26
rect 33 15 38 26
rect 40 21 45 26
rect 40 19 47 21
rect 40 17 43 19
rect 45 17 47 19
rect 40 15 47 17
rect 13 7 22 15
rect 13 5 16 7
rect 18 5 22 7
rect 13 3 22 5
<< pdif >>
rect 13 67 19 69
rect 13 65 15 67
rect 17 65 19 67
rect 13 63 19 65
rect 33 67 39 69
rect 33 65 35 67
rect 37 65 39 67
rect 13 58 17 63
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 52 9 54
rect 4 46 9 52
rect 11 57 17 58
rect 33 58 39 65
rect 33 57 41 58
rect 11 46 19 57
rect 21 50 29 57
rect 21 48 24 50
rect 26 48 29 50
rect 21 46 29 48
rect 31 47 41 57
rect 43 56 50 58
rect 43 54 46 56
rect 48 54 50 56
rect 43 52 50 54
rect 43 47 48 52
rect 31 46 39 47
<< alu1 >>
rect -2 67 58 72
rect -2 65 15 67
rect 17 65 25 67
rect 27 65 35 67
rect 37 65 58 67
rect -2 64 58 65
rect 2 56 14 59
rect 2 54 4 56
rect 6 54 14 56
rect 2 53 14 54
rect 2 24 6 53
rect 33 46 47 50
rect 33 42 37 46
rect 25 41 37 42
rect 25 39 33 41
rect 35 39 37 41
rect 25 38 37 39
rect 41 34 47 42
rect 2 22 4 24
rect 2 13 6 22
rect 17 33 30 34
rect 17 31 21 33
rect 23 31 30 33
rect 17 30 30 31
rect 26 21 30 30
rect 34 33 47 34
rect 34 31 43 33
rect 45 31 47 33
rect 34 30 47 31
rect 34 21 38 30
rect -2 7 58 8
rect -2 5 5 7
rect 7 5 16 7
rect 18 5 37 7
rect 39 5 45 7
rect 47 5 58 7
rect -2 0 58 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 35 7 49 9
rect 35 5 37 7
rect 39 5 45 7
rect 47 5 49 7
rect 35 3 49 5
<< ntie >>
rect 23 67 29 69
rect 23 65 25 67
rect 27 65 29 67
rect 23 63 29 65
<< nmos >>
rect 9 20 11 26
rect 24 15 26 26
rect 31 15 33 26
rect 38 15 40 26
<< pmos >>
rect 9 46 11 58
rect 19 46 21 57
rect 29 46 31 57
rect 41 47 43 58
<< polyct0 >>
rect 11 32 13 34
<< polyct1 >>
rect 33 39 35 41
rect 21 31 23 33
rect 43 31 45 33
<< ndifct0 >>
rect 43 17 45 19
<< ndifct1 >>
rect 4 22 6 24
rect 16 5 18 7
<< ntiect1 >>
rect 25 65 27 67
<< ptiect1 >>
rect 5 5 7 7
rect 37 5 39 7
rect 45 5 47 7
<< pdifct0 >>
rect 24 48 26 50
rect 46 54 48 56
<< pdifct1 >>
rect 15 65 17 67
rect 35 65 37 67
rect 4 54 6 56
<< alu0 >>
rect 23 56 50 57
rect 23 54 46 56
rect 48 54 50 56
rect 23 53 50 54
rect 23 50 27 53
rect 10 48 24 50
rect 26 48 27 50
rect 10 46 27 48
rect 10 34 14 46
rect 10 32 11 34
rect 13 32 14 34
rect 6 20 7 26
rect 10 25 14 32
rect 10 21 19 25
rect 15 17 19 21
rect 42 19 46 21
rect 42 17 43 19
rect 45 17 46 19
rect 15 13 46 17
<< labels >>
rlabel alu0 12 35 12 35 6 zn
rlabel alu0 25 51 25 51 6 zn
rlabel alu0 44 17 44 17 6 zn
rlabel alu0 36 55 36 55 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 32 20 32 6 a
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 24 28 24 6 a
rlabel alu1 36 24 36 24 6 c
rlabel alu1 28 40 28 40 6 b
rlabel alu1 36 48 36 48 6 b
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 36 44 36 6 c
rlabel alu1 44 48 44 48 6 b
<< end >>
