magic
tech scmos
timestamp 1199203539
<< ab >>
rect 0 0 160 72
<< nwell >>
rect -5 32 165 77
<< pwell >>
rect -5 -5 165 32
<< poly >>
rect 22 66 24 70
rect 29 66 31 70
rect 39 66 41 70
rect 46 66 48 70
rect 56 66 58 70
rect 66 66 68 70
rect 76 66 78 70
rect 86 66 88 70
rect 93 66 95 70
rect 104 68 130 70
rect 104 60 106 68
rect 111 60 113 64
rect 121 60 123 64
rect 128 60 130 68
rect 139 66 141 70
rect 149 66 151 70
rect 22 35 24 38
rect 20 32 24 35
rect 29 35 31 38
rect 39 35 41 38
rect 29 33 42 35
rect 20 26 22 32
rect 29 31 31 33
rect 33 31 38 33
rect 40 31 42 33
rect 29 29 42 31
rect 46 31 48 38
rect 56 35 58 38
rect 66 35 68 38
rect 76 35 78 38
rect 86 35 88 38
rect 56 33 78 35
rect 82 33 88 35
rect 93 35 95 38
rect 104 35 106 38
rect 93 33 106 35
rect 46 29 52 31
rect 30 26 32 29
rect 40 26 42 29
rect 50 26 52 29
rect 72 27 74 33
rect 82 31 84 33
rect 86 31 88 33
rect 82 29 88 31
rect 72 25 78 27
rect 72 23 74 25
rect 76 23 78 25
rect 72 21 78 23
rect 82 19 84 29
rect 104 24 106 33
rect 111 35 113 38
rect 121 35 123 38
rect 128 35 130 38
rect 139 35 141 38
rect 149 35 151 38
rect 111 33 123 35
rect 127 33 133 35
rect 111 31 113 33
rect 115 31 117 33
rect 111 29 117 31
rect 127 31 129 33
rect 131 31 133 33
rect 127 29 133 31
rect 137 33 151 35
rect 137 31 139 33
rect 141 31 143 33
rect 137 29 143 31
rect 92 22 106 24
rect 92 19 94 22
rect 104 19 106 22
rect 114 19 116 29
rect 137 24 139 29
rect 127 22 139 24
rect 127 19 129 22
rect 137 19 139 22
rect 59 16 65 18
rect 59 14 61 16
rect 63 14 65 16
rect 59 12 65 14
rect 20 4 22 12
rect 30 8 32 12
rect 40 8 42 12
rect 50 9 52 12
rect 59 9 61 12
rect 50 7 61 9
rect 50 4 52 7
rect 20 2 52 4
rect 82 2 84 7
rect 92 2 94 7
rect 104 2 106 7
rect 114 2 116 7
rect 127 2 129 6
rect 137 2 139 6
<< ndif >>
rect 13 24 20 26
rect 13 22 15 24
rect 17 22 20 24
rect 13 20 20 22
rect 15 12 20 20
rect 22 24 30 26
rect 22 22 25 24
rect 27 22 30 24
rect 22 17 30 22
rect 22 15 25 17
rect 27 15 30 17
rect 22 12 30 15
rect 32 16 40 26
rect 32 14 35 16
rect 37 14 40 16
rect 32 12 40 14
rect 42 24 50 26
rect 42 22 45 24
rect 47 22 50 24
rect 42 12 50 22
rect 52 24 59 26
rect 52 22 55 24
rect 57 22 59 24
rect 52 20 59 22
rect 52 12 57 20
rect 74 7 82 19
rect 84 16 92 19
rect 84 14 87 16
rect 89 14 92 16
rect 84 7 92 14
rect 94 7 104 19
rect 106 16 114 19
rect 106 14 109 16
rect 111 14 114 16
rect 106 7 114 14
rect 116 7 127 19
rect 74 5 76 7
rect 78 5 80 7
rect 74 3 80 5
rect 96 5 98 7
rect 100 5 102 7
rect 96 3 102 5
rect 118 5 120 7
rect 122 6 127 7
rect 129 16 137 19
rect 129 14 132 16
rect 134 14 137 16
rect 129 6 137 14
rect 139 7 147 19
rect 139 6 143 7
rect 122 5 124 6
rect 118 3 124 5
rect 141 5 143 6
rect 145 5 147 7
rect 141 3 147 5
<< pdif >>
rect 17 51 22 66
rect 15 49 22 51
rect 15 47 17 49
rect 19 47 22 49
rect 15 42 22 47
rect 15 40 17 42
rect 19 40 22 42
rect 15 38 22 40
rect 24 38 29 66
rect 31 64 39 66
rect 31 62 34 64
rect 36 62 39 64
rect 31 56 39 62
rect 31 54 34 56
rect 36 54 39 56
rect 31 38 39 54
rect 41 38 46 66
rect 48 57 56 66
rect 48 55 51 57
rect 53 55 56 57
rect 48 38 56 55
rect 58 42 66 66
rect 58 40 61 42
rect 63 40 66 42
rect 58 38 66 40
rect 68 57 76 66
rect 68 55 71 57
rect 73 55 76 57
rect 68 38 76 55
rect 78 42 86 66
rect 78 40 81 42
rect 83 40 86 42
rect 78 38 86 40
rect 88 38 93 66
rect 95 64 102 66
rect 95 62 98 64
rect 100 62 102 64
rect 95 60 102 62
rect 132 64 139 66
rect 132 62 134 64
rect 136 62 139 64
rect 132 60 139 62
rect 95 38 104 60
rect 106 38 111 60
rect 113 49 121 60
rect 113 47 116 49
rect 118 47 121 49
rect 113 42 121 47
rect 113 40 116 42
rect 118 40 121 42
rect 113 38 121 40
rect 123 38 128 60
rect 130 57 139 60
rect 130 55 134 57
rect 136 55 139 57
rect 130 38 139 55
rect 141 57 149 66
rect 141 55 144 57
rect 146 55 149 57
rect 141 50 149 55
rect 141 48 144 50
rect 146 48 149 50
rect 141 38 149 48
rect 151 59 158 66
rect 151 57 154 59
rect 156 57 158 59
rect 151 38 158 57
<< alu1 >>
rect -2 67 162 72
rect -2 65 5 67
rect 7 65 162 67
rect -2 64 162 65
rect 42 57 79 58
rect 42 55 51 57
rect 53 55 71 57
rect 73 55 79 57
rect 42 54 79 55
rect 2 42 20 43
rect 42 42 46 54
rect 2 40 17 42
rect 19 40 46 42
rect 2 38 46 40
rect 2 17 6 38
rect 24 24 49 26
rect 24 22 25 24
rect 27 22 45 24
rect 47 22 49 24
rect 24 21 49 22
rect 24 17 28 21
rect 105 34 111 42
rect 130 34 134 43
rect 81 33 117 34
rect 81 31 84 33
rect 86 31 113 33
rect 115 31 117 33
rect 81 30 117 31
rect 121 33 134 34
rect 121 31 129 33
rect 131 31 134 33
rect 121 30 134 31
rect 138 33 142 43
rect 138 31 139 33
rect 141 31 142 33
rect 138 26 142 31
rect 72 25 142 26
rect 72 23 74 25
rect 76 23 142 25
rect 72 22 142 23
rect 2 15 25 17
rect 27 15 28 17
rect 2 13 28 15
rect 122 13 126 22
rect -2 7 162 8
rect -2 5 5 7
rect 7 5 66 7
rect 68 5 76 7
rect 78 5 98 7
rect 100 5 120 7
rect 122 5 143 7
rect 145 5 153 7
rect 155 5 162 7
rect -2 0 162 5
<< ptie >>
rect 3 7 9 26
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 64 7 70 9
rect 64 5 66 7
rect 68 5 70 7
rect 64 3 70 5
rect 151 7 157 26
rect 151 5 153 7
rect 155 5 157 7
rect 151 3 157 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 38 9 65
<< nmos >>
rect 20 12 22 26
rect 30 12 32 26
rect 40 12 42 26
rect 50 12 52 26
rect 82 7 84 19
rect 92 7 94 19
rect 104 7 106 19
rect 114 7 116 19
rect 127 6 129 19
rect 137 6 139 19
<< pmos >>
rect 22 38 24 66
rect 29 38 31 66
rect 39 38 41 66
rect 46 38 48 66
rect 56 38 58 66
rect 66 38 68 66
rect 76 38 78 66
rect 86 38 88 66
rect 93 38 95 66
rect 104 38 106 60
rect 111 38 113 60
rect 121 38 123 60
rect 128 38 130 60
rect 139 38 141 66
rect 149 38 151 66
<< polyct0 >>
rect 31 31 33 33
rect 38 31 40 33
rect 61 14 63 16
<< polyct1 >>
rect 84 31 86 33
rect 74 23 76 25
rect 113 31 115 33
rect 129 31 131 33
rect 139 31 141 33
<< ndifct0 >>
rect 15 22 17 24
rect 35 14 37 16
rect 55 22 57 24
rect 87 14 89 16
rect 109 14 111 16
rect 132 14 134 16
<< ndifct1 >>
rect 25 22 27 24
rect 25 15 27 17
rect 45 22 47 24
rect 76 5 78 7
rect 98 5 100 7
rect 120 5 122 7
rect 143 5 145 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
rect 66 5 68 7
rect 153 5 155 7
<< pdifct0 >>
rect 17 47 19 49
rect 34 62 36 64
rect 34 54 36 56
rect 61 40 63 42
rect 81 40 83 42
rect 98 62 100 64
rect 134 62 136 64
rect 116 47 118 49
rect 116 40 118 42
rect 134 55 136 57
rect 144 55 146 57
rect 144 48 146 50
rect 154 57 156 59
<< pdifct1 >>
rect 17 40 19 42
rect 51 55 53 57
rect 71 55 73 57
<< alu0 >>
rect 33 62 34 64
rect 36 62 37 64
rect 33 56 37 62
rect 96 62 98 64
rect 100 62 102 64
rect 96 61 102 62
rect 132 62 134 64
rect 136 62 138 64
rect 33 54 34 56
rect 36 54 37 56
rect 33 52 37 54
rect 86 54 128 58
rect 132 57 138 62
rect 153 59 157 64
rect 132 55 134 57
rect 136 55 138 57
rect 132 54 138 55
rect 143 57 148 58
rect 143 55 144 57
rect 146 55 148 57
rect 153 57 154 59
rect 156 57 157 59
rect 153 55 157 57
rect 16 49 20 51
rect 16 47 17 49
rect 19 47 20 49
rect 16 43 20 47
rect 86 51 90 54
rect 50 47 90 51
rect 124 51 128 54
rect 143 51 148 55
rect 124 50 150 51
rect 94 49 120 50
rect 94 47 116 49
rect 118 47 120 49
rect 124 48 144 50
rect 146 48 150 50
rect 124 47 150 48
rect 50 34 54 47
rect 94 46 120 47
rect 94 43 98 46
rect 59 42 98 43
rect 115 42 120 46
rect 59 40 61 42
rect 63 40 81 42
rect 83 40 98 42
rect 59 39 98 40
rect 13 33 59 34
rect 13 31 31 33
rect 33 31 38 33
rect 40 31 59 33
rect 13 30 59 31
rect 13 24 19 30
rect 13 22 15 24
rect 17 22 19 24
rect 13 21 19 22
rect 53 24 59 30
rect 53 22 55 24
rect 57 22 59 24
rect 53 21 59 22
rect 64 17 68 39
rect 115 40 116 42
rect 118 40 120 42
rect 115 38 120 40
rect 33 16 113 17
rect 33 14 35 16
rect 37 14 61 16
rect 63 14 87 16
rect 89 14 109 16
rect 111 14 113 16
rect 33 13 113 14
rect 146 17 150 47
rect 130 16 150 17
rect 130 14 132 16
rect 134 14 150 16
rect 130 13 150 14
<< labels >>
rlabel alu0 16 27 16 27 6 bn
rlabel alu0 56 27 56 27 6 bn
rlabel alu0 73 15 73 15 6 an
rlabel alu0 78 41 78 41 6 an
rlabel alu0 140 15 140 15 6 bn
rlabel alu0 117 44 117 44 6 an
rlabel alu0 137 49 137 49 6 bn
rlabel alu0 145 52 145 52 6 bn
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 36 24 36 24 6 z
rlabel alu1 44 24 44 24 6 z
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 40 36 40 6 z
rlabel alu1 44 48 44 48 6 z
rlabel pdifct1 52 56 52 56 6 z
rlabel alu1 60 56 60 56 6 z
rlabel alu1 80 4 80 4 6 vss
rlabel alu1 76 24 76 24 6 b
rlabel alu1 84 24 84 24 6 b
rlabel alu1 92 24 92 24 6 b
rlabel alu1 84 32 84 32 6 a2
rlabel alu1 92 32 92 32 6 a2
rlabel alu1 68 56 68 56 6 z
rlabel alu1 76 56 76 56 6 z
rlabel alu1 80 68 80 68 6 vdd
rlabel alu1 100 24 100 24 6 b
rlabel alu1 108 24 108 24 6 b
rlabel alu1 116 24 116 24 6 b
rlabel alu1 124 20 124 20 6 b
rlabel alu1 124 32 124 32 6 a1
rlabel alu1 100 32 100 32 6 a2
rlabel alu1 108 36 108 36 6 a2
rlabel alu1 132 24 132 24 6 b
rlabel alu1 132 40 132 40 6 a1
rlabel alu1 140 36 140 36 6 b
<< end >>
