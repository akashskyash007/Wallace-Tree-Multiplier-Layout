magic
tech scmos
timestamp 1199202426
<< ab >>
rect 0 0 24 72
<< nwell >>
rect -5 32 29 77
<< pwell >>
rect -5 -5 29 32
<< poly >>
rect 13 56 15 61
rect 13 35 15 41
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 9 25 11 29
rect 9 13 11 18
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 18 9 21
rect 11 18 19 25
rect 13 17 19 18
rect 13 15 15 17
rect 17 15 19 17
rect 13 13 19 15
<< pdif >>
rect 5 57 11 59
rect 5 55 7 57
rect 9 56 11 57
rect 9 55 13 56
rect 5 41 13 55
rect 15 51 20 56
rect 15 49 22 51
rect 15 47 18 49
rect 20 47 22 49
rect 15 45 22 47
rect 15 41 20 45
<< alu1 >>
rect -2 67 26 72
rect -2 65 5 67
rect 7 65 17 67
rect 19 65 26 67
rect -2 64 26 65
rect 2 49 22 50
rect 2 47 18 49
rect 20 47 22 49
rect 2 46 22 47
rect 2 25 6 46
rect 10 33 22 35
rect 10 31 11 33
rect 13 31 22 33
rect 10 29 22 31
rect 2 23 7 25
rect 2 21 4 23
rect 6 21 7 23
rect 18 21 22 29
rect 2 19 7 21
rect -2 7 26 8
rect -2 5 5 7
rect 7 5 17 7
rect 19 5 26 7
rect -2 0 26 5
<< ptie >>
rect 3 7 21 9
rect 3 5 5 7
rect 7 5 17 7
rect 19 5 21 7
rect 3 3 21 5
<< ntie >>
rect 3 67 21 69
rect 3 65 5 67
rect 7 65 17 67
rect 19 65 21 67
rect 3 63 21 65
<< nmos >>
rect 9 18 11 25
<< pmos >>
rect 13 41 15 56
<< polyct1 >>
rect 11 31 13 33
<< ndifct0 >>
rect 15 15 17 17
<< ndifct1 >>
rect 4 21 6 23
<< ntiect1 >>
rect 5 65 7 67
rect 17 65 19 67
<< ptiect1 >>
rect 5 5 7 7
rect 17 5 19 7
<< pdifct0 >>
rect 7 55 9 57
<< pdifct1 >>
rect 18 47 20 49
<< alu0 >>
rect 5 57 11 64
rect 5 55 7 57
rect 9 55 11 57
rect 5 54 11 55
rect 13 17 19 18
rect 13 15 15 17
rect 17 15 19 17
rect 13 8 19 15
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 4 12 4 6 vss
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 12 48 12 48 6 z
rlabel alu1 12 68 12 68 6 vdd
rlabel alu1 20 28 20 28 6 a
<< end >>
