magic
tech scmos
timestamp 1635220242
<< ab >>
rect 5 -67 149 77
rect 153 -67 297 77
rect 301 -67 445 77
rect 449 -67 593 77
rect 597 -67 741 77
rect 745 -67 1037 77
rect 1041 -67 1185 77
rect 124 -139 148 -67
<< nwell >>
rect 0 37 1190 82
rect 0 -72 1190 -27
rect 119 -107 153 -72
<< pwell >>
rect 0 -27 1190 37
rect 119 -144 153 -107
<< poly >>
rect 14 71 16 75
rect 60 73 116 75
rect 60 65 62 73
rect 70 65 72 69
rect 80 65 82 69
rect 87 65 89 73
rect 97 65 99 69
rect 104 65 106 69
rect 24 57 26 62
rect 43 59 45 64
rect 50 59 52 64
rect 14 39 16 43
rect 24 40 26 43
rect 14 37 20 39
rect 24 38 39 40
rect 14 35 16 37
rect 18 35 20 37
rect 14 33 20 35
rect 32 36 35 38
rect 37 36 39 38
rect 32 34 39 36
rect 14 29 16 33
rect 32 31 34 34
rect 43 24 45 53
rect 50 49 52 53
rect 50 47 56 49
rect 50 45 52 47
rect 54 45 56 47
rect 50 43 56 45
rect 60 39 62 53
rect 50 37 62 39
rect 50 24 52 37
rect 70 34 72 53
rect 80 49 82 59
rect 76 47 82 49
rect 76 45 78 47
rect 80 45 82 47
rect 76 43 82 45
rect 56 31 62 33
rect 56 29 58 31
rect 60 29 62 31
rect 56 27 62 29
rect 60 24 62 27
rect 70 32 76 34
rect 70 30 72 32
rect 74 30 76 32
rect 70 28 76 30
rect 70 24 72 28
rect 80 24 82 43
rect 87 39 89 59
rect 114 63 116 73
rect 162 71 164 75
rect 134 64 136 69
rect 97 49 99 52
rect 93 47 99 49
rect 93 45 95 47
rect 97 45 99 47
rect 93 43 99 45
rect 104 40 106 52
rect 114 49 116 52
rect 134 50 136 54
rect 114 47 122 49
rect 120 40 122 47
rect 127 48 136 50
rect 127 46 129 48
rect 131 46 136 48
rect 127 44 136 46
rect 87 37 99 39
rect 87 31 93 33
rect 87 29 89 31
rect 91 29 93 31
rect 87 27 93 29
rect 87 24 89 27
rect 97 24 99 37
rect 104 38 110 40
rect 104 36 106 38
rect 108 36 110 38
rect 104 34 110 36
rect 120 38 126 40
rect 120 36 122 38
rect 124 36 126 38
rect 120 34 126 36
rect 104 24 106 34
rect 124 31 126 34
rect 134 31 136 44
rect 208 73 264 75
rect 208 65 210 73
rect 218 65 220 69
rect 228 65 230 69
rect 235 65 237 73
rect 245 65 247 69
rect 252 65 254 69
rect 172 57 174 62
rect 191 59 193 64
rect 198 59 200 64
rect 162 39 164 43
rect 172 40 174 43
rect 162 37 168 39
rect 172 38 187 40
rect 162 35 164 37
rect 166 35 168 37
rect 162 33 168 35
rect 180 36 183 38
rect 185 36 187 38
rect 180 34 187 36
rect 32 19 34 24
rect 124 20 126 25
rect 162 29 164 33
rect 180 31 182 34
rect 134 19 136 24
rect 14 12 16 15
rect 43 12 45 18
rect 50 13 52 18
rect 14 10 45 12
rect 60 9 62 18
rect 70 13 72 18
rect 80 13 82 18
rect 87 9 89 18
rect 97 13 99 18
rect 104 13 106 18
rect 191 24 193 53
rect 198 49 200 53
rect 198 47 204 49
rect 198 45 200 47
rect 202 45 204 47
rect 198 43 204 45
rect 208 39 210 53
rect 198 37 210 39
rect 198 24 200 37
rect 218 34 220 53
rect 228 49 230 59
rect 224 47 230 49
rect 224 45 226 47
rect 228 45 230 47
rect 224 43 230 45
rect 204 31 210 33
rect 204 29 206 31
rect 208 29 210 31
rect 204 27 210 29
rect 208 24 210 27
rect 218 32 224 34
rect 218 30 220 32
rect 222 30 224 32
rect 218 28 224 30
rect 218 24 220 28
rect 228 24 230 43
rect 235 39 237 59
rect 262 63 264 73
rect 310 71 312 75
rect 282 64 284 69
rect 245 49 247 52
rect 241 47 247 49
rect 241 45 243 47
rect 245 45 247 47
rect 241 43 247 45
rect 252 40 254 52
rect 262 49 264 52
rect 282 50 284 54
rect 262 47 270 49
rect 268 40 270 47
rect 275 48 284 50
rect 275 46 277 48
rect 279 46 284 48
rect 275 44 284 46
rect 235 37 247 39
rect 235 31 241 33
rect 235 29 237 31
rect 239 29 241 31
rect 235 27 241 29
rect 235 24 237 27
rect 245 24 247 37
rect 252 38 258 40
rect 252 36 254 38
rect 256 36 258 38
rect 252 34 258 36
rect 268 38 274 40
rect 268 36 270 38
rect 272 36 274 38
rect 268 34 274 36
rect 252 24 254 34
rect 272 31 274 34
rect 282 31 284 44
rect 356 73 412 75
rect 356 65 358 73
rect 366 65 368 69
rect 376 65 378 69
rect 383 65 385 73
rect 393 65 395 69
rect 400 65 402 69
rect 320 57 322 62
rect 339 59 341 64
rect 346 59 348 64
rect 310 39 312 43
rect 320 40 322 43
rect 310 37 316 39
rect 320 38 335 40
rect 310 35 312 37
rect 314 35 316 37
rect 310 33 316 35
rect 328 36 331 38
rect 333 36 335 38
rect 328 34 335 36
rect 180 19 182 24
rect 272 20 274 25
rect 310 29 312 33
rect 328 31 330 34
rect 282 19 284 24
rect 60 7 89 9
rect 162 12 164 15
rect 191 12 193 18
rect 198 13 200 18
rect 162 10 193 12
rect 208 9 210 18
rect 218 13 220 18
rect 228 13 230 18
rect 235 9 237 18
rect 245 13 247 18
rect 252 13 254 18
rect 339 24 341 53
rect 346 49 348 53
rect 346 47 352 49
rect 346 45 348 47
rect 350 45 352 47
rect 346 43 352 45
rect 356 39 358 53
rect 346 37 358 39
rect 346 24 348 37
rect 366 34 368 53
rect 376 49 378 59
rect 372 47 378 49
rect 372 45 374 47
rect 376 45 378 47
rect 372 43 378 45
rect 352 31 358 33
rect 352 29 354 31
rect 356 29 358 31
rect 352 27 358 29
rect 356 24 358 27
rect 366 32 372 34
rect 366 30 368 32
rect 370 30 372 32
rect 366 28 372 30
rect 366 24 368 28
rect 376 24 378 43
rect 383 39 385 59
rect 410 63 412 73
rect 458 71 460 75
rect 430 64 432 69
rect 393 49 395 52
rect 389 47 395 49
rect 389 45 391 47
rect 393 45 395 47
rect 389 43 395 45
rect 400 40 402 52
rect 410 49 412 52
rect 430 50 432 54
rect 410 47 418 49
rect 416 40 418 47
rect 423 48 432 50
rect 423 46 425 48
rect 427 46 432 48
rect 423 44 432 46
rect 383 37 395 39
rect 383 31 389 33
rect 383 29 385 31
rect 387 29 389 31
rect 383 27 389 29
rect 383 24 385 27
rect 393 24 395 37
rect 400 38 406 40
rect 400 36 402 38
rect 404 36 406 38
rect 400 34 406 36
rect 416 38 422 40
rect 416 36 418 38
rect 420 36 422 38
rect 416 34 422 36
rect 400 24 402 34
rect 420 31 422 34
rect 430 31 432 44
rect 504 73 560 75
rect 504 65 506 73
rect 514 65 516 69
rect 524 65 526 69
rect 531 65 533 73
rect 541 65 543 69
rect 548 65 550 69
rect 468 57 470 62
rect 487 59 489 64
rect 494 59 496 64
rect 458 39 460 43
rect 468 40 470 43
rect 458 37 464 39
rect 468 38 483 40
rect 458 35 460 37
rect 462 35 464 37
rect 458 33 464 35
rect 476 36 479 38
rect 481 36 483 38
rect 476 34 483 36
rect 328 19 330 24
rect 420 20 422 25
rect 458 29 460 33
rect 476 31 478 34
rect 430 19 432 24
rect 208 7 237 9
rect 310 12 312 15
rect 339 12 341 18
rect 346 13 348 18
rect 310 10 341 12
rect 356 9 358 18
rect 366 13 368 18
rect 376 13 378 18
rect 383 9 385 18
rect 393 13 395 18
rect 400 13 402 18
rect 487 24 489 53
rect 494 49 496 53
rect 494 47 500 49
rect 494 45 496 47
rect 498 45 500 47
rect 494 43 500 45
rect 504 39 506 53
rect 494 37 506 39
rect 494 24 496 37
rect 514 34 516 53
rect 524 49 526 59
rect 520 47 526 49
rect 520 45 522 47
rect 524 45 526 47
rect 520 43 526 45
rect 500 31 506 33
rect 500 29 502 31
rect 504 29 506 31
rect 500 27 506 29
rect 504 24 506 27
rect 514 32 520 34
rect 514 30 516 32
rect 518 30 520 32
rect 514 28 520 30
rect 514 24 516 28
rect 524 24 526 43
rect 531 39 533 59
rect 558 63 560 73
rect 606 71 608 75
rect 578 64 580 69
rect 541 49 543 52
rect 537 47 543 49
rect 537 45 539 47
rect 541 45 543 47
rect 537 43 543 45
rect 548 40 550 52
rect 558 49 560 52
rect 578 50 580 54
rect 558 47 566 49
rect 564 40 566 47
rect 571 48 580 50
rect 571 46 573 48
rect 575 46 580 48
rect 571 44 580 46
rect 531 37 543 39
rect 531 31 537 33
rect 531 29 533 31
rect 535 29 537 31
rect 531 27 537 29
rect 531 24 533 27
rect 541 24 543 37
rect 548 38 554 40
rect 548 36 550 38
rect 552 36 554 38
rect 548 34 554 36
rect 564 38 570 40
rect 564 36 566 38
rect 568 36 570 38
rect 564 34 570 36
rect 548 24 550 34
rect 568 31 570 34
rect 578 31 580 44
rect 652 73 708 75
rect 652 65 654 73
rect 662 65 664 69
rect 672 65 674 69
rect 679 65 681 73
rect 689 65 691 69
rect 696 65 698 69
rect 616 57 618 62
rect 635 59 637 64
rect 642 59 644 64
rect 606 39 608 43
rect 616 40 618 43
rect 606 37 612 39
rect 616 38 631 40
rect 606 35 608 37
rect 610 35 612 37
rect 606 33 612 35
rect 624 36 627 38
rect 629 36 631 38
rect 624 34 631 36
rect 476 19 478 24
rect 568 20 570 25
rect 606 29 608 33
rect 624 31 626 34
rect 578 19 580 24
rect 356 7 385 9
rect 458 12 460 15
rect 487 12 489 18
rect 494 13 496 18
rect 458 10 489 12
rect 504 9 506 18
rect 514 13 516 18
rect 524 13 526 18
rect 531 9 533 18
rect 541 13 543 18
rect 548 13 550 18
rect 635 24 637 53
rect 642 49 644 53
rect 642 47 648 49
rect 642 45 644 47
rect 646 45 648 47
rect 642 43 648 45
rect 652 39 654 53
rect 642 37 654 39
rect 642 24 644 37
rect 662 34 664 53
rect 672 49 674 59
rect 668 47 674 49
rect 668 45 670 47
rect 672 45 674 47
rect 668 43 674 45
rect 648 31 654 33
rect 648 29 650 31
rect 652 29 654 31
rect 648 27 654 29
rect 652 24 654 27
rect 662 32 668 34
rect 662 30 664 32
rect 666 30 668 32
rect 662 28 668 30
rect 662 24 664 28
rect 672 24 674 43
rect 679 39 681 59
rect 706 63 708 73
rect 754 71 756 75
rect 726 64 728 69
rect 689 49 691 52
rect 685 47 691 49
rect 685 45 687 47
rect 689 45 691 47
rect 685 43 691 45
rect 696 40 698 52
rect 706 49 708 52
rect 726 50 728 54
rect 706 47 714 49
rect 712 40 714 47
rect 719 48 728 50
rect 719 46 721 48
rect 723 46 728 48
rect 719 44 728 46
rect 679 37 691 39
rect 679 31 685 33
rect 679 29 681 31
rect 683 29 685 31
rect 679 27 685 29
rect 679 24 681 27
rect 689 24 691 37
rect 696 38 702 40
rect 696 36 698 38
rect 700 36 702 38
rect 696 34 702 36
rect 712 38 718 40
rect 712 36 714 38
rect 716 36 718 38
rect 712 34 718 36
rect 696 24 698 34
rect 716 31 718 34
rect 726 31 728 44
rect 800 73 856 75
rect 800 65 802 73
rect 810 65 812 69
rect 820 65 822 69
rect 827 65 829 73
rect 837 65 839 69
rect 844 65 846 69
rect 764 57 766 62
rect 783 59 785 64
rect 790 59 792 64
rect 754 39 756 43
rect 764 40 766 43
rect 754 37 760 39
rect 764 38 779 40
rect 754 35 756 37
rect 758 35 760 37
rect 754 33 760 35
rect 772 36 775 38
rect 777 36 779 38
rect 772 34 779 36
rect 624 19 626 24
rect 716 20 718 25
rect 754 29 756 33
rect 772 31 774 34
rect 726 19 728 24
rect 504 7 533 9
rect 606 12 608 15
rect 635 12 637 18
rect 642 13 644 18
rect 606 10 637 12
rect 652 9 654 18
rect 662 13 664 18
rect 672 13 674 18
rect 679 9 681 18
rect 689 13 691 18
rect 696 13 698 18
rect 783 24 785 53
rect 790 49 792 53
rect 790 47 796 49
rect 790 45 792 47
rect 794 45 796 47
rect 790 43 796 45
rect 800 39 802 53
rect 790 37 802 39
rect 790 24 792 37
rect 810 34 812 53
rect 820 49 822 59
rect 816 47 822 49
rect 816 45 818 47
rect 820 45 822 47
rect 816 43 822 45
rect 796 31 802 33
rect 796 29 798 31
rect 800 29 802 31
rect 796 27 802 29
rect 800 24 802 27
rect 810 32 816 34
rect 810 30 812 32
rect 814 30 816 32
rect 810 28 816 30
rect 810 24 812 28
rect 820 24 822 43
rect 827 39 829 59
rect 854 63 856 73
rect 902 71 904 75
rect 874 64 876 69
rect 837 49 839 52
rect 833 47 839 49
rect 833 45 835 47
rect 837 45 839 47
rect 833 43 839 45
rect 844 40 846 52
rect 854 49 856 52
rect 874 50 876 54
rect 854 47 862 49
rect 860 40 862 47
rect 867 48 876 50
rect 867 46 869 48
rect 871 46 876 48
rect 867 44 876 46
rect 827 37 839 39
rect 827 31 833 33
rect 827 29 829 31
rect 831 29 833 31
rect 827 27 833 29
rect 827 24 829 27
rect 837 24 839 37
rect 844 38 850 40
rect 844 36 846 38
rect 848 36 850 38
rect 844 34 850 36
rect 860 38 866 40
rect 860 36 862 38
rect 864 36 866 38
rect 860 34 866 36
rect 844 24 846 34
rect 864 31 866 34
rect 874 31 876 44
rect 948 73 1004 75
rect 948 65 950 73
rect 958 65 960 69
rect 968 65 970 69
rect 975 65 977 73
rect 985 65 987 69
rect 992 65 994 69
rect 912 57 914 62
rect 931 59 933 64
rect 938 59 940 64
rect 902 39 904 43
rect 912 40 914 43
rect 902 37 908 39
rect 912 38 927 40
rect 902 35 904 37
rect 906 35 908 37
rect 902 33 908 35
rect 920 36 923 38
rect 925 36 927 38
rect 920 34 927 36
rect 772 19 774 24
rect 864 20 866 25
rect 902 29 904 33
rect 920 31 922 34
rect 874 19 876 24
rect 652 7 681 9
rect 754 12 756 15
rect 783 12 785 18
rect 790 13 792 18
rect 754 10 785 12
rect 800 9 802 18
rect 810 13 812 18
rect 820 13 822 18
rect 827 9 829 18
rect 837 13 839 18
rect 844 13 846 18
rect 931 24 933 53
rect 938 49 940 53
rect 938 47 944 49
rect 938 45 940 47
rect 942 45 944 47
rect 938 43 944 45
rect 948 39 950 53
rect 938 37 950 39
rect 938 24 940 37
rect 958 34 960 53
rect 968 49 970 59
rect 964 47 970 49
rect 964 45 966 47
rect 968 45 970 47
rect 964 43 970 45
rect 944 31 950 33
rect 944 29 946 31
rect 948 29 950 31
rect 944 27 950 29
rect 948 24 950 27
rect 958 32 964 34
rect 958 30 960 32
rect 962 30 964 32
rect 958 28 964 30
rect 958 24 960 28
rect 968 24 970 43
rect 975 39 977 59
rect 1002 63 1004 73
rect 1050 71 1052 75
rect 1022 64 1024 69
rect 985 49 987 52
rect 981 47 987 49
rect 981 45 983 47
rect 985 45 987 47
rect 981 43 987 45
rect 992 40 994 52
rect 1002 49 1004 52
rect 1022 50 1024 54
rect 1002 47 1010 49
rect 1008 40 1010 47
rect 1015 48 1024 50
rect 1015 46 1017 48
rect 1019 46 1024 48
rect 1015 44 1024 46
rect 975 37 987 39
rect 975 31 981 33
rect 975 29 977 31
rect 979 29 981 31
rect 975 27 981 29
rect 975 24 977 27
rect 985 24 987 37
rect 992 38 998 40
rect 992 36 994 38
rect 996 36 998 38
rect 992 34 998 36
rect 1008 38 1014 40
rect 1008 36 1010 38
rect 1012 36 1014 38
rect 1008 34 1014 36
rect 992 24 994 34
rect 1012 31 1014 34
rect 1022 31 1024 44
rect 1096 73 1152 75
rect 1096 65 1098 73
rect 1106 65 1108 69
rect 1116 65 1118 69
rect 1123 65 1125 73
rect 1133 65 1135 69
rect 1140 65 1142 69
rect 1060 57 1062 62
rect 1079 59 1081 64
rect 1086 59 1088 64
rect 1050 39 1052 43
rect 1060 40 1062 43
rect 1050 37 1056 39
rect 1060 38 1075 40
rect 1050 35 1052 37
rect 1054 35 1056 37
rect 1050 33 1056 35
rect 1068 36 1071 38
rect 1073 36 1075 38
rect 1068 34 1075 36
rect 920 19 922 24
rect 1012 20 1014 25
rect 1050 29 1052 33
rect 1068 31 1070 34
rect 1022 19 1024 24
rect 800 7 829 9
rect 902 12 904 15
rect 931 12 933 18
rect 938 13 940 18
rect 902 10 933 12
rect 948 9 950 18
rect 958 13 960 18
rect 968 13 970 18
rect 975 9 977 18
rect 985 13 987 18
rect 992 13 994 18
rect 1079 24 1081 53
rect 1086 49 1088 53
rect 1086 47 1092 49
rect 1086 45 1088 47
rect 1090 45 1092 47
rect 1086 43 1092 45
rect 1096 39 1098 53
rect 1086 37 1098 39
rect 1086 24 1088 37
rect 1106 34 1108 53
rect 1116 49 1118 59
rect 1112 47 1118 49
rect 1112 45 1114 47
rect 1116 45 1118 47
rect 1112 43 1118 45
rect 1092 31 1098 33
rect 1092 29 1094 31
rect 1096 29 1098 31
rect 1092 27 1098 29
rect 1096 24 1098 27
rect 1106 32 1112 34
rect 1106 30 1108 32
rect 1110 30 1112 32
rect 1106 28 1112 30
rect 1106 24 1108 28
rect 1116 24 1118 43
rect 1123 39 1125 59
rect 1150 63 1152 73
rect 1170 64 1172 69
rect 1133 49 1135 52
rect 1129 47 1135 49
rect 1129 45 1131 47
rect 1133 45 1135 47
rect 1129 43 1135 45
rect 1140 40 1142 52
rect 1150 49 1152 52
rect 1170 50 1172 54
rect 1150 47 1158 49
rect 1156 40 1158 47
rect 1163 48 1172 50
rect 1163 46 1165 48
rect 1167 46 1172 48
rect 1163 44 1172 46
rect 1123 37 1135 39
rect 1123 31 1129 33
rect 1123 29 1125 31
rect 1127 29 1129 31
rect 1123 27 1129 29
rect 1123 24 1125 27
rect 1133 24 1135 37
rect 1140 38 1146 40
rect 1140 36 1142 38
rect 1144 36 1146 38
rect 1140 34 1146 36
rect 1156 38 1162 40
rect 1156 36 1158 38
rect 1160 36 1162 38
rect 1156 34 1162 36
rect 1140 24 1142 34
rect 1160 31 1162 34
rect 1170 31 1172 44
rect 1068 19 1070 24
rect 1160 20 1162 25
rect 1170 19 1172 24
rect 948 7 977 9
rect 1050 12 1052 15
rect 1079 12 1081 18
rect 1086 13 1088 18
rect 1050 10 1081 12
rect 1096 9 1098 18
rect 1106 13 1108 18
rect 1116 13 1118 18
rect 1123 9 1125 18
rect 1133 13 1135 18
rect 1140 13 1142 18
rect 1096 7 1125 9
rect 65 1 94 3
rect 48 -8 50 -3
rect 55 -8 57 -3
rect 65 -8 67 1
rect 72 -8 74 -3
rect 82 -8 84 -3
rect 92 -8 94 1
rect 109 -2 140 0
rect 102 -8 104 -3
rect 109 -8 111 -2
rect 138 -5 140 -2
rect 213 1 242 3
rect 18 -14 20 -9
rect 28 -15 30 -10
rect 120 -14 122 -9
rect 18 -34 20 -21
rect 28 -24 30 -21
rect 48 -24 50 -14
rect 28 -26 34 -24
rect 28 -28 30 -26
rect 32 -28 34 -26
rect 28 -30 34 -28
rect 44 -26 50 -24
rect 44 -28 46 -26
rect 48 -28 50 -26
rect 44 -30 50 -28
rect 55 -27 57 -14
rect 65 -17 67 -14
rect 61 -19 67 -17
rect 61 -21 63 -19
rect 65 -21 67 -19
rect 61 -23 67 -21
rect 55 -29 67 -27
rect 18 -36 27 -34
rect 18 -38 23 -36
rect 25 -38 27 -36
rect 18 -40 27 -38
rect 32 -37 34 -30
rect 32 -39 40 -37
rect 18 -44 20 -40
rect 38 -42 40 -39
rect 48 -42 50 -30
rect 55 -35 61 -33
rect 55 -37 57 -35
rect 59 -37 61 -35
rect 55 -39 61 -37
rect 55 -42 57 -39
rect 18 -59 20 -54
rect 38 -63 40 -53
rect 65 -49 67 -29
rect 72 -33 74 -14
rect 82 -18 84 -14
rect 78 -20 84 -18
rect 78 -22 80 -20
rect 82 -22 84 -20
rect 78 -24 84 -22
rect 92 -17 94 -14
rect 92 -19 98 -17
rect 92 -21 94 -19
rect 96 -21 98 -19
rect 92 -23 98 -21
rect 72 -35 78 -33
rect 72 -37 74 -35
rect 76 -37 78 -35
rect 72 -39 78 -37
rect 72 -49 74 -39
rect 82 -43 84 -24
rect 102 -27 104 -14
rect 92 -29 104 -27
rect 92 -43 94 -29
rect 98 -35 104 -33
rect 98 -37 100 -35
rect 102 -37 104 -35
rect 98 -39 104 -37
rect 102 -43 104 -39
rect 109 -43 111 -14
rect 196 -8 198 -3
rect 203 -8 205 -3
rect 213 -8 215 1
rect 220 -8 222 -3
rect 230 -8 232 -3
rect 240 -8 242 1
rect 257 -2 288 0
rect 250 -8 252 -3
rect 257 -8 259 -2
rect 286 -5 288 -2
rect 361 1 390 3
rect 166 -14 168 -9
rect 120 -24 122 -21
rect 138 -23 140 -19
rect 176 -15 178 -10
rect 268 -14 270 -9
rect 115 -26 122 -24
rect 115 -28 117 -26
rect 119 -28 122 -26
rect 134 -25 140 -23
rect 134 -27 136 -25
rect 138 -27 140 -25
rect 115 -30 130 -28
rect 134 -29 140 -27
rect 128 -33 130 -30
rect 138 -33 140 -29
rect 102 -54 104 -49
rect 109 -54 111 -49
rect 128 -52 130 -47
rect 48 -59 50 -55
rect 55 -59 57 -55
rect 65 -63 67 -55
rect 72 -59 74 -55
rect 82 -59 84 -55
rect 92 -63 94 -55
rect 38 -65 94 -63
rect 166 -34 168 -21
rect 176 -24 178 -21
rect 196 -24 198 -14
rect 176 -26 182 -24
rect 176 -28 178 -26
rect 180 -28 182 -26
rect 176 -30 182 -28
rect 192 -26 198 -24
rect 192 -28 194 -26
rect 196 -28 198 -26
rect 192 -30 198 -28
rect 203 -27 205 -14
rect 213 -17 215 -14
rect 209 -19 215 -17
rect 209 -21 211 -19
rect 213 -21 215 -19
rect 209 -23 215 -21
rect 203 -29 215 -27
rect 166 -36 175 -34
rect 166 -38 171 -36
rect 173 -38 175 -36
rect 166 -40 175 -38
rect 180 -37 182 -30
rect 180 -39 188 -37
rect 166 -44 168 -40
rect 186 -42 188 -39
rect 196 -42 198 -30
rect 203 -35 209 -33
rect 203 -37 205 -35
rect 207 -37 209 -35
rect 203 -39 209 -37
rect 203 -42 205 -39
rect 166 -59 168 -54
rect 138 -65 140 -61
rect 186 -63 188 -53
rect 213 -49 215 -29
rect 220 -33 222 -14
rect 230 -18 232 -14
rect 226 -20 232 -18
rect 226 -22 228 -20
rect 230 -22 232 -20
rect 226 -24 232 -22
rect 240 -17 242 -14
rect 240 -19 246 -17
rect 240 -21 242 -19
rect 244 -21 246 -19
rect 240 -23 246 -21
rect 220 -35 226 -33
rect 220 -37 222 -35
rect 224 -37 226 -35
rect 220 -39 226 -37
rect 220 -49 222 -39
rect 230 -43 232 -24
rect 250 -27 252 -14
rect 240 -29 252 -27
rect 240 -43 242 -29
rect 246 -35 252 -33
rect 246 -37 248 -35
rect 250 -37 252 -35
rect 246 -39 252 -37
rect 250 -43 252 -39
rect 257 -43 259 -14
rect 344 -8 346 -3
rect 351 -8 353 -3
rect 361 -8 363 1
rect 368 -8 370 -3
rect 378 -8 380 -3
rect 388 -8 390 1
rect 405 -2 436 0
rect 398 -8 400 -3
rect 405 -8 407 -2
rect 434 -5 436 -2
rect 509 1 538 3
rect 314 -14 316 -9
rect 268 -24 270 -21
rect 286 -23 288 -19
rect 324 -15 326 -10
rect 416 -14 418 -9
rect 263 -26 270 -24
rect 263 -28 265 -26
rect 267 -28 270 -26
rect 282 -25 288 -23
rect 282 -27 284 -25
rect 286 -27 288 -25
rect 263 -30 278 -28
rect 282 -29 288 -27
rect 276 -33 278 -30
rect 286 -33 288 -29
rect 250 -54 252 -49
rect 257 -54 259 -49
rect 276 -52 278 -47
rect 196 -59 198 -55
rect 203 -59 205 -55
rect 213 -63 215 -55
rect 220 -59 222 -55
rect 230 -59 232 -55
rect 240 -63 242 -55
rect 186 -65 242 -63
rect 314 -34 316 -21
rect 324 -24 326 -21
rect 344 -24 346 -14
rect 324 -26 330 -24
rect 324 -28 326 -26
rect 328 -28 330 -26
rect 324 -30 330 -28
rect 340 -26 346 -24
rect 340 -28 342 -26
rect 344 -28 346 -26
rect 340 -30 346 -28
rect 351 -27 353 -14
rect 361 -17 363 -14
rect 357 -19 363 -17
rect 357 -21 359 -19
rect 361 -21 363 -19
rect 357 -23 363 -21
rect 351 -29 363 -27
rect 314 -36 323 -34
rect 314 -38 319 -36
rect 321 -38 323 -36
rect 314 -40 323 -38
rect 328 -37 330 -30
rect 328 -39 336 -37
rect 314 -44 316 -40
rect 334 -42 336 -39
rect 344 -42 346 -30
rect 351 -35 357 -33
rect 351 -37 353 -35
rect 355 -37 357 -35
rect 351 -39 357 -37
rect 351 -42 353 -39
rect 314 -59 316 -54
rect 286 -65 288 -61
rect 334 -63 336 -53
rect 361 -49 363 -29
rect 368 -33 370 -14
rect 378 -18 380 -14
rect 374 -20 380 -18
rect 374 -22 376 -20
rect 378 -22 380 -20
rect 374 -24 380 -22
rect 388 -17 390 -14
rect 388 -19 394 -17
rect 388 -21 390 -19
rect 392 -21 394 -19
rect 388 -23 394 -21
rect 368 -35 374 -33
rect 368 -37 370 -35
rect 372 -37 374 -35
rect 368 -39 374 -37
rect 368 -49 370 -39
rect 378 -43 380 -24
rect 398 -27 400 -14
rect 388 -29 400 -27
rect 388 -43 390 -29
rect 394 -35 400 -33
rect 394 -37 396 -35
rect 398 -37 400 -35
rect 394 -39 400 -37
rect 398 -43 400 -39
rect 405 -43 407 -14
rect 492 -8 494 -3
rect 499 -8 501 -3
rect 509 -8 511 1
rect 516 -8 518 -3
rect 526 -8 528 -3
rect 536 -8 538 1
rect 553 -2 584 0
rect 546 -8 548 -3
rect 553 -8 555 -2
rect 582 -5 584 -2
rect 657 1 686 3
rect 462 -14 464 -9
rect 416 -24 418 -21
rect 434 -23 436 -19
rect 472 -15 474 -10
rect 564 -14 566 -9
rect 411 -26 418 -24
rect 411 -28 413 -26
rect 415 -28 418 -26
rect 430 -25 436 -23
rect 430 -27 432 -25
rect 434 -27 436 -25
rect 411 -30 426 -28
rect 430 -29 436 -27
rect 424 -33 426 -30
rect 434 -33 436 -29
rect 398 -54 400 -49
rect 405 -54 407 -49
rect 424 -52 426 -47
rect 344 -59 346 -55
rect 351 -59 353 -55
rect 361 -63 363 -55
rect 368 -59 370 -55
rect 378 -59 380 -55
rect 388 -63 390 -55
rect 334 -65 390 -63
rect 462 -34 464 -21
rect 472 -24 474 -21
rect 492 -24 494 -14
rect 472 -26 478 -24
rect 472 -28 474 -26
rect 476 -28 478 -26
rect 472 -30 478 -28
rect 488 -26 494 -24
rect 488 -28 490 -26
rect 492 -28 494 -26
rect 488 -30 494 -28
rect 499 -27 501 -14
rect 509 -17 511 -14
rect 505 -19 511 -17
rect 505 -21 507 -19
rect 509 -21 511 -19
rect 505 -23 511 -21
rect 499 -29 511 -27
rect 462 -36 471 -34
rect 462 -38 467 -36
rect 469 -38 471 -36
rect 462 -40 471 -38
rect 476 -37 478 -30
rect 476 -39 484 -37
rect 462 -44 464 -40
rect 482 -42 484 -39
rect 492 -42 494 -30
rect 499 -35 505 -33
rect 499 -37 501 -35
rect 503 -37 505 -35
rect 499 -39 505 -37
rect 499 -42 501 -39
rect 462 -59 464 -54
rect 434 -65 436 -61
rect 482 -63 484 -53
rect 509 -49 511 -29
rect 516 -33 518 -14
rect 526 -18 528 -14
rect 522 -20 528 -18
rect 522 -22 524 -20
rect 526 -22 528 -20
rect 522 -24 528 -22
rect 536 -17 538 -14
rect 536 -19 542 -17
rect 536 -21 538 -19
rect 540 -21 542 -19
rect 536 -23 542 -21
rect 516 -35 522 -33
rect 516 -37 518 -35
rect 520 -37 522 -35
rect 516 -39 522 -37
rect 516 -49 518 -39
rect 526 -43 528 -24
rect 546 -27 548 -14
rect 536 -29 548 -27
rect 536 -43 538 -29
rect 542 -35 548 -33
rect 542 -37 544 -35
rect 546 -37 548 -35
rect 542 -39 548 -37
rect 546 -43 548 -39
rect 553 -43 555 -14
rect 640 -8 642 -3
rect 647 -8 649 -3
rect 657 -8 659 1
rect 664 -8 666 -3
rect 674 -8 676 -3
rect 684 -8 686 1
rect 701 -2 732 0
rect 694 -8 696 -3
rect 701 -8 703 -2
rect 730 -5 732 -2
rect 805 1 834 3
rect 610 -14 612 -9
rect 564 -24 566 -21
rect 582 -23 584 -19
rect 620 -15 622 -10
rect 712 -14 714 -9
rect 559 -26 566 -24
rect 559 -28 561 -26
rect 563 -28 566 -26
rect 578 -25 584 -23
rect 578 -27 580 -25
rect 582 -27 584 -25
rect 559 -30 574 -28
rect 578 -29 584 -27
rect 572 -33 574 -30
rect 582 -33 584 -29
rect 546 -54 548 -49
rect 553 -54 555 -49
rect 572 -52 574 -47
rect 492 -59 494 -55
rect 499 -59 501 -55
rect 509 -63 511 -55
rect 516 -59 518 -55
rect 526 -59 528 -55
rect 536 -63 538 -55
rect 482 -65 538 -63
rect 610 -34 612 -21
rect 620 -24 622 -21
rect 640 -24 642 -14
rect 620 -26 626 -24
rect 620 -28 622 -26
rect 624 -28 626 -26
rect 620 -30 626 -28
rect 636 -26 642 -24
rect 636 -28 638 -26
rect 640 -28 642 -26
rect 636 -30 642 -28
rect 647 -27 649 -14
rect 657 -17 659 -14
rect 653 -19 659 -17
rect 653 -21 655 -19
rect 657 -21 659 -19
rect 653 -23 659 -21
rect 647 -29 659 -27
rect 610 -36 619 -34
rect 610 -38 615 -36
rect 617 -38 619 -36
rect 610 -40 619 -38
rect 624 -37 626 -30
rect 624 -39 632 -37
rect 610 -44 612 -40
rect 630 -42 632 -39
rect 640 -42 642 -30
rect 647 -35 653 -33
rect 647 -37 649 -35
rect 651 -37 653 -35
rect 647 -39 653 -37
rect 647 -42 649 -39
rect 610 -59 612 -54
rect 582 -65 584 -61
rect 630 -63 632 -53
rect 657 -49 659 -29
rect 664 -33 666 -14
rect 674 -18 676 -14
rect 670 -20 676 -18
rect 670 -22 672 -20
rect 674 -22 676 -20
rect 670 -24 676 -22
rect 684 -17 686 -14
rect 684 -19 690 -17
rect 684 -21 686 -19
rect 688 -21 690 -19
rect 684 -23 690 -21
rect 664 -35 670 -33
rect 664 -37 666 -35
rect 668 -37 670 -35
rect 664 -39 670 -37
rect 664 -49 666 -39
rect 674 -43 676 -24
rect 694 -27 696 -14
rect 684 -29 696 -27
rect 684 -43 686 -29
rect 690 -35 696 -33
rect 690 -37 692 -35
rect 694 -37 696 -35
rect 690 -39 696 -37
rect 694 -43 696 -39
rect 701 -43 703 -14
rect 788 -8 790 -3
rect 795 -8 797 -3
rect 805 -8 807 1
rect 812 -8 814 -3
rect 822 -8 824 -3
rect 832 -8 834 1
rect 849 -2 880 0
rect 842 -8 844 -3
rect 849 -8 851 -2
rect 878 -5 880 -2
rect 953 1 982 3
rect 758 -14 760 -9
rect 712 -24 714 -21
rect 730 -23 732 -19
rect 768 -15 770 -10
rect 860 -14 862 -9
rect 707 -26 714 -24
rect 707 -28 709 -26
rect 711 -28 714 -26
rect 726 -25 732 -23
rect 726 -27 728 -25
rect 730 -27 732 -25
rect 707 -30 722 -28
rect 726 -29 732 -27
rect 720 -33 722 -30
rect 730 -33 732 -29
rect 694 -54 696 -49
rect 701 -54 703 -49
rect 720 -52 722 -47
rect 640 -59 642 -55
rect 647 -59 649 -55
rect 657 -63 659 -55
rect 664 -59 666 -55
rect 674 -59 676 -55
rect 684 -63 686 -55
rect 630 -65 686 -63
rect 758 -34 760 -21
rect 768 -24 770 -21
rect 788 -24 790 -14
rect 768 -26 774 -24
rect 768 -28 770 -26
rect 772 -28 774 -26
rect 768 -30 774 -28
rect 784 -26 790 -24
rect 784 -28 786 -26
rect 788 -28 790 -26
rect 784 -30 790 -28
rect 795 -27 797 -14
rect 805 -17 807 -14
rect 801 -19 807 -17
rect 801 -21 803 -19
rect 805 -21 807 -19
rect 801 -23 807 -21
rect 795 -29 807 -27
rect 758 -36 767 -34
rect 758 -38 763 -36
rect 765 -38 767 -36
rect 758 -40 767 -38
rect 772 -37 774 -30
rect 772 -39 780 -37
rect 758 -44 760 -40
rect 778 -42 780 -39
rect 788 -42 790 -30
rect 795 -35 801 -33
rect 795 -37 797 -35
rect 799 -37 801 -35
rect 795 -39 801 -37
rect 795 -42 797 -39
rect 758 -59 760 -54
rect 730 -65 732 -61
rect 778 -63 780 -53
rect 805 -49 807 -29
rect 812 -33 814 -14
rect 822 -18 824 -14
rect 818 -20 824 -18
rect 818 -22 820 -20
rect 822 -22 824 -20
rect 818 -24 824 -22
rect 832 -17 834 -14
rect 832 -19 838 -17
rect 832 -21 834 -19
rect 836 -21 838 -19
rect 832 -23 838 -21
rect 812 -35 818 -33
rect 812 -37 814 -35
rect 816 -37 818 -35
rect 812 -39 818 -37
rect 812 -49 814 -39
rect 822 -43 824 -24
rect 842 -27 844 -14
rect 832 -29 844 -27
rect 832 -43 834 -29
rect 838 -35 844 -33
rect 838 -37 840 -35
rect 842 -37 844 -35
rect 838 -39 844 -37
rect 842 -43 844 -39
rect 849 -43 851 -14
rect 936 -8 938 -3
rect 943 -8 945 -3
rect 953 -8 955 1
rect 960 -8 962 -3
rect 970 -8 972 -3
rect 980 -8 982 1
rect 997 -2 1028 0
rect 990 -8 992 -3
rect 997 -8 999 -2
rect 1026 -5 1028 -2
rect 1101 1 1130 3
rect 906 -14 908 -9
rect 860 -24 862 -21
rect 878 -23 880 -19
rect 916 -15 918 -10
rect 1008 -14 1010 -9
rect 855 -26 862 -24
rect 855 -28 857 -26
rect 859 -28 862 -26
rect 874 -25 880 -23
rect 874 -27 876 -25
rect 878 -27 880 -25
rect 855 -30 870 -28
rect 874 -29 880 -27
rect 868 -33 870 -30
rect 878 -33 880 -29
rect 842 -54 844 -49
rect 849 -54 851 -49
rect 868 -52 870 -47
rect 788 -59 790 -55
rect 795 -59 797 -55
rect 805 -63 807 -55
rect 812 -59 814 -55
rect 822 -59 824 -55
rect 832 -63 834 -55
rect 778 -65 834 -63
rect 906 -34 908 -21
rect 916 -24 918 -21
rect 936 -24 938 -14
rect 916 -26 922 -24
rect 916 -28 918 -26
rect 920 -28 922 -26
rect 916 -30 922 -28
rect 932 -26 938 -24
rect 932 -28 934 -26
rect 936 -28 938 -26
rect 932 -30 938 -28
rect 943 -27 945 -14
rect 953 -17 955 -14
rect 949 -19 955 -17
rect 949 -21 951 -19
rect 953 -21 955 -19
rect 949 -23 955 -21
rect 943 -29 955 -27
rect 906 -36 915 -34
rect 906 -38 911 -36
rect 913 -38 915 -36
rect 906 -40 915 -38
rect 920 -37 922 -30
rect 920 -39 928 -37
rect 906 -44 908 -40
rect 926 -42 928 -39
rect 936 -42 938 -30
rect 943 -35 949 -33
rect 943 -37 945 -35
rect 947 -37 949 -35
rect 943 -39 949 -37
rect 943 -42 945 -39
rect 906 -59 908 -54
rect 878 -65 880 -61
rect 926 -63 928 -53
rect 953 -49 955 -29
rect 960 -33 962 -14
rect 970 -18 972 -14
rect 966 -20 972 -18
rect 966 -22 968 -20
rect 970 -22 972 -20
rect 966 -24 972 -22
rect 980 -17 982 -14
rect 980 -19 986 -17
rect 980 -21 982 -19
rect 984 -21 986 -19
rect 980 -23 986 -21
rect 960 -35 966 -33
rect 960 -37 962 -35
rect 964 -37 966 -35
rect 960 -39 966 -37
rect 960 -49 962 -39
rect 970 -43 972 -24
rect 990 -27 992 -14
rect 980 -29 992 -27
rect 980 -43 982 -29
rect 986 -35 992 -33
rect 986 -37 988 -35
rect 990 -37 992 -35
rect 986 -39 992 -37
rect 990 -43 992 -39
rect 997 -43 999 -14
rect 1084 -8 1086 -3
rect 1091 -8 1093 -3
rect 1101 -8 1103 1
rect 1108 -8 1110 -3
rect 1118 -8 1120 -3
rect 1128 -8 1130 1
rect 1145 -2 1176 0
rect 1138 -8 1140 -3
rect 1145 -8 1147 -2
rect 1174 -5 1176 -2
rect 1054 -14 1056 -9
rect 1008 -24 1010 -21
rect 1026 -23 1028 -19
rect 1064 -15 1066 -10
rect 1156 -14 1158 -9
rect 1003 -26 1010 -24
rect 1003 -28 1005 -26
rect 1007 -28 1010 -26
rect 1022 -25 1028 -23
rect 1022 -27 1024 -25
rect 1026 -27 1028 -25
rect 1003 -30 1018 -28
rect 1022 -29 1028 -27
rect 1016 -33 1018 -30
rect 1026 -33 1028 -29
rect 990 -54 992 -49
rect 997 -54 999 -49
rect 1016 -52 1018 -47
rect 936 -59 938 -55
rect 943 -59 945 -55
rect 953 -63 955 -55
rect 960 -59 962 -55
rect 970 -59 972 -55
rect 980 -63 982 -55
rect 926 -65 982 -63
rect 1054 -34 1056 -21
rect 1064 -24 1066 -21
rect 1084 -24 1086 -14
rect 1064 -26 1070 -24
rect 1064 -28 1066 -26
rect 1068 -28 1070 -26
rect 1064 -30 1070 -28
rect 1080 -26 1086 -24
rect 1080 -28 1082 -26
rect 1084 -28 1086 -26
rect 1080 -30 1086 -28
rect 1091 -27 1093 -14
rect 1101 -17 1103 -14
rect 1097 -19 1103 -17
rect 1097 -21 1099 -19
rect 1101 -21 1103 -19
rect 1097 -23 1103 -21
rect 1091 -29 1103 -27
rect 1054 -36 1063 -34
rect 1054 -38 1059 -36
rect 1061 -38 1063 -36
rect 1054 -40 1063 -38
rect 1068 -37 1070 -30
rect 1068 -39 1076 -37
rect 1054 -44 1056 -40
rect 1074 -42 1076 -39
rect 1084 -42 1086 -30
rect 1091 -35 1097 -33
rect 1091 -37 1093 -35
rect 1095 -37 1097 -35
rect 1091 -39 1097 -37
rect 1091 -42 1093 -39
rect 1054 -59 1056 -54
rect 1026 -65 1028 -61
rect 1074 -63 1076 -53
rect 1101 -49 1103 -29
rect 1108 -33 1110 -14
rect 1118 -18 1120 -14
rect 1114 -20 1120 -18
rect 1114 -22 1116 -20
rect 1118 -22 1120 -20
rect 1114 -24 1120 -22
rect 1128 -17 1130 -14
rect 1128 -19 1134 -17
rect 1128 -21 1130 -19
rect 1132 -21 1134 -19
rect 1128 -23 1134 -21
rect 1108 -35 1114 -33
rect 1108 -37 1110 -35
rect 1112 -37 1114 -35
rect 1108 -39 1114 -37
rect 1108 -49 1110 -39
rect 1118 -43 1120 -24
rect 1138 -27 1140 -14
rect 1128 -29 1140 -27
rect 1128 -43 1130 -29
rect 1134 -35 1140 -33
rect 1134 -37 1136 -35
rect 1138 -37 1140 -35
rect 1134 -39 1140 -37
rect 1138 -43 1140 -39
rect 1145 -43 1147 -14
rect 1156 -24 1158 -21
rect 1174 -23 1176 -19
rect 1151 -26 1158 -24
rect 1151 -28 1153 -26
rect 1155 -28 1158 -26
rect 1170 -25 1176 -23
rect 1170 -27 1172 -25
rect 1174 -27 1176 -25
rect 1151 -30 1166 -28
rect 1170 -29 1176 -27
rect 1164 -33 1166 -30
rect 1174 -33 1176 -29
rect 1138 -54 1140 -49
rect 1145 -54 1147 -49
rect 1164 -52 1166 -47
rect 1084 -59 1086 -55
rect 1091 -59 1093 -55
rect 1101 -63 1103 -55
rect 1108 -59 1110 -55
rect 1118 -59 1120 -55
rect 1128 -63 1130 -55
rect 1074 -65 1130 -63
rect 1174 -65 1176 -61
rect 133 -83 135 -78
rect 133 -104 135 -101
rect 133 -106 139 -104
rect 133 -108 135 -106
rect 137 -108 139 -106
rect 133 -110 139 -108
rect 133 -113 135 -110
rect 133 -127 135 -122
<< ndif >>
rect 25 29 32 31
rect 7 27 14 29
rect 7 25 9 27
rect 11 25 14 27
rect 7 23 14 25
rect 9 15 14 23
rect 16 21 21 29
rect 25 27 27 29
rect 29 27 32 29
rect 25 25 32 27
rect 27 24 32 25
rect 34 24 41 31
rect 117 29 124 31
rect 117 27 119 29
rect 121 27 124 29
rect 117 25 124 27
rect 126 29 134 31
rect 126 27 129 29
rect 131 27 134 29
rect 126 25 134 27
rect 16 19 23 21
rect 36 22 43 24
rect 36 20 38 22
rect 40 20 43 22
rect 16 17 19 19
rect 21 17 23 19
rect 36 18 43 20
rect 45 18 50 24
rect 52 22 60 24
rect 52 20 55 22
rect 57 20 60 22
rect 52 18 60 20
rect 62 22 70 24
rect 62 20 65 22
rect 67 20 70 22
rect 62 18 70 20
rect 72 22 80 24
rect 72 20 75 22
rect 77 20 80 22
rect 72 18 80 20
rect 82 18 87 24
rect 89 22 97 24
rect 89 20 92 22
rect 94 20 97 22
rect 89 18 97 20
rect 99 18 104 24
rect 106 22 113 24
rect 106 20 109 22
rect 111 20 113 22
rect 128 24 134 25
rect 136 29 143 31
rect 173 29 180 31
rect 136 27 139 29
rect 141 27 143 29
rect 136 24 143 27
rect 155 27 162 29
rect 155 25 157 27
rect 159 25 162 27
rect 106 18 113 20
rect 155 23 162 25
rect 16 15 23 17
rect 157 15 162 23
rect 164 21 169 29
rect 173 27 175 29
rect 177 27 180 29
rect 173 25 180 27
rect 175 24 180 25
rect 182 24 189 31
rect 265 29 272 31
rect 265 27 267 29
rect 269 27 272 29
rect 265 25 272 27
rect 274 29 282 31
rect 274 27 277 29
rect 279 27 282 29
rect 274 25 282 27
rect 164 19 171 21
rect 184 22 191 24
rect 184 20 186 22
rect 188 20 191 22
rect 164 17 167 19
rect 169 17 171 19
rect 184 18 191 20
rect 193 18 198 24
rect 200 22 208 24
rect 200 20 203 22
rect 205 20 208 22
rect 200 18 208 20
rect 210 22 218 24
rect 210 20 213 22
rect 215 20 218 22
rect 210 18 218 20
rect 220 22 228 24
rect 220 20 223 22
rect 225 20 228 22
rect 220 18 228 20
rect 230 18 235 24
rect 237 22 245 24
rect 237 20 240 22
rect 242 20 245 22
rect 237 18 245 20
rect 247 18 252 24
rect 254 22 261 24
rect 254 20 257 22
rect 259 20 261 22
rect 276 24 282 25
rect 284 29 291 31
rect 321 29 328 31
rect 284 27 287 29
rect 289 27 291 29
rect 284 24 291 27
rect 303 27 310 29
rect 303 25 305 27
rect 307 25 310 27
rect 254 18 261 20
rect 303 23 310 25
rect 164 15 171 17
rect 305 15 310 23
rect 312 21 317 29
rect 321 27 323 29
rect 325 27 328 29
rect 321 25 328 27
rect 323 24 328 25
rect 330 24 337 31
rect 413 29 420 31
rect 413 27 415 29
rect 417 27 420 29
rect 413 25 420 27
rect 422 29 430 31
rect 422 27 425 29
rect 427 27 430 29
rect 422 25 430 27
rect 312 19 319 21
rect 332 22 339 24
rect 332 20 334 22
rect 336 20 339 22
rect 312 17 315 19
rect 317 17 319 19
rect 332 18 339 20
rect 341 18 346 24
rect 348 22 356 24
rect 348 20 351 22
rect 353 20 356 22
rect 348 18 356 20
rect 358 22 366 24
rect 358 20 361 22
rect 363 20 366 22
rect 358 18 366 20
rect 368 22 376 24
rect 368 20 371 22
rect 373 20 376 22
rect 368 18 376 20
rect 378 18 383 24
rect 385 22 393 24
rect 385 20 388 22
rect 390 20 393 22
rect 385 18 393 20
rect 395 18 400 24
rect 402 22 409 24
rect 402 20 405 22
rect 407 20 409 22
rect 424 24 430 25
rect 432 29 439 31
rect 469 29 476 31
rect 432 27 435 29
rect 437 27 439 29
rect 432 24 439 27
rect 451 27 458 29
rect 451 25 453 27
rect 455 25 458 27
rect 402 18 409 20
rect 451 23 458 25
rect 312 15 319 17
rect 453 15 458 23
rect 460 21 465 29
rect 469 27 471 29
rect 473 27 476 29
rect 469 25 476 27
rect 471 24 476 25
rect 478 24 485 31
rect 561 29 568 31
rect 561 27 563 29
rect 565 27 568 29
rect 561 25 568 27
rect 570 29 578 31
rect 570 27 573 29
rect 575 27 578 29
rect 570 25 578 27
rect 460 19 467 21
rect 480 22 487 24
rect 480 20 482 22
rect 484 20 487 22
rect 460 17 463 19
rect 465 17 467 19
rect 480 18 487 20
rect 489 18 494 24
rect 496 22 504 24
rect 496 20 499 22
rect 501 20 504 22
rect 496 18 504 20
rect 506 22 514 24
rect 506 20 509 22
rect 511 20 514 22
rect 506 18 514 20
rect 516 22 524 24
rect 516 20 519 22
rect 521 20 524 22
rect 516 18 524 20
rect 526 18 531 24
rect 533 22 541 24
rect 533 20 536 22
rect 538 20 541 22
rect 533 18 541 20
rect 543 18 548 24
rect 550 22 557 24
rect 550 20 553 22
rect 555 20 557 22
rect 572 24 578 25
rect 580 29 587 31
rect 617 29 624 31
rect 580 27 583 29
rect 585 27 587 29
rect 580 24 587 27
rect 599 27 606 29
rect 599 25 601 27
rect 603 25 606 27
rect 550 18 557 20
rect 599 23 606 25
rect 460 15 467 17
rect 601 15 606 23
rect 608 21 613 29
rect 617 27 619 29
rect 621 27 624 29
rect 617 25 624 27
rect 619 24 624 25
rect 626 24 633 31
rect 709 29 716 31
rect 709 27 711 29
rect 713 27 716 29
rect 709 25 716 27
rect 718 29 726 31
rect 718 27 721 29
rect 723 27 726 29
rect 718 25 726 27
rect 608 19 615 21
rect 628 22 635 24
rect 628 20 630 22
rect 632 20 635 22
rect 608 17 611 19
rect 613 17 615 19
rect 628 18 635 20
rect 637 18 642 24
rect 644 22 652 24
rect 644 20 647 22
rect 649 20 652 22
rect 644 18 652 20
rect 654 22 662 24
rect 654 20 657 22
rect 659 20 662 22
rect 654 18 662 20
rect 664 22 672 24
rect 664 20 667 22
rect 669 20 672 22
rect 664 18 672 20
rect 674 18 679 24
rect 681 22 689 24
rect 681 20 684 22
rect 686 20 689 22
rect 681 18 689 20
rect 691 18 696 24
rect 698 22 705 24
rect 698 20 701 22
rect 703 20 705 22
rect 720 24 726 25
rect 728 29 735 31
rect 765 29 772 31
rect 728 27 731 29
rect 733 27 735 29
rect 728 24 735 27
rect 747 27 754 29
rect 747 25 749 27
rect 751 25 754 27
rect 698 18 705 20
rect 747 23 754 25
rect 608 15 615 17
rect 749 15 754 23
rect 756 21 761 29
rect 765 27 767 29
rect 769 27 772 29
rect 765 25 772 27
rect 767 24 772 25
rect 774 24 781 31
rect 857 29 864 31
rect 857 27 859 29
rect 861 27 864 29
rect 857 25 864 27
rect 866 29 874 31
rect 866 27 869 29
rect 871 27 874 29
rect 866 25 874 27
rect 756 19 763 21
rect 776 22 783 24
rect 776 20 778 22
rect 780 20 783 22
rect 756 17 759 19
rect 761 17 763 19
rect 776 18 783 20
rect 785 18 790 24
rect 792 22 800 24
rect 792 20 795 22
rect 797 20 800 22
rect 792 18 800 20
rect 802 22 810 24
rect 802 20 805 22
rect 807 20 810 22
rect 802 18 810 20
rect 812 22 820 24
rect 812 20 815 22
rect 817 20 820 22
rect 812 18 820 20
rect 822 18 827 24
rect 829 22 837 24
rect 829 20 832 22
rect 834 20 837 22
rect 829 18 837 20
rect 839 18 844 24
rect 846 22 853 24
rect 846 20 849 22
rect 851 20 853 22
rect 868 24 874 25
rect 876 29 883 31
rect 913 29 920 31
rect 876 27 879 29
rect 881 27 883 29
rect 876 24 883 27
rect 895 27 902 29
rect 895 25 897 27
rect 899 25 902 27
rect 846 18 853 20
rect 895 23 902 25
rect 756 15 763 17
rect 897 15 902 23
rect 904 21 909 29
rect 913 27 915 29
rect 917 27 920 29
rect 913 25 920 27
rect 915 24 920 25
rect 922 24 929 31
rect 1005 29 1012 31
rect 1005 27 1007 29
rect 1009 27 1012 29
rect 1005 25 1012 27
rect 1014 29 1022 31
rect 1014 27 1017 29
rect 1019 27 1022 29
rect 1014 25 1022 27
rect 904 19 911 21
rect 924 22 931 24
rect 924 20 926 22
rect 928 20 931 22
rect 904 17 907 19
rect 909 17 911 19
rect 924 18 931 20
rect 933 18 938 24
rect 940 22 948 24
rect 940 20 943 22
rect 945 20 948 22
rect 940 18 948 20
rect 950 22 958 24
rect 950 20 953 22
rect 955 20 958 22
rect 950 18 958 20
rect 960 22 968 24
rect 960 20 963 22
rect 965 20 968 22
rect 960 18 968 20
rect 970 18 975 24
rect 977 22 985 24
rect 977 20 980 22
rect 982 20 985 22
rect 977 18 985 20
rect 987 18 992 24
rect 994 22 1001 24
rect 994 20 997 22
rect 999 20 1001 22
rect 1016 24 1022 25
rect 1024 29 1031 31
rect 1061 29 1068 31
rect 1024 27 1027 29
rect 1029 27 1031 29
rect 1024 24 1031 27
rect 1043 27 1050 29
rect 1043 25 1045 27
rect 1047 25 1050 27
rect 994 18 1001 20
rect 1043 23 1050 25
rect 904 15 911 17
rect 1045 15 1050 23
rect 1052 21 1057 29
rect 1061 27 1063 29
rect 1065 27 1068 29
rect 1061 25 1068 27
rect 1063 24 1068 25
rect 1070 24 1077 31
rect 1153 29 1160 31
rect 1153 27 1155 29
rect 1157 27 1160 29
rect 1153 25 1160 27
rect 1162 29 1170 31
rect 1162 27 1165 29
rect 1167 27 1170 29
rect 1162 25 1170 27
rect 1052 19 1059 21
rect 1072 22 1079 24
rect 1072 20 1074 22
rect 1076 20 1079 22
rect 1052 17 1055 19
rect 1057 17 1059 19
rect 1072 18 1079 20
rect 1081 18 1086 24
rect 1088 22 1096 24
rect 1088 20 1091 22
rect 1093 20 1096 22
rect 1088 18 1096 20
rect 1098 22 1106 24
rect 1098 20 1101 22
rect 1103 20 1106 22
rect 1098 18 1106 20
rect 1108 22 1116 24
rect 1108 20 1111 22
rect 1113 20 1116 22
rect 1108 18 1116 20
rect 1118 18 1123 24
rect 1125 22 1133 24
rect 1125 20 1128 22
rect 1130 20 1133 22
rect 1125 18 1133 20
rect 1135 18 1140 24
rect 1142 22 1149 24
rect 1142 20 1145 22
rect 1147 20 1149 22
rect 1164 24 1170 25
rect 1172 29 1179 31
rect 1172 27 1175 29
rect 1177 27 1179 29
rect 1172 24 1179 27
rect 1142 18 1149 20
rect 1052 15 1059 17
rect 131 -7 138 -5
rect 41 -10 48 -8
rect 11 -17 18 -14
rect 11 -19 13 -17
rect 15 -19 18 -17
rect 11 -21 18 -19
rect 20 -15 26 -14
rect 41 -12 43 -10
rect 45 -12 48 -10
rect 41 -14 48 -12
rect 50 -14 55 -8
rect 57 -10 65 -8
rect 57 -12 60 -10
rect 62 -12 65 -10
rect 57 -14 65 -12
rect 67 -14 72 -8
rect 74 -10 82 -8
rect 74 -12 77 -10
rect 79 -12 82 -10
rect 74 -14 82 -12
rect 84 -10 92 -8
rect 84 -12 87 -10
rect 89 -12 92 -10
rect 84 -14 92 -12
rect 94 -10 102 -8
rect 94 -12 97 -10
rect 99 -12 102 -10
rect 94 -14 102 -12
rect 104 -14 109 -8
rect 111 -10 118 -8
rect 131 -9 133 -7
rect 135 -9 138 -7
rect 111 -12 114 -10
rect 116 -12 118 -10
rect 111 -14 118 -12
rect 131 -11 138 -9
rect 20 -17 28 -15
rect 20 -19 23 -17
rect 25 -19 28 -17
rect 20 -21 28 -19
rect 30 -17 37 -15
rect 30 -19 33 -17
rect 35 -19 37 -17
rect 30 -21 37 -19
rect 113 -21 120 -14
rect 122 -15 127 -14
rect 122 -17 129 -15
rect 122 -19 125 -17
rect 127 -19 129 -17
rect 133 -19 138 -11
rect 140 -13 145 -5
rect 279 -7 286 -5
rect 140 -15 147 -13
rect 189 -10 196 -8
rect 140 -17 143 -15
rect 145 -17 147 -15
rect 140 -19 147 -17
rect 159 -17 166 -14
rect 159 -19 161 -17
rect 163 -19 166 -17
rect 122 -21 129 -19
rect 159 -21 166 -19
rect 168 -15 174 -14
rect 189 -12 191 -10
rect 193 -12 196 -10
rect 189 -14 196 -12
rect 198 -14 203 -8
rect 205 -10 213 -8
rect 205 -12 208 -10
rect 210 -12 213 -10
rect 205 -14 213 -12
rect 215 -14 220 -8
rect 222 -10 230 -8
rect 222 -12 225 -10
rect 227 -12 230 -10
rect 222 -14 230 -12
rect 232 -10 240 -8
rect 232 -12 235 -10
rect 237 -12 240 -10
rect 232 -14 240 -12
rect 242 -10 250 -8
rect 242 -12 245 -10
rect 247 -12 250 -10
rect 242 -14 250 -12
rect 252 -14 257 -8
rect 259 -10 266 -8
rect 279 -9 281 -7
rect 283 -9 286 -7
rect 259 -12 262 -10
rect 264 -12 266 -10
rect 259 -14 266 -12
rect 279 -11 286 -9
rect 168 -17 176 -15
rect 168 -19 171 -17
rect 173 -19 176 -17
rect 168 -21 176 -19
rect 178 -17 185 -15
rect 178 -19 181 -17
rect 183 -19 185 -17
rect 178 -21 185 -19
rect 261 -21 268 -14
rect 270 -15 275 -14
rect 270 -17 277 -15
rect 270 -19 273 -17
rect 275 -19 277 -17
rect 281 -19 286 -11
rect 288 -13 293 -5
rect 427 -7 434 -5
rect 288 -15 295 -13
rect 337 -10 344 -8
rect 288 -17 291 -15
rect 293 -17 295 -15
rect 288 -19 295 -17
rect 307 -17 314 -14
rect 307 -19 309 -17
rect 311 -19 314 -17
rect 270 -21 277 -19
rect 307 -21 314 -19
rect 316 -15 322 -14
rect 337 -12 339 -10
rect 341 -12 344 -10
rect 337 -14 344 -12
rect 346 -14 351 -8
rect 353 -10 361 -8
rect 353 -12 356 -10
rect 358 -12 361 -10
rect 353 -14 361 -12
rect 363 -14 368 -8
rect 370 -10 378 -8
rect 370 -12 373 -10
rect 375 -12 378 -10
rect 370 -14 378 -12
rect 380 -10 388 -8
rect 380 -12 383 -10
rect 385 -12 388 -10
rect 380 -14 388 -12
rect 390 -10 398 -8
rect 390 -12 393 -10
rect 395 -12 398 -10
rect 390 -14 398 -12
rect 400 -14 405 -8
rect 407 -10 414 -8
rect 427 -9 429 -7
rect 431 -9 434 -7
rect 407 -12 410 -10
rect 412 -12 414 -10
rect 407 -14 414 -12
rect 427 -11 434 -9
rect 316 -17 324 -15
rect 316 -19 319 -17
rect 321 -19 324 -17
rect 316 -21 324 -19
rect 326 -17 333 -15
rect 326 -19 329 -17
rect 331 -19 333 -17
rect 326 -21 333 -19
rect 409 -21 416 -14
rect 418 -15 423 -14
rect 418 -17 425 -15
rect 418 -19 421 -17
rect 423 -19 425 -17
rect 429 -19 434 -11
rect 436 -13 441 -5
rect 575 -7 582 -5
rect 436 -15 443 -13
rect 485 -10 492 -8
rect 436 -17 439 -15
rect 441 -17 443 -15
rect 436 -19 443 -17
rect 455 -17 462 -14
rect 455 -19 457 -17
rect 459 -19 462 -17
rect 418 -21 425 -19
rect 455 -21 462 -19
rect 464 -15 470 -14
rect 485 -12 487 -10
rect 489 -12 492 -10
rect 485 -14 492 -12
rect 494 -14 499 -8
rect 501 -10 509 -8
rect 501 -12 504 -10
rect 506 -12 509 -10
rect 501 -14 509 -12
rect 511 -14 516 -8
rect 518 -10 526 -8
rect 518 -12 521 -10
rect 523 -12 526 -10
rect 518 -14 526 -12
rect 528 -10 536 -8
rect 528 -12 531 -10
rect 533 -12 536 -10
rect 528 -14 536 -12
rect 538 -10 546 -8
rect 538 -12 541 -10
rect 543 -12 546 -10
rect 538 -14 546 -12
rect 548 -14 553 -8
rect 555 -10 562 -8
rect 575 -9 577 -7
rect 579 -9 582 -7
rect 555 -12 558 -10
rect 560 -12 562 -10
rect 555 -14 562 -12
rect 575 -11 582 -9
rect 464 -17 472 -15
rect 464 -19 467 -17
rect 469 -19 472 -17
rect 464 -21 472 -19
rect 474 -17 481 -15
rect 474 -19 477 -17
rect 479 -19 481 -17
rect 474 -21 481 -19
rect 557 -21 564 -14
rect 566 -15 571 -14
rect 566 -17 573 -15
rect 566 -19 569 -17
rect 571 -19 573 -17
rect 577 -19 582 -11
rect 584 -13 589 -5
rect 723 -7 730 -5
rect 584 -15 591 -13
rect 633 -10 640 -8
rect 584 -17 587 -15
rect 589 -17 591 -15
rect 584 -19 591 -17
rect 603 -17 610 -14
rect 603 -19 605 -17
rect 607 -19 610 -17
rect 566 -21 573 -19
rect 603 -21 610 -19
rect 612 -15 618 -14
rect 633 -12 635 -10
rect 637 -12 640 -10
rect 633 -14 640 -12
rect 642 -14 647 -8
rect 649 -10 657 -8
rect 649 -12 652 -10
rect 654 -12 657 -10
rect 649 -14 657 -12
rect 659 -14 664 -8
rect 666 -10 674 -8
rect 666 -12 669 -10
rect 671 -12 674 -10
rect 666 -14 674 -12
rect 676 -10 684 -8
rect 676 -12 679 -10
rect 681 -12 684 -10
rect 676 -14 684 -12
rect 686 -10 694 -8
rect 686 -12 689 -10
rect 691 -12 694 -10
rect 686 -14 694 -12
rect 696 -14 701 -8
rect 703 -10 710 -8
rect 723 -9 725 -7
rect 727 -9 730 -7
rect 703 -12 706 -10
rect 708 -12 710 -10
rect 703 -14 710 -12
rect 723 -11 730 -9
rect 612 -17 620 -15
rect 612 -19 615 -17
rect 617 -19 620 -17
rect 612 -21 620 -19
rect 622 -17 629 -15
rect 622 -19 625 -17
rect 627 -19 629 -17
rect 622 -21 629 -19
rect 705 -21 712 -14
rect 714 -15 719 -14
rect 714 -17 721 -15
rect 714 -19 717 -17
rect 719 -19 721 -17
rect 725 -19 730 -11
rect 732 -13 737 -5
rect 871 -7 878 -5
rect 732 -15 739 -13
rect 781 -10 788 -8
rect 732 -17 735 -15
rect 737 -17 739 -15
rect 732 -19 739 -17
rect 751 -17 758 -14
rect 751 -19 753 -17
rect 755 -19 758 -17
rect 714 -21 721 -19
rect 751 -21 758 -19
rect 760 -15 766 -14
rect 781 -12 783 -10
rect 785 -12 788 -10
rect 781 -14 788 -12
rect 790 -14 795 -8
rect 797 -10 805 -8
rect 797 -12 800 -10
rect 802 -12 805 -10
rect 797 -14 805 -12
rect 807 -14 812 -8
rect 814 -10 822 -8
rect 814 -12 817 -10
rect 819 -12 822 -10
rect 814 -14 822 -12
rect 824 -10 832 -8
rect 824 -12 827 -10
rect 829 -12 832 -10
rect 824 -14 832 -12
rect 834 -10 842 -8
rect 834 -12 837 -10
rect 839 -12 842 -10
rect 834 -14 842 -12
rect 844 -14 849 -8
rect 851 -10 858 -8
rect 871 -9 873 -7
rect 875 -9 878 -7
rect 851 -12 854 -10
rect 856 -12 858 -10
rect 851 -14 858 -12
rect 871 -11 878 -9
rect 760 -17 768 -15
rect 760 -19 763 -17
rect 765 -19 768 -17
rect 760 -21 768 -19
rect 770 -17 777 -15
rect 770 -19 773 -17
rect 775 -19 777 -17
rect 770 -21 777 -19
rect 853 -21 860 -14
rect 862 -15 867 -14
rect 862 -17 869 -15
rect 862 -19 865 -17
rect 867 -19 869 -17
rect 873 -19 878 -11
rect 880 -13 885 -5
rect 1019 -7 1026 -5
rect 880 -15 887 -13
rect 929 -10 936 -8
rect 880 -17 883 -15
rect 885 -17 887 -15
rect 880 -19 887 -17
rect 899 -17 906 -14
rect 899 -19 901 -17
rect 903 -19 906 -17
rect 862 -21 869 -19
rect 899 -21 906 -19
rect 908 -15 914 -14
rect 929 -12 931 -10
rect 933 -12 936 -10
rect 929 -14 936 -12
rect 938 -14 943 -8
rect 945 -10 953 -8
rect 945 -12 948 -10
rect 950 -12 953 -10
rect 945 -14 953 -12
rect 955 -14 960 -8
rect 962 -10 970 -8
rect 962 -12 965 -10
rect 967 -12 970 -10
rect 962 -14 970 -12
rect 972 -10 980 -8
rect 972 -12 975 -10
rect 977 -12 980 -10
rect 972 -14 980 -12
rect 982 -10 990 -8
rect 982 -12 985 -10
rect 987 -12 990 -10
rect 982 -14 990 -12
rect 992 -14 997 -8
rect 999 -10 1006 -8
rect 1019 -9 1021 -7
rect 1023 -9 1026 -7
rect 999 -12 1002 -10
rect 1004 -12 1006 -10
rect 999 -14 1006 -12
rect 1019 -11 1026 -9
rect 908 -17 916 -15
rect 908 -19 911 -17
rect 913 -19 916 -17
rect 908 -21 916 -19
rect 918 -17 925 -15
rect 918 -19 921 -17
rect 923 -19 925 -17
rect 918 -21 925 -19
rect 1001 -21 1008 -14
rect 1010 -15 1015 -14
rect 1010 -17 1017 -15
rect 1010 -19 1013 -17
rect 1015 -19 1017 -17
rect 1021 -19 1026 -11
rect 1028 -13 1033 -5
rect 1167 -7 1174 -5
rect 1028 -15 1035 -13
rect 1077 -10 1084 -8
rect 1028 -17 1031 -15
rect 1033 -17 1035 -15
rect 1028 -19 1035 -17
rect 1047 -17 1054 -14
rect 1047 -19 1049 -17
rect 1051 -19 1054 -17
rect 1010 -21 1017 -19
rect 1047 -21 1054 -19
rect 1056 -15 1062 -14
rect 1077 -12 1079 -10
rect 1081 -12 1084 -10
rect 1077 -14 1084 -12
rect 1086 -14 1091 -8
rect 1093 -10 1101 -8
rect 1093 -12 1096 -10
rect 1098 -12 1101 -10
rect 1093 -14 1101 -12
rect 1103 -14 1108 -8
rect 1110 -10 1118 -8
rect 1110 -12 1113 -10
rect 1115 -12 1118 -10
rect 1110 -14 1118 -12
rect 1120 -10 1128 -8
rect 1120 -12 1123 -10
rect 1125 -12 1128 -10
rect 1120 -14 1128 -12
rect 1130 -10 1138 -8
rect 1130 -12 1133 -10
rect 1135 -12 1138 -10
rect 1130 -14 1138 -12
rect 1140 -14 1145 -8
rect 1147 -10 1154 -8
rect 1167 -9 1169 -7
rect 1171 -9 1174 -7
rect 1147 -12 1150 -10
rect 1152 -12 1154 -10
rect 1147 -14 1154 -12
rect 1167 -11 1174 -9
rect 1056 -17 1064 -15
rect 1056 -19 1059 -17
rect 1061 -19 1064 -17
rect 1056 -21 1064 -19
rect 1066 -17 1073 -15
rect 1066 -19 1069 -17
rect 1071 -19 1073 -17
rect 1066 -21 1073 -19
rect 1149 -21 1156 -14
rect 1158 -15 1163 -14
rect 1158 -17 1165 -15
rect 1158 -19 1161 -17
rect 1163 -19 1165 -17
rect 1169 -19 1174 -11
rect 1176 -13 1181 -5
rect 1176 -15 1183 -13
rect 1176 -17 1179 -15
rect 1181 -17 1183 -15
rect 1176 -19 1183 -17
rect 1158 -21 1165 -19
rect 126 -115 133 -113
rect 126 -117 128 -115
rect 130 -117 133 -115
rect 126 -119 133 -117
rect 128 -122 133 -119
rect 135 -118 146 -113
rect 135 -120 142 -118
rect 144 -120 146 -118
rect 135 -122 146 -120
<< pdif >>
rect 9 57 14 71
rect 7 54 14 57
rect 7 52 9 54
rect 11 52 14 54
rect 7 47 14 52
rect 7 45 9 47
rect 11 45 14 47
rect 7 43 14 45
rect 16 69 23 71
rect 16 67 19 69
rect 21 67 23 69
rect 16 65 23 67
rect 16 57 22 65
rect 55 59 60 65
rect 35 57 43 59
rect 16 55 24 57
rect 16 53 19 55
rect 21 53 24 55
rect 16 43 24 53
rect 26 49 31 57
rect 35 55 37 57
rect 39 55 43 57
rect 35 53 43 55
rect 45 53 50 59
rect 52 57 60 59
rect 52 55 55 57
rect 57 55 60 57
rect 52 53 60 55
rect 62 57 70 65
rect 62 55 65 57
rect 67 55 70 57
rect 62 53 70 55
rect 72 63 80 65
rect 72 61 75 63
rect 77 61 80 63
rect 72 59 80 61
rect 82 59 87 65
rect 89 63 97 65
rect 89 61 92 63
rect 94 61 97 63
rect 89 59 97 61
rect 72 53 78 59
rect 26 47 33 49
rect 26 45 29 47
rect 31 45 33 47
rect 26 43 33 45
rect 92 52 97 59
rect 99 52 104 65
rect 106 63 111 65
rect 106 61 114 63
rect 106 59 109 61
rect 111 59 114 61
rect 106 52 114 59
rect 116 58 121 63
rect 127 62 134 64
rect 127 60 129 62
rect 131 60 134 62
rect 116 56 123 58
rect 116 54 119 56
rect 121 54 123 56
rect 127 54 134 60
rect 136 60 141 64
rect 136 58 143 60
rect 136 56 139 58
rect 141 56 143 58
rect 157 57 162 71
rect 136 54 143 56
rect 155 54 162 57
rect 116 52 123 54
rect 155 52 157 54
rect 159 52 162 54
rect 155 47 162 52
rect 155 45 157 47
rect 159 45 162 47
rect 155 43 162 45
rect 164 69 171 71
rect 164 67 167 69
rect 169 67 171 69
rect 164 65 171 67
rect 164 57 170 65
rect 203 59 208 65
rect 183 57 191 59
rect 164 55 172 57
rect 164 53 167 55
rect 169 53 172 55
rect 164 43 172 53
rect 174 49 179 57
rect 183 55 185 57
rect 187 55 191 57
rect 183 53 191 55
rect 193 53 198 59
rect 200 57 208 59
rect 200 55 203 57
rect 205 55 208 57
rect 200 53 208 55
rect 210 57 218 65
rect 210 55 213 57
rect 215 55 218 57
rect 210 53 218 55
rect 220 63 228 65
rect 220 61 223 63
rect 225 61 228 63
rect 220 59 228 61
rect 230 59 235 65
rect 237 63 245 65
rect 237 61 240 63
rect 242 61 245 63
rect 237 59 245 61
rect 220 53 226 59
rect 174 47 181 49
rect 174 45 177 47
rect 179 45 181 47
rect 174 43 181 45
rect 240 52 245 59
rect 247 52 252 65
rect 254 63 259 65
rect 254 61 262 63
rect 254 59 257 61
rect 259 59 262 61
rect 254 52 262 59
rect 264 58 269 63
rect 275 62 282 64
rect 275 60 277 62
rect 279 60 282 62
rect 264 56 271 58
rect 264 54 267 56
rect 269 54 271 56
rect 275 54 282 60
rect 284 60 289 64
rect 284 58 291 60
rect 284 56 287 58
rect 289 56 291 58
rect 305 57 310 71
rect 284 54 291 56
rect 303 54 310 57
rect 264 52 271 54
rect 303 52 305 54
rect 307 52 310 54
rect 303 47 310 52
rect 303 45 305 47
rect 307 45 310 47
rect 303 43 310 45
rect 312 69 319 71
rect 312 67 315 69
rect 317 67 319 69
rect 312 65 319 67
rect 312 57 318 65
rect 351 59 356 65
rect 331 57 339 59
rect 312 55 320 57
rect 312 53 315 55
rect 317 53 320 55
rect 312 43 320 53
rect 322 49 327 57
rect 331 55 333 57
rect 335 55 339 57
rect 331 53 339 55
rect 341 53 346 59
rect 348 57 356 59
rect 348 55 351 57
rect 353 55 356 57
rect 348 53 356 55
rect 358 57 366 65
rect 358 55 361 57
rect 363 55 366 57
rect 358 53 366 55
rect 368 63 376 65
rect 368 61 371 63
rect 373 61 376 63
rect 368 59 376 61
rect 378 59 383 65
rect 385 63 393 65
rect 385 61 388 63
rect 390 61 393 63
rect 385 59 393 61
rect 368 53 374 59
rect 322 47 329 49
rect 322 45 325 47
rect 327 45 329 47
rect 322 43 329 45
rect 388 52 393 59
rect 395 52 400 65
rect 402 63 407 65
rect 402 61 410 63
rect 402 59 405 61
rect 407 59 410 61
rect 402 52 410 59
rect 412 58 417 63
rect 423 62 430 64
rect 423 60 425 62
rect 427 60 430 62
rect 412 56 419 58
rect 412 54 415 56
rect 417 54 419 56
rect 423 54 430 60
rect 432 60 437 64
rect 432 58 439 60
rect 432 56 435 58
rect 437 56 439 58
rect 453 57 458 71
rect 432 54 439 56
rect 451 54 458 57
rect 412 52 419 54
rect 451 52 453 54
rect 455 52 458 54
rect 451 47 458 52
rect 451 45 453 47
rect 455 45 458 47
rect 451 43 458 45
rect 460 69 467 71
rect 460 67 463 69
rect 465 67 467 69
rect 460 65 467 67
rect 460 57 466 65
rect 499 59 504 65
rect 479 57 487 59
rect 460 55 468 57
rect 460 53 463 55
rect 465 53 468 55
rect 460 43 468 53
rect 470 49 475 57
rect 479 55 481 57
rect 483 55 487 57
rect 479 53 487 55
rect 489 53 494 59
rect 496 57 504 59
rect 496 55 499 57
rect 501 55 504 57
rect 496 53 504 55
rect 506 57 514 65
rect 506 55 509 57
rect 511 55 514 57
rect 506 53 514 55
rect 516 63 524 65
rect 516 61 519 63
rect 521 61 524 63
rect 516 59 524 61
rect 526 59 531 65
rect 533 63 541 65
rect 533 61 536 63
rect 538 61 541 63
rect 533 59 541 61
rect 516 53 522 59
rect 470 47 477 49
rect 470 45 473 47
rect 475 45 477 47
rect 470 43 477 45
rect 536 52 541 59
rect 543 52 548 65
rect 550 63 555 65
rect 550 61 558 63
rect 550 59 553 61
rect 555 59 558 61
rect 550 52 558 59
rect 560 58 565 63
rect 571 62 578 64
rect 571 60 573 62
rect 575 60 578 62
rect 560 56 567 58
rect 560 54 563 56
rect 565 54 567 56
rect 571 54 578 60
rect 580 60 585 64
rect 580 58 587 60
rect 580 56 583 58
rect 585 56 587 58
rect 601 57 606 71
rect 580 54 587 56
rect 599 54 606 57
rect 560 52 567 54
rect 599 52 601 54
rect 603 52 606 54
rect 599 47 606 52
rect 599 45 601 47
rect 603 45 606 47
rect 599 43 606 45
rect 608 69 615 71
rect 608 67 611 69
rect 613 67 615 69
rect 608 65 615 67
rect 608 57 614 65
rect 647 59 652 65
rect 627 57 635 59
rect 608 55 616 57
rect 608 53 611 55
rect 613 53 616 55
rect 608 43 616 53
rect 618 49 623 57
rect 627 55 629 57
rect 631 55 635 57
rect 627 53 635 55
rect 637 53 642 59
rect 644 57 652 59
rect 644 55 647 57
rect 649 55 652 57
rect 644 53 652 55
rect 654 57 662 65
rect 654 55 657 57
rect 659 55 662 57
rect 654 53 662 55
rect 664 63 672 65
rect 664 61 667 63
rect 669 61 672 63
rect 664 59 672 61
rect 674 59 679 65
rect 681 63 689 65
rect 681 61 684 63
rect 686 61 689 63
rect 681 59 689 61
rect 664 53 670 59
rect 618 47 625 49
rect 618 45 621 47
rect 623 45 625 47
rect 618 43 625 45
rect 684 52 689 59
rect 691 52 696 65
rect 698 63 703 65
rect 698 61 706 63
rect 698 59 701 61
rect 703 59 706 61
rect 698 52 706 59
rect 708 58 713 63
rect 719 62 726 64
rect 719 60 721 62
rect 723 60 726 62
rect 708 56 715 58
rect 708 54 711 56
rect 713 54 715 56
rect 719 54 726 60
rect 728 60 733 64
rect 728 58 735 60
rect 728 56 731 58
rect 733 56 735 58
rect 749 57 754 71
rect 728 54 735 56
rect 747 54 754 57
rect 708 52 715 54
rect 747 52 749 54
rect 751 52 754 54
rect 747 47 754 52
rect 747 45 749 47
rect 751 45 754 47
rect 747 43 754 45
rect 756 69 763 71
rect 756 67 759 69
rect 761 67 763 69
rect 756 65 763 67
rect 756 57 762 65
rect 795 59 800 65
rect 775 57 783 59
rect 756 55 764 57
rect 756 53 759 55
rect 761 53 764 55
rect 756 43 764 53
rect 766 49 771 57
rect 775 55 777 57
rect 779 55 783 57
rect 775 53 783 55
rect 785 53 790 59
rect 792 57 800 59
rect 792 55 795 57
rect 797 55 800 57
rect 792 53 800 55
rect 802 57 810 65
rect 802 55 805 57
rect 807 55 810 57
rect 802 53 810 55
rect 812 63 820 65
rect 812 61 815 63
rect 817 61 820 63
rect 812 59 820 61
rect 822 59 827 65
rect 829 63 837 65
rect 829 61 832 63
rect 834 61 837 63
rect 829 59 837 61
rect 812 53 818 59
rect 766 47 773 49
rect 766 45 769 47
rect 771 45 773 47
rect 766 43 773 45
rect 832 52 837 59
rect 839 52 844 65
rect 846 63 851 65
rect 846 61 854 63
rect 846 59 849 61
rect 851 59 854 61
rect 846 52 854 59
rect 856 58 861 63
rect 867 62 874 64
rect 867 60 869 62
rect 871 60 874 62
rect 856 56 863 58
rect 856 54 859 56
rect 861 54 863 56
rect 867 54 874 60
rect 876 60 881 64
rect 876 58 883 60
rect 876 56 879 58
rect 881 56 883 58
rect 897 57 902 71
rect 876 54 883 56
rect 895 54 902 57
rect 856 52 863 54
rect 895 52 897 54
rect 899 52 902 54
rect 895 47 902 52
rect 895 45 897 47
rect 899 45 902 47
rect 895 43 902 45
rect 904 69 911 71
rect 904 67 907 69
rect 909 67 911 69
rect 904 65 911 67
rect 904 57 910 65
rect 943 59 948 65
rect 923 57 931 59
rect 904 55 912 57
rect 904 53 907 55
rect 909 53 912 55
rect 904 43 912 53
rect 914 49 919 57
rect 923 55 925 57
rect 927 55 931 57
rect 923 53 931 55
rect 933 53 938 59
rect 940 57 948 59
rect 940 55 943 57
rect 945 55 948 57
rect 940 53 948 55
rect 950 57 958 65
rect 950 55 953 57
rect 955 55 958 57
rect 950 53 958 55
rect 960 63 968 65
rect 960 61 963 63
rect 965 61 968 63
rect 960 59 968 61
rect 970 59 975 65
rect 977 63 985 65
rect 977 61 980 63
rect 982 61 985 63
rect 977 59 985 61
rect 960 53 966 59
rect 914 47 921 49
rect 914 45 917 47
rect 919 45 921 47
rect 914 43 921 45
rect 980 52 985 59
rect 987 52 992 65
rect 994 63 999 65
rect 994 61 1002 63
rect 994 59 997 61
rect 999 59 1002 61
rect 994 52 1002 59
rect 1004 58 1009 63
rect 1015 62 1022 64
rect 1015 60 1017 62
rect 1019 60 1022 62
rect 1004 56 1011 58
rect 1004 54 1007 56
rect 1009 54 1011 56
rect 1015 54 1022 60
rect 1024 60 1029 64
rect 1024 58 1031 60
rect 1024 56 1027 58
rect 1029 56 1031 58
rect 1045 57 1050 71
rect 1024 54 1031 56
rect 1043 54 1050 57
rect 1004 52 1011 54
rect 1043 52 1045 54
rect 1047 52 1050 54
rect 1043 47 1050 52
rect 1043 45 1045 47
rect 1047 45 1050 47
rect 1043 43 1050 45
rect 1052 69 1059 71
rect 1052 67 1055 69
rect 1057 67 1059 69
rect 1052 65 1059 67
rect 1052 57 1058 65
rect 1091 59 1096 65
rect 1071 57 1079 59
rect 1052 55 1060 57
rect 1052 53 1055 55
rect 1057 53 1060 55
rect 1052 43 1060 53
rect 1062 49 1067 57
rect 1071 55 1073 57
rect 1075 55 1079 57
rect 1071 53 1079 55
rect 1081 53 1086 59
rect 1088 57 1096 59
rect 1088 55 1091 57
rect 1093 55 1096 57
rect 1088 53 1096 55
rect 1098 57 1106 65
rect 1098 55 1101 57
rect 1103 55 1106 57
rect 1098 53 1106 55
rect 1108 63 1116 65
rect 1108 61 1111 63
rect 1113 61 1116 63
rect 1108 59 1116 61
rect 1118 59 1123 65
rect 1125 63 1133 65
rect 1125 61 1128 63
rect 1130 61 1133 63
rect 1125 59 1133 61
rect 1108 53 1114 59
rect 1062 47 1069 49
rect 1062 45 1065 47
rect 1067 45 1069 47
rect 1062 43 1069 45
rect 1128 52 1133 59
rect 1135 52 1140 65
rect 1142 63 1147 65
rect 1142 61 1150 63
rect 1142 59 1145 61
rect 1147 59 1150 61
rect 1142 52 1150 59
rect 1152 58 1157 63
rect 1163 62 1170 64
rect 1163 60 1165 62
rect 1167 60 1170 62
rect 1152 56 1159 58
rect 1152 54 1155 56
rect 1157 54 1159 56
rect 1163 54 1170 60
rect 1172 60 1177 64
rect 1172 58 1179 60
rect 1172 56 1175 58
rect 1177 56 1179 58
rect 1172 54 1179 56
rect 1152 52 1159 54
rect 31 -44 38 -42
rect 11 -46 18 -44
rect 11 -48 13 -46
rect 15 -48 18 -46
rect 11 -50 18 -48
rect 13 -54 18 -50
rect 20 -50 27 -44
rect 31 -46 33 -44
rect 35 -46 38 -44
rect 31 -48 38 -46
rect 20 -52 23 -50
rect 25 -52 27 -50
rect 20 -54 27 -52
rect 33 -53 38 -48
rect 40 -49 48 -42
rect 40 -51 43 -49
rect 45 -51 48 -49
rect 40 -53 48 -51
rect 43 -55 48 -53
rect 50 -55 55 -42
rect 57 -49 62 -42
rect 121 -35 128 -33
rect 121 -37 123 -35
rect 125 -37 128 -35
rect 121 -39 128 -37
rect 76 -49 82 -43
rect 57 -51 65 -49
rect 57 -53 60 -51
rect 62 -53 65 -51
rect 57 -55 65 -53
rect 67 -55 72 -49
rect 74 -51 82 -49
rect 74 -53 77 -51
rect 79 -53 82 -51
rect 74 -55 82 -53
rect 84 -45 92 -43
rect 84 -47 87 -45
rect 89 -47 92 -45
rect 84 -55 92 -47
rect 94 -45 102 -43
rect 94 -47 97 -45
rect 99 -47 102 -45
rect 94 -49 102 -47
rect 104 -49 109 -43
rect 111 -45 119 -43
rect 111 -47 115 -45
rect 117 -47 119 -45
rect 123 -47 128 -39
rect 130 -43 138 -33
rect 130 -45 133 -43
rect 135 -45 138 -43
rect 130 -47 138 -45
rect 111 -49 119 -47
rect 94 -55 99 -49
rect 132 -55 138 -47
rect 131 -57 138 -55
rect 131 -59 133 -57
rect 135 -59 138 -57
rect 131 -61 138 -59
rect 140 -35 147 -33
rect 140 -37 143 -35
rect 145 -37 147 -35
rect 140 -42 147 -37
rect 140 -44 143 -42
rect 145 -44 147 -42
rect 179 -44 186 -42
rect 140 -47 147 -44
rect 159 -46 166 -44
rect 140 -61 145 -47
rect 159 -48 161 -46
rect 163 -48 166 -46
rect 159 -50 166 -48
rect 161 -54 166 -50
rect 168 -50 175 -44
rect 179 -46 181 -44
rect 183 -46 186 -44
rect 179 -48 186 -46
rect 168 -52 171 -50
rect 173 -52 175 -50
rect 168 -54 175 -52
rect 181 -53 186 -48
rect 188 -49 196 -42
rect 188 -51 191 -49
rect 193 -51 196 -49
rect 188 -53 196 -51
rect 191 -55 196 -53
rect 198 -55 203 -42
rect 205 -49 210 -42
rect 269 -35 276 -33
rect 269 -37 271 -35
rect 273 -37 276 -35
rect 269 -39 276 -37
rect 224 -49 230 -43
rect 205 -51 213 -49
rect 205 -53 208 -51
rect 210 -53 213 -51
rect 205 -55 213 -53
rect 215 -55 220 -49
rect 222 -51 230 -49
rect 222 -53 225 -51
rect 227 -53 230 -51
rect 222 -55 230 -53
rect 232 -45 240 -43
rect 232 -47 235 -45
rect 237 -47 240 -45
rect 232 -55 240 -47
rect 242 -45 250 -43
rect 242 -47 245 -45
rect 247 -47 250 -45
rect 242 -49 250 -47
rect 252 -49 257 -43
rect 259 -45 267 -43
rect 259 -47 263 -45
rect 265 -47 267 -45
rect 271 -47 276 -39
rect 278 -43 286 -33
rect 278 -45 281 -43
rect 283 -45 286 -43
rect 278 -47 286 -45
rect 259 -49 267 -47
rect 242 -55 247 -49
rect 280 -55 286 -47
rect 279 -57 286 -55
rect 279 -59 281 -57
rect 283 -59 286 -57
rect 279 -61 286 -59
rect 288 -35 295 -33
rect 288 -37 291 -35
rect 293 -37 295 -35
rect 288 -42 295 -37
rect 288 -44 291 -42
rect 293 -44 295 -42
rect 327 -44 334 -42
rect 288 -47 295 -44
rect 307 -46 314 -44
rect 288 -61 293 -47
rect 307 -48 309 -46
rect 311 -48 314 -46
rect 307 -50 314 -48
rect 309 -54 314 -50
rect 316 -50 323 -44
rect 327 -46 329 -44
rect 331 -46 334 -44
rect 327 -48 334 -46
rect 316 -52 319 -50
rect 321 -52 323 -50
rect 316 -54 323 -52
rect 329 -53 334 -48
rect 336 -49 344 -42
rect 336 -51 339 -49
rect 341 -51 344 -49
rect 336 -53 344 -51
rect 339 -55 344 -53
rect 346 -55 351 -42
rect 353 -49 358 -42
rect 417 -35 424 -33
rect 417 -37 419 -35
rect 421 -37 424 -35
rect 417 -39 424 -37
rect 372 -49 378 -43
rect 353 -51 361 -49
rect 353 -53 356 -51
rect 358 -53 361 -51
rect 353 -55 361 -53
rect 363 -55 368 -49
rect 370 -51 378 -49
rect 370 -53 373 -51
rect 375 -53 378 -51
rect 370 -55 378 -53
rect 380 -45 388 -43
rect 380 -47 383 -45
rect 385 -47 388 -45
rect 380 -55 388 -47
rect 390 -45 398 -43
rect 390 -47 393 -45
rect 395 -47 398 -45
rect 390 -49 398 -47
rect 400 -49 405 -43
rect 407 -45 415 -43
rect 407 -47 411 -45
rect 413 -47 415 -45
rect 419 -47 424 -39
rect 426 -43 434 -33
rect 426 -45 429 -43
rect 431 -45 434 -43
rect 426 -47 434 -45
rect 407 -49 415 -47
rect 390 -55 395 -49
rect 428 -55 434 -47
rect 427 -57 434 -55
rect 427 -59 429 -57
rect 431 -59 434 -57
rect 427 -61 434 -59
rect 436 -35 443 -33
rect 436 -37 439 -35
rect 441 -37 443 -35
rect 436 -42 443 -37
rect 436 -44 439 -42
rect 441 -44 443 -42
rect 475 -44 482 -42
rect 436 -47 443 -44
rect 455 -46 462 -44
rect 436 -61 441 -47
rect 455 -48 457 -46
rect 459 -48 462 -46
rect 455 -50 462 -48
rect 457 -54 462 -50
rect 464 -50 471 -44
rect 475 -46 477 -44
rect 479 -46 482 -44
rect 475 -48 482 -46
rect 464 -52 467 -50
rect 469 -52 471 -50
rect 464 -54 471 -52
rect 477 -53 482 -48
rect 484 -49 492 -42
rect 484 -51 487 -49
rect 489 -51 492 -49
rect 484 -53 492 -51
rect 487 -55 492 -53
rect 494 -55 499 -42
rect 501 -49 506 -42
rect 565 -35 572 -33
rect 565 -37 567 -35
rect 569 -37 572 -35
rect 565 -39 572 -37
rect 520 -49 526 -43
rect 501 -51 509 -49
rect 501 -53 504 -51
rect 506 -53 509 -51
rect 501 -55 509 -53
rect 511 -55 516 -49
rect 518 -51 526 -49
rect 518 -53 521 -51
rect 523 -53 526 -51
rect 518 -55 526 -53
rect 528 -45 536 -43
rect 528 -47 531 -45
rect 533 -47 536 -45
rect 528 -55 536 -47
rect 538 -45 546 -43
rect 538 -47 541 -45
rect 543 -47 546 -45
rect 538 -49 546 -47
rect 548 -49 553 -43
rect 555 -45 563 -43
rect 555 -47 559 -45
rect 561 -47 563 -45
rect 567 -47 572 -39
rect 574 -43 582 -33
rect 574 -45 577 -43
rect 579 -45 582 -43
rect 574 -47 582 -45
rect 555 -49 563 -47
rect 538 -55 543 -49
rect 576 -55 582 -47
rect 575 -57 582 -55
rect 575 -59 577 -57
rect 579 -59 582 -57
rect 575 -61 582 -59
rect 584 -35 591 -33
rect 584 -37 587 -35
rect 589 -37 591 -35
rect 584 -42 591 -37
rect 584 -44 587 -42
rect 589 -44 591 -42
rect 623 -44 630 -42
rect 584 -47 591 -44
rect 603 -46 610 -44
rect 584 -61 589 -47
rect 603 -48 605 -46
rect 607 -48 610 -46
rect 603 -50 610 -48
rect 605 -54 610 -50
rect 612 -50 619 -44
rect 623 -46 625 -44
rect 627 -46 630 -44
rect 623 -48 630 -46
rect 612 -52 615 -50
rect 617 -52 619 -50
rect 612 -54 619 -52
rect 625 -53 630 -48
rect 632 -49 640 -42
rect 632 -51 635 -49
rect 637 -51 640 -49
rect 632 -53 640 -51
rect 635 -55 640 -53
rect 642 -55 647 -42
rect 649 -49 654 -42
rect 713 -35 720 -33
rect 713 -37 715 -35
rect 717 -37 720 -35
rect 713 -39 720 -37
rect 668 -49 674 -43
rect 649 -51 657 -49
rect 649 -53 652 -51
rect 654 -53 657 -51
rect 649 -55 657 -53
rect 659 -55 664 -49
rect 666 -51 674 -49
rect 666 -53 669 -51
rect 671 -53 674 -51
rect 666 -55 674 -53
rect 676 -45 684 -43
rect 676 -47 679 -45
rect 681 -47 684 -45
rect 676 -55 684 -47
rect 686 -45 694 -43
rect 686 -47 689 -45
rect 691 -47 694 -45
rect 686 -49 694 -47
rect 696 -49 701 -43
rect 703 -45 711 -43
rect 703 -47 707 -45
rect 709 -47 711 -45
rect 715 -47 720 -39
rect 722 -43 730 -33
rect 722 -45 725 -43
rect 727 -45 730 -43
rect 722 -47 730 -45
rect 703 -49 711 -47
rect 686 -55 691 -49
rect 724 -55 730 -47
rect 723 -57 730 -55
rect 723 -59 725 -57
rect 727 -59 730 -57
rect 723 -61 730 -59
rect 732 -35 739 -33
rect 732 -37 735 -35
rect 737 -37 739 -35
rect 732 -42 739 -37
rect 732 -44 735 -42
rect 737 -44 739 -42
rect 771 -44 778 -42
rect 732 -47 739 -44
rect 751 -46 758 -44
rect 732 -61 737 -47
rect 751 -48 753 -46
rect 755 -48 758 -46
rect 751 -50 758 -48
rect 753 -54 758 -50
rect 760 -50 767 -44
rect 771 -46 773 -44
rect 775 -46 778 -44
rect 771 -48 778 -46
rect 760 -52 763 -50
rect 765 -52 767 -50
rect 760 -54 767 -52
rect 773 -53 778 -48
rect 780 -49 788 -42
rect 780 -51 783 -49
rect 785 -51 788 -49
rect 780 -53 788 -51
rect 783 -55 788 -53
rect 790 -55 795 -42
rect 797 -49 802 -42
rect 861 -35 868 -33
rect 861 -37 863 -35
rect 865 -37 868 -35
rect 861 -39 868 -37
rect 816 -49 822 -43
rect 797 -51 805 -49
rect 797 -53 800 -51
rect 802 -53 805 -51
rect 797 -55 805 -53
rect 807 -55 812 -49
rect 814 -51 822 -49
rect 814 -53 817 -51
rect 819 -53 822 -51
rect 814 -55 822 -53
rect 824 -45 832 -43
rect 824 -47 827 -45
rect 829 -47 832 -45
rect 824 -55 832 -47
rect 834 -45 842 -43
rect 834 -47 837 -45
rect 839 -47 842 -45
rect 834 -49 842 -47
rect 844 -49 849 -43
rect 851 -45 859 -43
rect 851 -47 855 -45
rect 857 -47 859 -45
rect 863 -47 868 -39
rect 870 -43 878 -33
rect 870 -45 873 -43
rect 875 -45 878 -43
rect 870 -47 878 -45
rect 851 -49 859 -47
rect 834 -55 839 -49
rect 872 -55 878 -47
rect 871 -57 878 -55
rect 871 -59 873 -57
rect 875 -59 878 -57
rect 871 -61 878 -59
rect 880 -35 887 -33
rect 880 -37 883 -35
rect 885 -37 887 -35
rect 880 -42 887 -37
rect 880 -44 883 -42
rect 885 -44 887 -42
rect 919 -44 926 -42
rect 880 -47 887 -44
rect 899 -46 906 -44
rect 880 -61 885 -47
rect 899 -48 901 -46
rect 903 -48 906 -46
rect 899 -50 906 -48
rect 901 -54 906 -50
rect 908 -50 915 -44
rect 919 -46 921 -44
rect 923 -46 926 -44
rect 919 -48 926 -46
rect 908 -52 911 -50
rect 913 -52 915 -50
rect 908 -54 915 -52
rect 921 -53 926 -48
rect 928 -49 936 -42
rect 928 -51 931 -49
rect 933 -51 936 -49
rect 928 -53 936 -51
rect 931 -55 936 -53
rect 938 -55 943 -42
rect 945 -49 950 -42
rect 1009 -35 1016 -33
rect 1009 -37 1011 -35
rect 1013 -37 1016 -35
rect 1009 -39 1016 -37
rect 964 -49 970 -43
rect 945 -51 953 -49
rect 945 -53 948 -51
rect 950 -53 953 -51
rect 945 -55 953 -53
rect 955 -55 960 -49
rect 962 -51 970 -49
rect 962 -53 965 -51
rect 967 -53 970 -51
rect 962 -55 970 -53
rect 972 -45 980 -43
rect 972 -47 975 -45
rect 977 -47 980 -45
rect 972 -55 980 -47
rect 982 -45 990 -43
rect 982 -47 985 -45
rect 987 -47 990 -45
rect 982 -49 990 -47
rect 992 -49 997 -43
rect 999 -45 1007 -43
rect 999 -47 1003 -45
rect 1005 -47 1007 -45
rect 1011 -47 1016 -39
rect 1018 -43 1026 -33
rect 1018 -45 1021 -43
rect 1023 -45 1026 -43
rect 1018 -47 1026 -45
rect 999 -49 1007 -47
rect 982 -55 987 -49
rect 1020 -55 1026 -47
rect 1019 -57 1026 -55
rect 1019 -59 1021 -57
rect 1023 -59 1026 -57
rect 1019 -61 1026 -59
rect 1028 -35 1035 -33
rect 1028 -37 1031 -35
rect 1033 -37 1035 -35
rect 1028 -42 1035 -37
rect 1028 -44 1031 -42
rect 1033 -44 1035 -42
rect 1067 -44 1074 -42
rect 1028 -47 1035 -44
rect 1047 -46 1054 -44
rect 1028 -61 1033 -47
rect 1047 -48 1049 -46
rect 1051 -48 1054 -46
rect 1047 -50 1054 -48
rect 1049 -54 1054 -50
rect 1056 -50 1063 -44
rect 1067 -46 1069 -44
rect 1071 -46 1074 -44
rect 1067 -48 1074 -46
rect 1056 -52 1059 -50
rect 1061 -52 1063 -50
rect 1056 -54 1063 -52
rect 1069 -53 1074 -48
rect 1076 -49 1084 -42
rect 1076 -51 1079 -49
rect 1081 -51 1084 -49
rect 1076 -53 1084 -51
rect 1079 -55 1084 -53
rect 1086 -55 1091 -42
rect 1093 -49 1098 -42
rect 1157 -35 1164 -33
rect 1157 -37 1159 -35
rect 1161 -37 1164 -35
rect 1157 -39 1164 -37
rect 1112 -49 1118 -43
rect 1093 -51 1101 -49
rect 1093 -53 1096 -51
rect 1098 -53 1101 -51
rect 1093 -55 1101 -53
rect 1103 -55 1108 -49
rect 1110 -51 1118 -49
rect 1110 -53 1113 -51
rect 1115 -53 1118 -51
rect 1110 -55 1118 -53
rect 1120 -45 1128 -43
rect 1120 -47 1123 -45
rect 1125 -47 1128 -45
rect 1120 -55 1128 -47
rect 1130 -45 1138 -43
rect 1130 -47 1133 -45
rect 1135 -47 1138 -45
rect 1130 -49 1138 -47
rect 1140 -49 1145 -43
rect 1147 -45 1155 -43
rect 1147 -47 1151 -45
rect 1153 -47 1155 -45
rect 1159 -47 1164 -39
rect 1166 -43 1174 -33
rect 1166 -45 1169 -43
rect 1171 -45 1174 -43
rect 1166 -47 1174 -45
rect 1147 -49 1155 -47
rect 1130 -55 1135 -49
rect 1168 -55 1174 -47
rect 1167 -57 1174 -55
rect 1167 -59 1169 -57
rect 1171 -59 1174 -57
rect 1167 -61 1174 -59
rect 1176 -35 1183 -33
rect 1176 -37 1179 -35
rect 1181 -37 1183 -35
rect 1176 -42 1183 -37
rect 1176 -44 1179 -42
rect 1181 -44 1183 -42
rect 1176 -47 1183 -44
rect 1176 -61 1181 -47
rect 137 -82 144 -80
rect 137 -83 139 -82
rect 128 -88 133 -83
rect 126 -90 133 -88
rect 126 -92 128 -90
rect 130 -92 133 -90
rect 126 -97 133 -92
rect 126 -99 128 -97
rect 130 -99 133 -97
rect 126 -101 133 -99
rect 135 -84 139 -83
rect 141 -84 144 -82
rect 135 -101 144 -84
<< alu1 >>
rect 3 72 1187 77
rect 3 70 33 72
rect 35 70 43 72
rect 45 70 124 72
rect 126 70 181 72
rect 183 70 191 72
rect 193 70 272 72
rect 274 70 329 72
rect 331 70 339 72
rect 341 70 420 72
rect 422 70 477 72
rect 479 70 487 72
rect 489 70 568 72
rect 570 70 625 72
rect 627 70 635 72
rect 637 70 716 72
rect 718 70 773 72
rect 775 70 783 72
rect 785 70 864 72
rect 866 70 921 72
rect 923 70 931 72
rect 933 70 1012 72
rect 1014 70 1069 72
rect 1071 70 1079 72
rect 1081 70 1160 72
rect 1162 70 1187 72
rect 3 69 1187 70
rect 7 54 12 56
rect 7 52 9 54
rect 11 52 12 54
rect 7 47 12 52
rect 7 45 9 47
rect 11 45 20 47
rect 7 43 20 45
rect 7 29 11 43
rect 7 27 12 29
rect 7 25 9 27
rect 11 25 12 27
rect 7 23 12 25
rect 126 48 132 55
rect 126 47 129 48
rect 102 39 108 47
rect 118 46 129 47
rect 131 46 132 48
rect 118 43 132 46
rect 102 38 116 39
rect 102 36 106 38
rect 108 36 116 38
rect 102 35 116 36
rect 155 54 160 56
rect 155 52 157 54
rect 159 52 160 54
rect 155 47 160 52
rect 155 45 157 47
rect 159 45 168 47
rect 155 43 168 45
rect 155 29 159 43
rect 155 27 160 29
rect 155 25 157 27
rect 159 25 160 27
rect 155 23 160 25
rect 274 48 280 55
rect 274 47 277 48
rect 250 39 256 47
rect 266 46 277 47
rect 279 46 280 48
rect 266 43 280 46
rect 250 38 264 39
rect 250 36 254 38
rect 256 36 264 38
rect 250 35 264 36
rect 303 54 308 56
rect 303 52 305 54
rect 307 52 308 54
rect 303 47 308 52
rect 303 45 305 47
rect 307 45 316 47
rect 303 43 316 45
rect 303 29 307 43
rect 303 27 308 29
rect 303 25 305 27
rect 307 25 308 27
rect 303 23 308 25
rect 422 48 428 55
rect 422 47 425 48
rect 398 39 404 47
rect 414 46 425 47
rect 427 46 428 48
rect 414 43 428 46
rect 398 38 412 39
rect 398 36 402 38
rect 404 36 412 38
rect 398 35 412 36
rect 451 54 456 56
rect 451 52 453 54
rect 455 52 456 54
rect 451 47 456 52
rect 451 45 453 47
rect 455 45 464 47
rect 451 43 464 45
rect 451 29 455 43
rect 451 27 456 29
rect 451 25 453 27
rect 455 25 456 27
rect 451 23 456 25
rect 570 48 576 55
rect 570 47 573 48
rect 546 39 552 47
rect 562 46 573 47
rect 575 46 576 48
rect 562 43 576 46
rect 546 38 560 39
rect 546 36 550 38
rect 552 36 560 38
rect 546 35 560 36
rect 599 54 604 56
rect 599 52 601 54
rect 603 52 604 54
rect 599 47 604 52
rect 599 45 601 47
rect 603 45 612 47
rect 599 43 612 45
rect 599 29 603 43
rect 599 27 604 29
rect 599 25 601 27
rect 603 25 604 27
rect 599 23 604 25
rect 718 48 724 55
rect 718 47 721 48
rect 694 39 700 47
rect 710 46 721 47
rect 723 46 724 48
rect 710 43 724 46
rect 694 38 708 39
rect 694 36 698 38
rect 700 36 708 38
rect 694 35 708 36
rect 747 54 752 56
rect 747 52 749 54
rect 751 52 752 54
rect 747 47 752 52
rect 747 45 749 47
rect 751 45 760 47
rect 747 43 760 45
rect 747 29 751 43
rect 747 27 752 29
rect 747 25 749 27
rect 751 25 752 27
rect 747 23 752 25
rect 866 48 872 55
rect 866 47 869 48
rect 842 39 848 47
rect 858 46 869 47
rect 871 46 872 48
rect 858 43 872 46
rect 842 38 856 39
rect 842 36 846 38
rect 848 36 856 38
rect 842 35 856 36
rect 895 54 900 56
rect 895 52 897 54
rect 899 52 900 54
rect 895 47 900 52
rect 895 45 897 47
rect 899 45 908 47
rect 895 43 908 45
rect 895 29 899 43
rect 895 27 900 29
rect 895 25 897 27
rect 899 25 900 27
rect 895 23 900 25
rect 1014 48 1020 55
rect 1014 47 1017 48
rect 990 39 996 47
rect 1006 46 1017 47
rect 1019 46 1020 48
rect 1006 43 1020 46
rect 990 38 1004 39
rect 990 36 994 38
rect 996 36 1004 38
rect 990 35 1004 36
rect 1043 54 1048 56
rect 1043 52 1045 54
rect 1047 52 1048 54
rect 1043 47 1048 52
rect 1043 45 1045 47
rect 1047 45 1056 47
rect 1043 43 1056 45
rect 1043 29 1047 43
rect 1043 27 1048 29
rect 1043 25 1045 27
rect 1047 25 1048 27
rect 1043 23 1048 25
rect 1162 48 1168 55
rect 1162 47 1165 48
rect 1138 39 1144 47
rect 1154 46 1165 47
rect 1167 46 1168 48
rect 1154 43 1168 46
rect 1138 38 1152 39
rect 1138 36 1142 38
rect 1144 36 1152 38
rect 1138 35 1152 36
rect 3 12 1187 13
rect 3 10 125 12
rect 127 10 136 12
rect 138 10 273 12
rect 275 10 284 12
rect 286 10 421 12
rect 423 10 432 12
rect 434 10 569 12
rect 571 10 580 12
rect 582 10 717 12
rect 719 10 728 12
rect 730 10 865 12
rect 867 10 876 12
rect 878 10 1013 12
rect 1015 10 1024 12
rect 1026 10 1161 12
rect 1163 10 1172 12
rect 1174 10 1187 12
rect 3 0 1187 10
rect 3 -2 16 0
rect 18 -2 27 0
rect 29 -2 164 0
rect 166 -2 175 0
rect 177 -2 312 0
rect 314 -2 323 0
rect 325 -2 460 0
rect 462 -2 471 0
rect 473 -2 608 0
rect 610 -2 619 0
rect 621 -2 756 0
rect 758 -2 767 0
rect 769 -2 904 0
rect 906 -2 915 0
rect 917 -2 1052 0
rect 1054 -2 1063 0
rect 1065 -2 1187 0
rect 3 -3 1187 -2
rect 38 -26 52 -25
rect 38 -28 46 -26
rect 48 -28 52 -26
rect 38 -29 52 -28
rect 22 -36 36 -33
rect 22 -38 23 -36
rect 25 -37 36 -36
rect 46 -37 52 -29
rect 25 -38 28 -37
rect 22 -45 28 -38
rect 142 -15 147 -13
rect 142 -17 143 -15
rect 145 -17 147 -15
rect 142 -19 147 -17
rect 143 -33 147 -19
rect 134 -35 147 -33
rect 134 -37 143 -35
rect 145 -37 147 -35
rect 142 -38 147 -37
rect 142 -40 143 -38
rect 145 -40 147 -38
rect 142 -42 147 -40
rect 142 -44 143 -42
rect 145 -44 147 -42
rect 142 -46 147 -44
rect 186 -26 200 -25
rect 186 -28 194 -26
rect 196 -28 200 -26
rect 186 -29 200 -28
rect 170 -36 184 -33
rect 170 -38 171 -36
rect 173 -37 184 -36
rect 194 -37 200 -29
rect 173 -38 176 -37
rect 170 -45 176 -38
rect 290 -15 295 -13
rect 290 -17 291 -15
rect 293 -17 295 -15
rect 290 -19 295 -17
rect 291 -33 295 -19
rect 282 -35 295 -33
rect 282 -37 291 -35
rect 293 -37 295 -35
rect 290 -42 295 -37
rect 290 -44 291 -42
rect 293 -44 295 -42
rect 290 -46 295 -44
rect 334 -26 348 -25
rect 334 -28 342 -26
rect 344 -28 348 -26
rect 334 -29 348 -28
rect 318 -36 332 -33
rect 318 -38 319 -36
rect 321 -37 332 -36
rect 342 -37 348 -29
rect 321 -38 324 -37
rect 318 -45 324 -38
rect 438 -15 443 -13
rect 438 -17 439 -15
rect 441 -17 443 -15
rect 438 -19 443 -17
rect 439 -33 443 -19
rect 430 -35 443 -33
rect 430 -37 439 -35
rect 441 -37 443 -35
rect 438 -42 443 -37
rect 438 -44 439 -42
rect 441 -44 443 -42
rect 438 -46 443 -44
rect 482 -26 496 -25
rect 482 -28 490 -26
rect 492 -28 496 -26
rect 482 -29 496 -28
rect 466 -36 480 -33
rect 466 -38 467 -36
rect 469 -37 480 -36
rect 490 -37 496 -29
rect 469 -38 472 -37
rect 466 -45 472 -38
rect 586 -15 591 -13
rect 586 -17 587 -15
rect 589 -17 591 -15
rect 586 -19 591 -17
rect 587 -33 591 -19
rect 578 -35 591 -33
rect 578 -37 587 -35
rect 589 -37 591 -35
rect 586 -42 591 -37
rect 586 -44 587 -42
rect 589 -44 591 -42
rect 586 -46 591 -44
rect 630 -26 644 -25
rect 630 -28 638 -26
rect 640 -28 644 -26
rect 630 -29 644 -28
rect 614 -36 628 -33
rect 614 -38 615 -36
rect 617 -37 628 -36
rect 638 -37 644 -29
rect 617 -38 620 -37
rect 614 -45 620 -38
rect 734 -15 739 -13
rect 734 -17 735 -15
rect 737 -17 739 -15
rect 734 -19 739 -17
rect 735 -33 739 -19
rect 726 -35 739 -33
rect 726 -37 735 -35
rect 737 -37 739 -35
rect 734 -42 739 -37
rect 734 -44 735 -42
rect 737 -44 739 -42
rect 734 -46 739 -44
rect 778 -26 792 -25
rect 778 -28 786 -26
rect 788 -28 792 -26
rect 778 -29 792 -28
rect 762 -36 776 -33
rect 762 -38 763 -36
rect 765 -37 776 -36
rect 786 -37 792 -29
rect 765 -38 768 -37
rect 762 -45 768 -38
rect 882 -15 887 -13
rect 882 -17 883 -15
rect 885 -17 887 -15
rect 882 -19 887 -17
rect 883 -33 887 -19
rect 874 -35 887 -33
rect 874 -37 883 -35
rect 885 -37 887 -35
rect 882 -42 887 -37
rect 882 -44 883 -42
rect 885 -44 887 -42
rect 882 -46 887 -44
rect 926 -26 940 -25
rect 926 -28 934 -26
rect 936 -28 940 -26
rect 926 -29 940 -28
rect 910 -36 924 -33
rect 910 -38 911 -36
rect 913 -37 924 -36
rect 934 -37 940 -29
rect 913 -38 916 -37
rect 910 -45 916 -38
rect 1030 -15 1035 -13
rect 1030 -17 1031 -15
rect 1033 -17 1035 -15
rect 1030 -19 1035 -17
rect 1031 -33 1035 -19
rect 1022 -35 1035 -33
rect 1022 -37 1031 -35
rect 1033 -37 1035 -35
rect 1030 -42 1035 -37
rect 1030 -44 1031 -42
rect 1033 -44 1035 -42
rect 1030 -46 1035 -44
rect 1074 -26 1088 -25
rect 1074 -28 1082 -26
rect 1084 -28 1088 -26
rect 1074 -29 1088 -28
rect 1058 -36 1072 -33
rect 1058 -38 1059 -36
rect 1061 -37 1072 -36
rect 1082 -37 1088 -29
rect 1061 -38 1064 -37
rect 1058 -45 1064 -38
rect 1178 -15 1183 -13
rect 1178 -17 1179 -15
rect 1181 -17 1183 -15
rect 1178 -19 1183 -17
rect 1179 -33 1183 -19
rect 1170 -35 1183 -33
rect 1170 -37 1179 -35
rect 1181 -37 1183 -35
rect 1178 -42 1183 -37
rect 1178 -44 1179 -42
rect 1181 -44 1183 -42
rect 1178 -46 1183 -44
rect 3 -60 1187 -59
rect 3 -62 28 -60
rect 30 -62 109 -60
rect 111 -62 119 -60
rect 121 -62 176 -60
rect 178 -62 257 -60
rect 259 -62 267 -60
rect 269 -62 324 -60
rect 326 -62 405 -60
rect 407 -62 415 -60
rect 417 -62 472 -60
rect 474 -62 553 -60
rect 555 -62 563 -60
rect 565 -62 620 -60
rect 622 -62 701 -60
rect 703 -62 711 -60
rect 713 -62 768 -60
rect 770 -62 849 -60
rect 851 -62 859 -60
rect 861 -62 916 -60
rect 918 -62 997 -60
rect 999 -62 1007 -60
rect 1009 -62 1064 -60
rect 1066 -62 1145 -60
rect 1147 -62 1155 -60
rect 1157 -62 1187 -60
rect 3 -67 1187 -62
rect 122 -72 150 -67
rect 122 -74 129 -72
rect 131 -74 141 -72
rect 143 -74 150 -72
rect 122 -75 150 -74
rect 126 -90 138 -88
rect 126 -92 128 -90
rect 130 -92 138 -90
rect 126 -94 138 -92
rect 126 -97 130 -94
rect 126 -99 128 -97
rect 126 -115 130 -99
rect 134 -106 146 -104
rect 134 -108 135 -106
rect 137 -107 146 -106
rect 137 -108 141 -107
rect 134 -109 141 -108
rect 143 -109 146 -107
rect 134 -110 146 -109
rect 126 -117 128 -115
rect 126 -126 130 -117
rect 134 -118 138 -110
rect 122 -132 150 -131
rect 122 -134 129 -132
rect 131 -134 141 -132
rect 143 -134 150 -132
rect 122 -139 150 -134
<< alu2 >>
rect 140 -38 146 -33
rect 140 -40 143 -38
rect 145 -40 146 -38
rect 140 -107 146 -40
rect 140 -109 141 -107
rect 143 -109 146 -107
rect 140 -110 146 -109
<< ptie >>
rect 117 12 146 14
rect 117 10 125 12
rect 127 10 136 12
rect 138 10 146 12
rect 117 8 146 10
rect 265 12 294 14
rect 265 10 273 12
rect 275 10 284 12
rect 286 10 294 12
rect 265 8 294 10
rect 413 12 442 14
rect 413 10 421 12
rect 423 10 432 12
rect 434 10 442 12
rect 413 8 442 10
rect 561 12 590 14
rect 561 10 569 12
rect 571 10 580 12
rect 582 10 590 12
rect 561 8 590 10
rect 709 12 738 14
rect 709 10 717 12
rect 719 10 728 12
rect 730 10 738 12
rect 709 8 738 10
rect 857 12 886 14
rect 857 10 865 12
rect 867 10 876 12
rect 878 10 886 12
rect 857 8 886 10
rect 1005 12 1034 14
rect 1005 10 1013 12
rect 1015 10 1024 12
rect 1026 10 1034 12
rect 1005 8 1034 10
rect 1153 12 1182 14
rect 1153 10 1161 12
rect 1163 10 1172 12
rect 1174 10 1182 12
rect 1153 8 1182 10
rect 8 0 37 2
rect 8 -2 16 0
rect 18 -2 27 0
rect 29 -2 37 0
rect 8 -4 37 -2
rect 156 0 185 2
rect 156 -2 164 0
rect 166 -2 175 0
rect 177 -2 185 0
rect 156 -4 185 -2
rect 304 0 333 2
rect 304 -2 312 0
rect 314 -2 323 0
rect 325 -2 333 0
rect 304 -4 333 -2
rect 452 0 481 2
rect 452 -2 460 0
rect 462 -2 471 0
rect 473 -2 481 0
rect 452 -4 481 -2
rect 600 0 629 2
rect 600 -2 608 0
rect 610 -2 619 0
rect 621 -2 629 0
rect 600 -4 629 -2
rect 748 0 777 2
rect 748 -2 756 0
rect 758 -2 767 0
rect 769 -2 777 0
rect 748 -4 777 -2
rect 896 0 925 2
rect 896 -2 904 0
rect 906 -2 915 0
rect 917 -2 925 0
rect 896 -4 925 -2
rect 1044 0 1073 2
rect 1044 -2 1052 0
rect 1054 -2 1063 0
rect 1065 -2 1073 0
rect 1044 -4 1073 -2
rect 127 -132 145 -130
rect 127 -134 129 -132
rect 131 -134 141 -132
rect 143 -134 145 -132
rect 127 -136 145 -134
<< ntie >>
rect 27 72 51 74
rect 27 70 33 72
rect 35 70 43 72
rect 45 70 51 72
rect 27 68 51 70
rect 122 72 128 74
rect 122 70 124 72
rect 126 70 128 72
rect 175 72 199 74
rect 122 68 128 70
rect 175 70 181 72
rect 183 70 191 72
rect 193 70 199 72
rect 175 68 199 70
rect 270 72 276 74
rect 270 70 272 72
rect 274 70 276 72
rect 323 72 347 74
rect 270 68 276 70
rect 323 70 329 72
rect 331 70 339 72
rect 341 70 347 72
rect 323 68 347 70
rect 418 72 424 74
rect 418 70 420 72
rect 422 70 424 72
rect 471 72 495 74
rect 418 68 424 70
rect 471 70 477 72
rect 479 70 487 72
rect 489 70 495 72
rect 471 68 495 70
rect 566 72 572 74
rect 566 70 568 72
rect 570 70 572 72
rect 619 72 643 74
rect 566 68 572 70
rect 619 70 625 72
rect 627 70 635 72
rect 637 70 643 72
rect 619 68 643 70
rect 714 72 720 74
rect 714 70 716 72
rect 718 70 720 72
rect 767 72 791 74
rect 714 68 720 70
rect 767 70 773 72
rect 775 70 783 72
rect 785 70 791 72
rect 767 68 791 70
rect 862 72 868 74
rect 862 70 864 72
rect 866 70 868 72
rect 915 72 939 74
rect 862 68 868 70
rect 915 70 921 72
rect 923 70 931 72
rect 933 70 939 72
rect 915 68 939 70
rect 1010 72 1016 74
rect 1010 70 1012 72
rect 1014 70 1016 72
rect 1063 72 1087 74
rect 1010 68 1016 70
rect 1063 70 1069 72
rect 1071 70 1079 72
rect 1081 70 1087 72
rect 1063 68 1087 70
rect 1158 72 1164 74
rect 1158 70 1160 72
rect 1162 70 1164 72
rect 1158 68 1164 70
rect 26 -60 32 -58
rect 26 -62 28 -60
rect 30 -62 32 -60
rect 26 -64 32 -62
rect 103 -60 127 -58
rect 103 -62 109 -60
rect 111 -62 119 -60
rect 121 -62 127 -60
rect 174 -60 180 -58
rect 103 -64 127 -62
rect 174 -62 176 -60
rect 178 -62 180 -60
rect 174 -64 180 -62
rect 251 -60 275 -58
rect 251 -62 257 -60
rect 259 -62 267 -60
rect 269 -62 275 -60
rect 322 -60 328 -58
rect 251 -64 275 -62
rect 322 -62 324 -60
rect 326 -62 328 -60
rect 322 -64 328 -62
rect 399 -60 423 -58
rect 399 -62 405 -60
rect 407 -62 415 -60
rect 417 -62 423 -60
rect 470 -60 476 -58
rect 399 -64 423 -62
rect 470 -62 472 -60
rect 474 -62 476 -60
rect 470 -64 476 -62
rect 547 -60 571 -58
rect 547 -62 553 -60
rect 555 -62 563 -60
rect 565 -62 571 -60
rect 618 -60 624 -58
rect 547 -64 571 -62
rect 618 -62 620 -60
rect 622 -62 624 -60
rect 618 -64 624 -62
rect 695 -60 719 -58
rect 695 -62 701 -60
rect 703 -62 711 -60
rect 713 -62 719 -60
rect 766 -60 772 -58
rect 695 -64 719 -62
rect 766 -62 768 -60
rect 770 -62 772 -60
rect 766 -64 772 -62
rect 843 -60 867 -58
rect 843 -62 849 -60
rect 851 -62 859 -60
rect 861 -62 867 -60
rect 914 -60 920 -58
rect 843 -64 867 -62
rect 914 -62 916 -60
rect 918 -62 920 -60
rect 914 -64 920 -62
rect 991 -60 1015 -58
rect 991 -62 997 -60
rect 999 -62 1007 -60
rect 1009 -62 1015 -60
rect 1062 -60 1068 -58
rect 991 -64 1015 -62
rect 1062 -62 1064 -60
rect 1066 -62 1068 -60
rect 1062 -64 1068 -62
rect 1139 -60 1163 -58
rect 1139 -62 1145 -60
rect 1147 -62 1155 -60
rect 1157 -62 1163 -60
rect 1139 -64 1163 -62
rect 127 -72 145 -70
rect 127 -74 129 -72
rect 131 -74 141 -72
rect 143 -74 145 -72
rect 127 -76 145 -74
<< nmos >>
rect 14 15 16 29
rect 32 24 34 31
rect 124 25 126 31
rect 43 18 45 24
rect 50 18 52 24
rect 60 18 62 24
rect 70 18 72 24
rect 80 18 82 24
rect 87 18 89 24
rect 97 18 99 24
rect 104 18 106 24
rect 134 24 136 31
rect 162 15 164 29
rect 180 24 182 31
rect 272 25 274 31
rect 191 18 193 24
rect 198 18 200 24
rect 208 18 210 24
rect 218 18 220 24
rect 228 18 230 24
rect 235 18 237 24
rect 245 18 247 24
rect 252 18 254 24
rect 282 24 284 31
rect 310 15 312 29
rect 328 24 330 31
rect 420 25 422 31
rect 339 18 341 24
rect 346 18 348 24
rect 356 18 358 24
rect 366 18 368 24
rect 376 18 378 24
rect 383 18 385 24
rect 393 18 395 24
rect 400 18 402 24
rect 430 24 432 31
rect 458 15 460 29
rect 476 24 478 31
rect 568 25 570 31
rect 487 18 489 24
rect 494 18 496 24
rect 504 18 506 24
rect 514 18 516 24
rect 524 18 526 24
rect 531 18 533 24
rect 541 18 543 24
rect 548 18 550 24
rect 578 24 580 31
rect 606 15 608 29
rect 624 24 626 31
rect 716 25 718 31
rect 635 18 637 24
rect 642 18 644 24
rect 652 18 654 24
rect 662 18 664 24
rect 672 18 674 24
rect 679 18 681 24
rect 689 18 691 24
rect 696 18 698 24
rect 726 24 728 31
rect 754 15 756 29
rect 772 24 774 31
rect 864 25 866 31
rect 783 18 785 24
rect 790 18 792 24
rect 800 18 802 24
rect 810 18 812 24
rect 820 18 822 24
rect 827 18 829 24
rect 837 18 839 24
rect 844 18 846 24
rect 874 24 876 31
rect 902 15 904 29
rect 920 24 922 31
rect 1012 25 1014 31
rect 931 18 933 24
rect 938 18 940 24
rect 948 18 950 24
rect 958 18 960 24
rect 968 18 970 24
rect 975 18 977 24
rect 985 18 987 24
rect 992 18 994 24
rect 1022 24 1024 31
rect 1050 15 1052 29
rect 1068 24 1070 31
rect 1160 25 1162 31
rect 1079 18 1081 24
rect 1086 18 1088 24
rect 1096 18 1098 24
rect 1106 18 1108 24
rect 1116 18 1118 24
rect 1123 18 1125 24
rect 1133 18 1135 24
rect 1140 18 1142 24
rect 1170 24 1172 31
rect 18 -21 20 -14
rect 48 -14 50 -8
rect 55 -14 57 -8
rect 65 -14 67 -8
rect 72 -14 74 -8
rect 82 -14 84 -8
rect 92 -14 94 -8
rect 102 -14 104 -8
rect 109 -14 111 -8
rect 28 -21 30 -15
rect 120 -21 122 -14
rect 138 -19 140 -5
rect 166 -21 168 -14
rect 196 -14 198 -8
rect 203 -14 205 -8
rect 213 -14 215 -8
rect 220 -14 222 -8
rect 230 -14 232 -8
rect 240 -14 242 -8
rect 250 -14 252 -8
rect 257 -14 259 -8
rect 176 -21 178 -15
rect 268 -21 270 -14
rect 286 -19 288 -5
rect 314 -21 316 -14
rect 344 -14 346 -8
rect 351 -14 353 -8
rect 361 -14 363 -8
rect 368 -14 370 -8
rect 378 -14 380 -8
rect 388 -14 390 -8
rect 398 -14 400 -8
rect 405 -14 407 -8
rect 324 -21 326 -15
rect 416 -21 418 -14
rect 434 -19 436 -5
rect 462 -21 464 -14
rect 492 -14 494 -8
rect 499 -14 501 -8
rect 509 -14 511 -8
rect 516 -14 518 -8
rect 526 -14 528 -8
rect 536 -14 538 -8
rect 546 -14 548 -8
rect 553 -14 555 -8
rect 472 -21 474 -15
rect 564 -21 566 -14
rect 582 -19 584 -5
rect 610 -21 612 -14
rect 640 -14 642 -8
rect 647 -14 649 -8
rect 657 -14 659 -8
rect 664 -14 666 -8
rect 674 -14 676 -8
rect 684 -14 686 -8
rect 694 -14 696 -8
rect 701 -14 703 -8
rect 620 -21 622 -15
rect 712 -21 714 -14
rect 730 -19 732 -5
rect 758 -21 760 -14
rect 788 -14 790 -8
rect 795 -14 797 -8
rect 805 -14 807 -8
rect 812 -14 814 -8
rect 822 -14 824 -8
rect 832 -14 834 -8
rect 842 -14 844 -8
rect 849 -14 851 -8
rect 768 -21 770 -15
rect 860 -21 862 -14
rect 878 -19 880 -5
rect 906 -21 908 -14
rect 936 -14 938 -8
rect 943 -14 945 -8
rect 953 -14 955 -8
rect 960 -14 962 -8
rect 970 -14 972 -8
rect 980 -14 982 -8
rect 990 -14 992 -8
rect 997 -14 999 -8
rect 916 -21 918 -15
rect 1008 -21 1010 -14
rect 1026 -19 1028 -5
rect 1054 -21 1056 -14
rect 1084 -14 1086 -8
rect 1091 -14 1093 -8
rect 1101 -14 1103 -8
rect 1108 -14 1110 -8
rect 1118 -14 1120 -8
rect 1128 -14 1130 -8
rect 1138 -14 1140 -8
rect 1145 -14 1147 -8
rect 1064 -21 1066 -15
rect 1156 -21 1158 -14
rect 1174 -19 1176 -5
rect 133 -122 135 -113
<< pmos >>
rect 14 43 16 71
rect 24 43 26 57
rect 43 53 45 59
rect 50 53 52 59
rect 60 53 62 65
rect 70 53 72 65
rect 80 59 82 65
rect 87 59 89 65
rect 97 52 99 65
rect 104 52 106 65
rect 114 52 116 63
rect 134 54 136 64
rect 162 43 164 71
rect 172 43 174 57
rect 191 53 193 59
rect 198 53 200 59
rect 208 53 210 65
rect 218 53 220 65
rect 228 59 230 65
rect 235 59 237 65
rect 245 52 247 65
rect 252 52 254 65
rect 262 52 264 63
rect 282 54 284 64
rect 310 43 312 71
rect 320 43 322 57
rect 339 53 341 59
rect 346 53 348 59
rect 356 53 358 65
rect 366 53 368 65
rect 376 59 378 65
rect 383 59 385 65
rect 393 52 395 65
rect 400 52 402 65
rect 410 52 412 63
rect 430 54 432 64
rect 458 43 460 71
rect 468 43 470 57
rect 487 53 489 59
rect 494 53 496 59
rect 504 53 506 65
rect 514 53 516 65
rect 524 59 526 65
rect 531 59 533 65
rect 541 52 543 65
rect 548 52 550 65
rect 558 52 560 63
rect 578 54 580 64
rect 606 43 608 71
rect 616 43 618 57
rect 635 53 637 59
rect 642 53 644 59
rect 652 53 654 65
rect 662 53 664 65
rect 672 59 674 65
rect 679 59 681 65
rect 689 52 691 65
rect 696 52 698 65
rect 706 52 708 63
rect 726 54 728 64
rect 754 43 756 71
rect 764 43 766 57
rect 783 53 785 59
rect 790 53 792 59
rect 800 53 802 65
rect 810 53 812 65
rect 820 59 822 65
rect 827 59 829 65
rect 837 52 839 65
rect 844 52 846 65
rect 854 52 856 63
rect 874 54 876 64
rect 902 43 904 71
rect 912 43 914 57
rect 931 53 933 59
rect 938 53 940 59
rect 948 53 950 65
rect 958 53 960 65
rect 968 59 970 65
rect 975 59 977 65
rect 985 52 987 65
rect 992 52 994 65
rect 1002 52 1004 63
rect 1022 54 1024 64
rect 1050 43 1052 71
rect 1060 43 1062 57
rect 1079 53 1081 59
rect 1086 53 1088 59
rect 1096 53 1098 65
rect 1106 53 1108 65
rect 1116 59 1118 65
rect 1123 59 1125 65
rect 1133 52 1135 65
rect 1140 52 1142 65
rect 1150 52 1152 63
rect 1170 54 1172 64
rect 18 -54 20 -44
rect 38 -53 40 -42
rect 48 -55 50 -42
rect 55 -55 57 -42
rect 65 -55 67 -49
rect 72 -55 74 -49
rect 82 -55 84 -43
rect 92 -55 94 -43
rect 102 -49 104 -43
rect 109 -49 111 -43
rect 128 -47 130 -33
rect 138 -61 140 -33
rect 166 -54 168 -44
rect 186 -53 188 -42
rect 196 -55 198 -42
rect 203 -55 205 -42
rect 213 -55 215 -49
rect 220 -55 222 -49
rect 230 -55 232 -43
rect 240 -55 242 -43
rect 250 -49 252 -43
rect 257 -49 259 -43
rect 276 -47 278 -33
rect 286 -61 288 -33
rect 314 -54 316 -44
rect 334 -53 336 -42
rect 344 -55 346 -42
rect 351 -55 353 -42
rect 361 -55 363 -49
rect 368 -55 370 -49
rect 378 -55 380 -43
rect 388 -55 390 -43
rect 398 -49 400 -43
rect 405 -49 407 -43
rect 424 -47 426 -33
rect 434 -61 436 -33
rect 462 -54 464 -44
rect 482 -53 484 -42
rect 492 -55 494 -42
rect 499 -55 501 -42
rect 509 -55 511 -49
rect 516 -55 518 -49
rect 526 -55 528 -43
rect 536 -55 538 -43
rect 546 -49 548 -43
rect 553 -49 555 -43
rect 572 -47 574 -33
rect 582 -61 584 -33
rect 610 -54 612 -44
rect 630 -53 632 -42
rect 640 -55 642 -42
rect 647 -55 649 -42
rect 657 -55 659 -49
rect 664 -55 666 -49
rect 674 -55 676 -43
rect 684 -55 686 -43
rect 694 -49 696 -43
rect 701 -49 703 -43
rect 720 -47 722 -33
rect 730 -61 732 -33
rect 758 -54 760 -44
rect 778 -53 780 -42
rect 788 -55 790 -42
rect 795 -55 797 -42
rect 805 -55 807 -49
rect 812 -55 814 -49
rect 822 -55 824 -43
rect 832 -55 834 -43
rect 842 -49 844 -43
rect 849 -49 851 -43
rect 868 -47 870 -33
rect 878 -61 880 -33
rect 906 -54 908 -44
rect 926 -53 928 -42
rect 936 -55 938 -42
rect 943 -55 945 -42
rect 953 -55 955 -49
rect 960 -55 962 -49
rect 970 -55 972 -43
rect 980 -55 982 -43
rect 990 -49 992 -43
rect 997 -49 999 -43
rect 1016 -47 1018 -33
rect 1026 -61 1028 -33
rect 1054 -54 1056 -44
rect 1074 -53 1076 -42
rect 1084 -55 1086 -42
rect 1091 -55 1093 -42
rect 1101 -55 1103 -49
rect 1108 -55 1110 -49
rect 1118 -55 1120 -43
rect 1128 -55 1130 -43
rect 1138 -49 1140 -43
rect 1145 -49 1147 -43
rect 1164 -47 1166 -33
rect 1174 -61 1176 -33
rect 133 -101 135 -83
<< polyct0 >>
rect 16 35 18 37
rect 35 36 37 38
rect 52 45 54 47
rect 78 45 80 47
rect 58 29 60 31
rect 72 30 74 32
rect 95 45 97 47
rect 89 29 91 31
rect 122 36 124 38
rect 164 35 166 37
rect 183 36 185 38
rect 200 45 202 47
rect 226 45 228 47
rect 206 29 208 31
rect 220 30 222 32
rect 243 45 245 47
rect 237 29 239 31
rect 270 36 272 38
rect 312 35 314 37
rect 331 36 333 38
rect 348 45 350 47
rect 374 45 376 47
rect 354 29 356 31
rect 368 30 370 32
rect 391 45 393 47
rect 385 29 387 31
rect 418 36 420 38
rect 460 35 462 37
rect 479 36 481 38
rect 496 45 498 47
rect 522 45 524 47
rect 502 29 504 31
rect 516 30 518 32
rect 539 45 541 47
rect 533 29 535 31
rect 566 36 568 38
rect 608 35 610 37
rect 627 36 629 38
rect 644 45 646 47
rect 670 45 672 47
rect 650 29 652 31
rect 664 30 666 32
rect 687 45 689 47
rect 681 29 683 31
rect 714 36 716 38
rect 756 35 758 37
rect 775 36 777 38
rect 792 45 794 47
rect 818 45 820 47
rect 798 29 800 31
rect 812 30 814 32
rect 835 45 837 47
rect 829 29 831 31
rect 862 36 864 38
rect 904 35 906 37
rect 923 36 925 38
rect 940 45 942 47
rect 966 45 968 47
rect 946 29 948 31
rect 960 30 962 32
rect 983 45 985 47
rect 977 29 979 31
rect 1010 36 1012 38
rect 1052 35 1054 37
rect 1071 36 1073 38
rect 1088 45 1090 47
rect 1114 45 1116 47
rect 1094 29 1096 31
rect 1108 30 1110 32
rect 1131 45 1133 47
rect 1125 29 1127 31
rect 1158 36 1160 38
rect 30 -28 32 -26
rect 63 -21 65 -19
rect 57 -37 59 -35
rect 80 -22 82 -20
rect 94 -21 96 -19
rect 74 -37 76 -35
rect 100 -37 102 -35
rect 117 -28 119 -26
rect 136 -27 138 -25
rect 178 -28 180 -26
rect 211 -21 213 -19
rect 205 -37 207 -35
rect 228 -22 230 -20
rect 242 -21 244 -19
rect 222 -37 224 -35
rect 248 -37 250 -35
rect 265 -28 267 -26
rect 284 -27 286 -25
rect 326 -28 328 -26
rect 359 -21 361 -19
rect 353 -37 355 -35
rect 376 -22 378 -20
rect 390 -21 392 -19
rect 370 -37 372 -35
rect 396 -37 398 -35
rect 413 -28 415 -26
rect 432 -27 434 -25
rect 474 -28 476 -26
rect 507 -21 509 -19
rect 501 -37 503 -35
rect 524 -22 526 -20
rect 538 -21 540 -19
rect 518 -37 520 -35
rect 544 -37 546 -35
rect 561 -28 563 -26
rect 580 -27 582 -25
rect 622 -28 624 -26
rect 655 -21 657 -19
rect 649 -37 651 -35
rect 672 -22 674 -20
rect 686 -21 688 -19
rect 666 -37 668 -35
rect 692 -37 694 -35
rect 709 -28 711 -26
rect 728 -27 730 -25
rect 770 -28 772 -26
rect 803 -21 805 -19
rect 797 -37 799 -35
rect 820 -22 822 -20
rect 834 -21 836 -19
rect 814 -37 816 -35
rect 840 -37 842 -35
rect 857 -28 859 -26
rect 876 -27 878 -25
rect 918 -28 920 -26
rect 951 -21 953 -19
rect 945 -37 947 -35
rect 968 -22 970 -20
rect 982 -21 984 -19
rect 962 -37 964 -35
rect 988 -37 990 -35
rect 1005 -28 1007 -26
rect 1024 -27 1026 -25
rect 1066 -28 1068 -26
rect 1099 -21 1101 -19
rect 1093 -37 1095 -35
rect 1116 -22 1118 -20
rect 1130 -21 1132 -19
rect 1110 -37 1112 -35
rect 1136 -37 1138 -35
rect 1153 -28 1155 -26
rect 1172 -27 1174 -25
<< polyct1 >>
rect 129 46 131 48
rect 106 36 108 38
rect 277 46 279 48
rect 254 36 256 38
rect 425 46 427 48
rect 402 36 404 38
rect 573 46 575 48
rect 550 36 552 38
rect 721 46 723 48
rect 698 36 700 38
rect 869 46 871 48
rect 846 36 848 38
rect 1017 46 1019 48
rect 994 36 996 38
rect 1165 46 1167 48
rect 1142 36 1144 38
rect 46 -28 48 -26
rect 23 -38 25 -36
rect 194 -28 196 -26
rect 171 -38 173 -36
rect 342 -28 344 -26
rect 319 -38 321 -36
rect 490 -28 492 -26
rect 467 -38 469 -36
rect 638 -28 640 -26
rect 615 -38 617 -36
rect 786 -28 788 -26
rect 763 -38 765 -36
rect 934 -28 936 -26
rect 911 -38 913 -36
rect 1082 -28 1084 -26
rect 1059 -38 1061 -36
rect 135 -108 137 -106
<< ndifct0 >>
rect 27 27 29 29
rect 119 27 121 29
rect 129 27 131 29
rect 38 20 40 22
rect 19 17 21 19
rect 55 20 57 22
rect 65 20 67 22
rect 75 20 77 22
rect 92 20 94 22
rect 109 20 111 22
rect 139 27 141 29
rect 175 27 177 29
rect 267 27 269 29
rect 277 27 279 29
rect 186 20 188 22
rect 167 17 169 19
rect 203 20 205 22
rect 213 20 215 22
rect 223 20 225 22
rect 240 20 242 22
rect 257 20 259 22
rect 287 27 289 29
rect 323 27 325 29
rect 415 27 417 29
rect 425 27 427 29
rect 334 20 336 22
rect 315 17 317 19
rect 351 20 353 22
rect 361 20 363 22
rect 371 20 373 22
rect 388 20 390 22
rect 405 20 407 22
rect 435 27 437 29
rect 471 27 473 29
rect 563 27 565 29
rect 573 27 575 29
rect 482 20 484 22
rect 463 17 465 19
rect 499 20 501 22
rect 509 20 511 22
rect 519 20 521 22
rect 536 20 538 22
rect 553 20 555 22
rect 583 27 585 29
rect 619 27 621 29
rect 711 27 713 29
rect 721 27 723 29
rect 630 20 632 22
rect 611 17 613 19
rect 647 20 649 22
rect 657 20 659 22
rect 667 20 669 22
rect 684 20 686 22
rect 701 20 703 22
rect 731 27 733 29
rect 767 27 769 29
rect 859 27 861 29
rect 869 27 871 29
rect 778 20 780 22
rect 759 17 761 19
rect 795 20 797 22
rect 805 20 807 22
rect 815 20 817 22
rect 832 20 834 22
rect 849 20 851 22
rect 879 27 881 29
rect 915 27 917 29
rect 1007 27 1009 29
rect 1017 27 1019 29
rect 926 20 928 22
rect 907 17 909 19
rect 943 20 945 22
rect 953 20 955 22
rect 963 20 965 22
rect 980 20 982 22
rect 997 20 999 22
rect 1027 27 1029 29
rect 1063 27 1065 29
rect 1155 27 1157 29
rect 1165 27 1167 29
rect 1074 20 1076 22
rect 1055 17 1057 19
rect 1091 20 1093 22
rect 1101 20 1103 22
rect 1111 20 1113 22
rect 1128 20 1130 22
rect 1145 20 1147 22
rect 1175 27 1177 29
rect 13 -19 15 -17
rect 43 -12 45 -10
rect 60 -12 62 -10
rect 77 -12 79 -10
rect 87 -12 89 -10
rect 97 -12 99 -10
rect 133 -9 135 -7
rect 114 -12 116 -10
rect 23 -19 25 -17
rect 33 -19 35 -17
rect 125 -19 127 -17
rect 161 -19 163 -17
rect 191 -12 193 -10
rect 208 -12 210 -10
rect 225 -12 227 -10
rect 235 -12 237 -10
rect 245 -12 247 -10
rect 281 -9 283 -7
rect 262 -12 264 -10
rect 171 -19 173 -17
rect 181 -19 183 -17
rect 273 -19 275 -17
rect 309 -19 311 -17
rect 339 -12 341 -10
rect 356 -12 358 -10
rect 373 -12 375 -10
rect 383 -12 385 -10
rect 393 -12 395 -10
rect 429 -9 431 -7
rect 410 -12 412 -10
rect 319 -19 321 -17
rect 329 -19 331 -17
rect 421 -19 423 -17
rect 457 -19 459 -17
rect 487 -12 489 -10
rect 504 -12 506 -10
rect 521 -12 523 -10
rect 531 -12 533 -10
rect 541 -12 543 -10
rect 577 -9 579 -7
rect 558 -12 560 -10
rect 467 -19 469 -17
rect 477 -19 479 -17
rect 569 -19 571 -17
rect 605 -19 607 -17
rect 635 -12 637 -10
rect 652 -12 654 -10
rect 669 -12 671 -10
rect 679 -12 681 -10
rect 689 -12 691 -10
rect 725 -9 727 -7
rect 706 -12 708 -10
rect 615 -19 617 -17
rect 625 -19 627 -17
rect 717 -19 719 -17
rect 753 -19 755 -17
rect 783 -12 785 -10
rect 800 -12 802 -10
rect 817 -12 819 -10
rect 827 -12 829 -10
rect 837 -12 839 -10
rect 873 -9 875 -7
rect 854 -12 856 -10
rect 763 -19 765 -17
rect 773 -19 775 -17
rect 865 -19 867 -17
rect 901 -19 903 -17
rect 931 -12 933 -10
rect 948 -12 950 -10
rect 965 -12 967 -10
rect 975 -12 977 -10
rect 985 -12 987 -10
rect 1021 -9 1023 -7
rect 1002 -12 1004 -10
rect 911 -19 913 -17
rect 921 -19 923 -17
rect 1013 -19 1015 -17
rect 1049 -19 1051 -17
rect 1079 -12 1081 -10
rect 1096 -12 1098 -10
rect 1113 -12 1115 -10
rect 1123 -12 1125 -10
rect 1133 -12 1135 -10
rect 1169 -9 1171 -7
rect 1150 -12 1152 -10
rect 1059 -19 1061 -17
rect 1069 -19 1071 -17
rect 1161 -19 1163 -17
rect 142 -120 144 -118
<< ndifct1 >>
rect 9 25 11 27
rect 157 25 159 27
rect 305 25 307 27
rect 453 25 455 27
rect 601 25 603 27
rect 749 25 751 27
rect 897 25 899 27
rect 1045 25 1047 27
rect 143 -17 145 -15
rect 291 -17 293 -15
rect 439 -17 441 -15
rect 587 -17 589 -15
rect 735 -17 737 -15
rect 883 -17 885 -15
rect 1031 -17 1033 -15
rect 1179 -17 1181 -15
rect 128 -117 130 -115
<< ntiect1 >>
rect 33 70 35 72
rect 43 70 45 72
rect 124 70 126 72
rect 181 70 183 72
rect 191 70 193 72
rect 272 70 274 72
rect 329 70 331 72
rect 339 70 341 72
rect 420 70 422 72
rect 477 70 479 72
rect 487 70 489 72
rect 568 70 570 72
rect 625 70 627 72
rect 635 70 637 72
rect 716 70 718 72
rect 773 70 775 72
rect 783 70 785 72
rect 864 70 866 72
rect 921 70 923 72
rect 931 70 933 72
rect 1012 70 1014 72
rect 1069 70 1071 72
rect 1079 70 1081 72
rect 1160 70 1162 72
rect 28 -62 30 -60
rect 109 -62 111 -60
rect 119 -62 121 -60
rect 176 -62 178 -60
rect 257 -62 259 -60
rect 267 -62 269 -60
rect 324 -62 326 -60
rect 405 -62 407 -60
rect 415 -62 417 -60
rect 472 -62 474 -60
rect 553 -62 555 -60
rect 563 -62 565 -60
rect 620 -62 622 -60
rect 701 -62 703 -60
rect 711 -62 713 -60
rect 768 -62 770 -60
rect 849 -62 851 -60
rect 859 -62 861 -60
rect 916 -62 918 -60
rect 997 -62 999 -60
rect 1007 -62 1009 -60
rect 1064 -62 1066 -60
rect 1145 -62 1147 -60
rect 1155 -62 1157 -60
rect 129 -74 131 -72
rect 141 -74 143 -72
<< ptiect1 >>
rect 125 10 127 12
rect 136 10 138 12
rect 273 10 275 12
rect 284 10 286 12
rect 421 10 423 12
rect 432 10 434 12
rect 569 10 571 12
rect 580 10 582 12
rect 717 10 719 12
rect 728 10 730 12
rect 865 10 867 12
rect 876 10 878 12
rect 1013 10 1015 12
rect 1024 10 1026 12
rect 1161 10 1163 12
rect 1172 10 1174 12
rect 16 -2 18 0
rect 27 -2 29 0
rect 164 -2 166 0
rect 175 -2 177 0
rect 312 -2 314 0
rect 323 -2 325 0
rect 460 -2 462 0
rect 471 -2 473 0
rect 608 -2 610 0
rect 619 -2 621 0
rect 756 -2 758 0
rect 767 -2 769 0
rect 904 -2 906 0
rect 915 -2 917 0
rect 1052 -2 1054 0
rect 1063 -2 1065 0
rect 129 -134 131 -132
rect 141 -134 143 -132
<< pdifct0 >>
rect 19 67 21 69
rect 19 53 21 55
rect 37 55 39 57
rect 55 55 57 57
rect 65 55 67 57
rect 75 61 77 63
rect 92 61 94 63
rect 29 45 31 47
rect 109 59 111 61
rect 129 60 131 62
rect 119 54 121 56
rect 139 56 141 58
rect 167 67 169 69
rect 167 53 169 55
rect 185 55 187 57
rect 203 55 205 57
rect 213 55 215 57
rect 223 61 225 63
rect 240 61 242 63
rect 177 45 179 47
rect 257 59 259 61
rect 277 60 279 62
rect 267 54 269 56
rect 287 56 289 58
rect 315 67 317 69
rect 315 53 317 55
rect 333 55 335 57
rect 351 55 353 57
rect 361 55 363 57
rect 371 61 373 63
rect 388 61 390 63
rect 325 45 327 47
rect 405 59 407 61
rect 425 60 427 62
rect 415 54 417 56
rect 435 56 437 58
rect 463 67 465 69
rect 463 53 465 55
rect 481 55 483 57
rect 499 55 501 57
rect 509 55 511 57
rect 519 61 521 63
rect 536 61 538 63
rect 473 45 475 47
rect 553 59 555 61
rect 573 60 575 62
rect 563 54 565 56
rect 583 56 585 58
rect 611 67 613 69
rect 611 53 613 55
rect 629 55 631 57
rect 647 55 649 57
rect 657 55 659 57
rect 667 61 669 63
rect 684 61 686 63
rect 621 45 623 47
rect 701 59 703 61
rect 721 60 723 62
rect 711 54 713 56
rect 731 56 733 58
rect 759 67 761 69
rect 759 53 761 55
rect 777 55 779 57
rect 795 55 797 57
rect 805 55 807 57
rect 815 61 817 63
rect 832 61 834 63
rect 769 45 771 47
rect 849 59 851 61
rect 869 60 871 62
rect 859 54 861 56
rect 879 56 881 58
rect 907 67 909 69
rect 907 53 909 55
rect 925 55 927 57
rect 943 55 945 57
rect 953 55 955 57
rect 963 61 965 63
rect 980 61 982 63
rect 917 45 919 47
rect 997 59 999 61
rect 1017 60 1019 62
rect 1007 54 1009 56
rect 1027 56 1029 58
rect 1055 67 1057 69
rect 1055 53 1057 55
rect 1073 55 1075 57
rect 1091 55 1093 57
rect 1101 55 1103 57
rect 1111 61 1113 63
rect 1128 61 1130 63
rect 1065 45 1067 47
rect 1145 59 1147 61
rect 1165 60 1167 62
rect 1155 54 1157 56
rect 1175 56 1177 58
rect 13 -48 15 -46
rect 33 -46 35 -44
rect 23 -52 25 -50
rect 43 -51 45 -49
rect 123 -37 125 -35
rect 60 -53 62 -51
rect 77 -53 79 -51
rect 87 -47 89 -45
rect 97 -47 99 -45
rect 115 -47 117 -45
rect 133 -45 135 -43
rect 133 -59 135 -57
rect 161 -48 163 -46
rect 181 -46 183 -44
rect 171 -52 173 -50
rect 191 -51 193 -49
rect 271 -37 273 -35
rect 208 -53 210 -51
rect 225 -53 227 -51
rect 235 -47 237 -45
rect 245 -47 247 -45
rect 263 -47 265 -45
rect 281 -45 283 -43
rect 281 -59 283 -57
rect 309 -48 311 -46
rect 329 -46 331 -44
rect 319 -52 321 -50
rect 339 -51 341 -49
rect 419 -37 421 -35
rect 356 -53 358 -51
rect 373 -53 375 -51
rect 383 -47 385 -45
rect 393 -47 395 -45
rect 411 -47 413 -45
rect 429 -45 431 -43
rect 429 -59 431 -57
rect 457 -48 459 -46
rect 477 -46 479 -44
rect 467 -52 469 -50
rect 487 -51 489 -49
rect 567 -37 569 -35
rect 504 -53 506 -51
rect 521 -53 523 -51
rect 531 -47 533 -45
rect 541 -47 543 -45
rect 559 -47 561 -45
rect 577 -45 579 -43
rect 577 -59 579 -57
rect 605 -48 607 -46
rect 625 -46 627 -44
rect 615 -52 617 -50
rect 635 -51 637 -49
rect 715 -37 717 -35
rect 652 -53 654 -51
rect 669 -53 671 -51
rect 679 -47 681 -45
rect 689 -47 691 -45
rect 707 -47 709 -45
rect 725 -45 727 -43
rect 725 -59 727 -57
rect 753 -48 755 -46
rect 773 -46 775 -44
rect 763 -52 765 -50
rect 783 -51 785 -49
rect 863 -37 865 -35
rect 800 -53 802 -51
rect 817 -53 819 -51
rect 827 -47 829 -45
rect 837 -47 839 -45
rect 855 -47 857 -45
rect 873 -45 875 -43
rect 873 -59 875 -57
rect 901 -48 903 -46
rect 921 -46 923 -44
rect 911 -52 913 -50
rect 931 -51 933 -49
rect 1011 -37 1013 -35
rect 948 -53 950 -51
rect 965 -53 967 -51
rect 975 -47 977 -45
rect 985 -47 987 -45
rect 1003 -47 1005 -45
rect 1021 -45 1023 -43
rect 1021 -59 1023 -57
rect 1049 -48 1051 -46
rect 1069 -46 1071 -44
rect 1059 -52 1061 -50
rect 1079 -51 1081 -49
rect 1159 -37 1161 -35
rect 1096 -53 1098 -51
rect 1113 -53 1115 -51
rect 1123 -47 1125 -45
rect 1133 -47 1135 -45
rect 1151 -47 1153 -45
rect 1169 -45 1171 -43
rect 1169 -59 1171 -57
rect 139 -84 141 -82
<< pdifct1 >>
rect 9 52 11 54
rect 9 45 11 47
rect 157 52 159 54
rect 157 45 159 47
rect 305 52 307 54
rect 305 45 307 47
rect 453 52 455 54
rect 453 45 455 47
rect 601 52 603 54
rect 601 45 603 47
rect 749 52 751 54
rect 749 45 751 47
rect 897 52 899 54
rect 897 45 899 47
rect 1045 52 1047 54
rect 1045 45 1047 47
rect 143 -37 145 -35
rect 143 -44 145 -42
rect 291 -37 293 -35
rect 291 -44 293 -42
rect 439 -37 441 -35
rect 439 -44 441 -42
rect 587 -37 589 -35
rect 587 -44 589 -42
rect 735 -37 737 -35
rect 735 -44 737 -42
rect 883 -37 885 -35
rect 883 -44 885 -42
rect 1031 -37 1033 -35
rect 1031 -44 1033 -42
rect 1179 -37 1181 -35
rect 1179 -44 1181 -42
rect 128 -92 130 -90
rect 128 -99 130 -97
<< alu0 >>
rect 18 67 19 69
rect 21 67 22 69
rect 18 55 22 67
rect 18 53 19 55
rect 21 53 22 55
rect 36 57 40 69
rect 74 63 78 69
rect 74 61 75 63
rect 77 61 78 63
rect 74 59 78 61
rect 86 63 96 64
rect 86 61 92 63
rect 94 61 96 63
rect 86 60 96 61
rect 107 61 113 69
rect 36 55 37 57
rect 39 55 40 57
rect 36 53 40 55
rect 43 57 59 58
rect 43 55 55 57
rect 57 55 59 57
rect 43 54 59 55
rect 64 57 68 59
rect 64 55 65 57
rect 67 55 68 57
rect 18 51 22 53
rect 26 47 33 48
rect 26 45 29 47
rect 31 45 33 47
rect 26 44 33 45
rect 26 38 30 44
rect 43 39 47 54
rect 64 48 68 55
rect 50 47 59 48
rect 50 45 52 47
rect 54 45 59 47
rect 50 44 59 45
rect 14 37 30 38
rect 14 35 16 37
rect 18 35 30 37
rect 33 38 49 39
rect 33 36 35 38
rect 37 36 49 38
rect 33 35 49 36
rect 14 34 30 35
rect 26 29 30 34
rect 26 27 27 29
rect 29 27 30 29
rect 26 25 30 27
rect 37 22 41 24
rect 18 19 22 21
rect 18 17 19 19
rect 21 17 22 19
rect 18 13 22 17
rect 37 20 38 22
rect 40 20 41 22
rect 37 13 41 20
rect 45 23 49 35
rect 55 33 59 44
rect 64 47 82 48
rect 64 45 78 47
rect 80 45 82 47
rect 64 44 82 45
rect 55 31 61 33
rect 55 29 58 31
rect 60 29 61 31
rect 55 27 61 29
rect 45 22 59 23
rect 45 20 55 22
rect 57 20 59 22
rect 45 19 59 20
rect 64 22 68 44
rect 86 41 90 60
rect 107 59 109 61
rect 111 59 113 61
rect 127 62 133 69
rect 127 60 129 62
rect 131 60 133 62
rect 166 67 167 69
rect 169 67 170 69
rect 127 59 133 60
rect 107 58 113 59
rect 138 58 142 60
rect 118 56 122 58
rect 118 55 119 56
rect 81 37 90 41
rect 94 54 119 55
rect 121 54 122 56
rect 138 56 139 58
rect 141 56 142 58
rect 94 51 122 54
rect 94 47 98 51
rect 94 45 95 47
rect 97 45 98 47
rect 81 34 85 37
rect 71 32 85 34
rect 94 33 98 45
rect 138 39 142 56
rect 120 38 142 39
rect 120 36 122 38
rect 124 36 142 38
rect 120 35 142 36
rect 71 30 72 32
rect 74 30 85 32
rect 71 28 85 30
rect 64 20 65 22
rect 67 20 68 22
rect 64 18 68 20
rect 74 22 78 24
rect 74 20 75 22
rect 77 20 78 22
rect 74 13 78 20
rect 81 23 85 28
rect 88 31 98 33
rect 88 29 89 31
rect 91 29 123 31
rect 88 27 119 29
rect 121 27 123 29
rect 117 26 123 27
rect 128 29 132 31
rect 128 27 129 29
rect 131 27 132 29
rect 81 22 96 23
rect 81 20 92 22
rect 94 20 96 22
rect 81 19 96 20
rect 107 22 113 23
rect 107 20 109 22
rect 111 20 113 22
rect 107 13 113 20
rect 128 13 132 27
rect 138 29 142 35
rect 138 27 139 29
rect 141 27 142 29
rect 138 25 142 27
rect 166 55 170 67
rect 166 53 167 55
rect 169 53 170 55
rect 184 57 188 69
rect 222 63 226 69
rect 222 61 223 63
rect 225 61 226 63
rect 222 59 226 61
rect 234 63 244 64
rect 234 61 240 63
rect 242 61 244 63
rect 234 60 244 61
rect 255 61 261 69
rect 184 55 185 57
rect 187 55 188 57
rect 184 53 188 55
rect 191 57 207 58
rect 191 55 203 57
rect 205 55 207 57
rect 191 54 207 55
rect 212 57 216 59
rect 212 55 213 57
rect 215 55 216 57
rect 166 51 170 53
rect 174 47 181 48
rect 174 45 177 47
rect 179 45 181 47
rect 174 44 181 45
rect 174 38 178 44
rect 191 39 195 54
rect 212 48 216 55
rect 198 47 207 48
rect 198 45 200 47
rect 202 45 207 47
rect 198 44 207 45
rect 162 37 178 38
rect 162 35 164 37
rect 166 35 178 37
rect 181 38 197 39
rect 181 36 183 38
rect 185 36 197 38
rect 181 35 197 36
rect 162 34 178 35
rect 174 29 178 34
rect 174 27 175 29
rect 177 27 178 29
rect 174 25 178 27
rect 185 22 189 24
rect 166 19 170 21
rect 166 17 167 19
rect 169 17 170 19
rect 166 13 170 17
rect 185 20 186 22
rect 188 20 189 22
rect 185 13 189 20
rect 193 23 197 35
rect 203 33 207 44
rect 212 47 230 48
rect 212 45 226 47
rect 228 45 230 47
rect 212 44 230 45
rect 203 31 209 33
rect 203 29 206 31
rect 208 29 209 31
rect 203 27 209 29
rect 193 22 207 23
rect 193 20 203 22
rect 205 20 207 22
rect 193 19 207 20
rect 212 22 216 44
rect 234 41 238 60
rect 255 59 257 61
rect 259 59 261 61
rect 275 62 281 69
rect 275 60 277 62
rect 279 60 281 62
rect 314 67 315 69
rect 317 67 318 69
rect 275 59 281 60
rect 255 58 261 59
rect 286 58 290 60
rect 266 56 270 58
rect 266 55 267 56
rect 229 37 238 41
rect 242 54 267 55
rect 269 54 270 56
rect 286 56 287 58
rect 289 56 290 58
rect 242 51 270 54
rect 242 47 246 51
rect 242 45 243 47
rect 245 45 246 47
rect 229 34 233 37
rect 219 32 233 34
rect 242 33 246 45
rect 286 39 290 56
rect 268 38 290 39
rect 268 36 270 38
rect 272 36 290 38
rect 268 35 290 36
rect 219 30 220 32
rect 222 30 233 32
rect 219 28 233 30
rect 212 20 213 22
rect 215 20 216 22
rect 212 18 216 20
rect 222 22 226 24
rect 222 20 223 22
rect 225 20 226 22
rect 222 13 226 20
rect 229 23 233 28
rect 236 31 246 33
rect 236 29 237 31
rect 239 29 271 31
rect 236 27 267 29
rect 269 27 271 29
rect 265 26 271 27
rect 276 29 280 31
rect 276 27 277 29
rect 279 27 280 29
rect 229 22 244 23
rect 229 20 240 22
rect 242 20 244 22
rect 229 19 244 20
rect 255 22 261 23
rect 255 20 257 22
rect 259 20 261 22
rect 255 13 261 20
rect 276 13 280 27
rect 286 29 290 35
rect 286 27 287 29
rect 289 27 290 29
rect 286 25 290 27
rect 314 55 318 67
rect 314 53 315 55
rect 317 53 318 55
rect 332 57 336 69
rect 370 63 374 69
rect 370 61 371 63
rect 373 61 374 63
rect 370 59 374 61
rect 382 63 392 64
rect 382 61 388 63
rect 390 61 392 63
rect 382 60 392 61
rect 403 61 409 69
rect 332 55 333 57
rect 335 55 336 57
rect 332 53 336 55
rect 339 57 355 58
rect 339 55 351 57
rect 353 55 355 57
rect 339 54 355 55
rect 360 57 364 59
rect 360 55 361 57
rect 363 55 364 57
rect 314 51 318 53
rect 322 47 329 48
rect 322 45 325 47
rect 327 45 329 47
rect 322 44 329 45
rect 322 38 326 44
rect 339 39 343 54
rect 360 48 364 55
rect 346 47 355 48
rect 346 45 348 47
rect 350 45 355 47
rect 346 44 355 45
rect 310 37 326 38
rect 310 35 312 37
rect 314 35 326 37
rect 329 38 345 39
rect 329 36 331 38
rect 333 36 345 38
rect 329 35 345 36
rect 310 34 326 35
rect 322 29 326 34
rect 322 27 323 29
rect 325 27 326 29
rect 322 25 326 27
rect 333 22 337 24
rect 314 19 318 21
rect 314 17 315 19
rect 317 17 318 19
rect 314 13 318 17
rect 333 20 334 22
rect 336 20 337 22
rect 333 13 337 20
rect 341 23 345 35
rect 351 33 355 44
rect 360 47 378 48
rect 360 45 374 47
rect 376 45 378 47
rect 360 44 378 45
rect 351 31 357 33
rect 351 29 354 31
rect 356 29 357 31
rect 351 27 357 29
rect 341 22 355 23
rect 341 20 351 22
rect 353 20 355 22
rect 341 19 355 20
rect 360 22 364 44
rect 382 41 386 60
rect 403 59 405 61
rect 407 59 409 61
rect 423 62 429 69
rect 423 60 425 62
rect 427 60 429 62
rect 462 67 463 69
rect 465 67 466 69
rect 423 59 429 60
rect 403 58 409 59
rect 434 58 438 60
rect 414 56 418 58
rect 414 55 415 56
rect 377 37 386 41
rect 390 54 415 55
rect 417 54 418 56
rect 434 56 435 58
rect 437 56 438 58
rect 390 51 418 54
rect 390 47 394 51
rect 390 45 391 47
rect 393 45 394 47
rect 377 34 381 37
rect 367 32 381 34
rect 390 33 394 45
rect 434 39 438 56
rect 416 38 438 39
rect 416 36 418 38
rect 420 36 438 38
rect 416 35 438 36
rect 367 30 368 32
rect 370 30 381 32
rect 367 28 381 30
rect 360 20 361 22
rect 363 20 364 22
rect 360 18 364 20
rect 370 22 374 24
rect 370 20 371 22
rect 373 20 374 22
rect 370 13 374 20
rect 377 23 381 28
rect 384 31 394 33
rect 384 29 385 31
rect 387 29 419 31
rect 384 27 415 29
rect 417 27 419 29
rect 413 26 419 27
rect 424 29 428 31
rect 424 27 425 29
rect 427 27 428 29
rect 377 22 392 23
rect 377 20 388 22
rect 390 20 392 22
rect 377 19 392 20
rect 403 22 409 23
rect 403 20 405 22
rect 407 20 409 22
rect 403 13 409 20
rect 424 13 428 27
rect 434 29 438 35
rect 434 27 435 29
rect 437 27 438 29
rect 434 25 438 27
rect 462 55 466 67
rect 462 53 463 55
rect 465 53 466 55
rect 480 57 484 69
rect 518 63 522 69
rect 518 61 519 63
rect 521 61 522 63
rect 518 59 522 61
rect 530 63 540 64
rect 530 61 536 63
rect 538 61 540 63
rect 530 60 540 61
rect 551 61 557 69
rect 480 55 481 57
rect 483 55 484 57
rect 480 53 484 55
rect 487 57 503 58
rect 487 55 499 57
rect 501 55 503 57
rect 487 54 503 55
rect 508 57 512 59
rect 508 55 509 57
rect 511 55 512 57
rect 462 51 466 53
rect 470 47 477 48
rect 470 45 473 47
rect 475 45 477 47
rect 470 44 477 45
rect 470 38 474 44
rect 487 39 491 54
rect 508 48 512 55
rect 494 47 503 48
rect 494 45 496 47
rect 498 45 503 47
rect 494 44 503 45
rect 458 37 474 38
rect 458 35 460 37
rect 462 35 474 37
rect 477 38 493 39
rect 477 36 479 38
rect 481 36 493 38
rect 477 35 493 36
rect 458 34 474 35
rect 470 29 474 34
rect 470 27 471 29
rect 473 27 474 29
rect 470 25 474 27
rect 481 22 485 24
rect 462 19 466 21
rect 462 17 463 19
rect 465 17 466 19
rect 462 13 466 17
rect 481 20 482 22
rect 484 20 485 22
rect 481 13 485 20
rect 489 23 493 35
rect 499 33 503 44
rect 508 47 526 48
rect 508 45 522 47
rect 524 45 526 47
rect 508 44 526 45
rect 499 31 505 33
rect 499 29 502 31
rect 504 29 505 31
rect 499 27 505 29
rect 489 22 503 23
rect 489 20 499 22
rect 501 20 503 22
rect 489 19 503 20
rect 508 22 512 44
rect 530 41 534 60
rect 551 59 553 61
rect 555 59 557 61
rect 571 62 577 69
rect 571 60 573 62
rect 575 60 577 62
rect 610 67 611 69
rect 613 67 614 69
rect 571 59 577 60
rect 551 58 557 59
rect 582 58 586 60
rect 562 56 566 58
rect 562 55 563 56
rect 525 37 534 41
rect 538 54 563 55
rect 565 54 566 56
rect 582 56 583 58
rect 585 56 586 58
rect 538 51 566 54
rect 538 47 542 51
rect 538 45 539 47
rect 541 45 542 47
rect 525 34 529 37
rect 515 32 529 34
rect 538 33 542 45
rect 582 39 586 56
rect 564 38 586 39
rect 564 36 566 38
rect 568 36 586 38
rect 564 35 586 36
rect 515 30 516 32
rect 518 30 529 32
rect 515 28 529 30
rect 508 20 509 22
rect 511 20 512 22
rect 508 18 512 20
rect 518 22 522 24
rect 518 20 519 22
rect 521 20 522 22
rect 518 13 522 20
rect 525 23 529 28
rect 532 31 542 33
rect 532 29 533 31
rect 535 29 567 31
rect 532 27 563 29
rect 565 27 567 29
rect 561 26 567 27
rect 572 29 576 31
rect 572 27 573 29
rect 575 27 576 29
rect 525 22 540 23
rect 525 20 536 22
rect 538 20 540 22
rect 525 19 540 20
rect 551 22 557 23
rect 551 20 553 22
rect 555 20 557 22
rect 551 13 557 20
rect 572 13 576 27
rect 582 29 586 35
rect 582 27 583 29
rect 585 27 586 29
rect 582 25 586 27
rect 610 55 614 67
rect 610 53 611 55
rect 613 53 614 55
rect 628 57 632 69
rect 666 63 670 69
rect 666 61 667 63
rect 669 61 670 63
rect 666 59 670 61
rect 678 63 688 64
rect 678 61 684 63
rect 686 61 688 63
rect 678 60 688 61
rect 699 61 705 69
rect 628 55 629 57
rect 631 55 632 57
rect 628 53 632 55
rect 635 57 651 58
rect 635 55 647 57
rect 649 55 651 57
rect 635 54 651 55
rect 656 57 660 59
rect 656 55 657 57
rect 659 55 660 57
rect 610 51 614 53
rect 618 47 625 48
rect 618 45 621 47
rect 623 45 625 47
rect 618 44 625 45
rect 618 38 622 44
rect 635 39 639 54
rect 656 48 660 55
rect 642 47 651 48
rect 642 45 644 47
rect 646 45 651 47
rect 642 44 651 45
rect 606 37 622 38
rect 606 35 608 37
rect 610 35 622 37
rect 625 38 641 39
rect 625 36 627 38
rect 629 36 641 38
rect 625 35 641 36
rect 606 34 622 35
rect 618 29 622 34
rect 618 27 619 29
rect 621 27 622 29
rect 618 25 622 27
rect 629 22 633 24
rect 610 19 614 21
rect 610 17 611 19
rect 613 17 614 19
rect 610 13 614 17
rect 629 20 630 22
rect 632 20 633 22
rect 629 13 633 20
rect 637 23 641 35
rect 647 33 651 44
rect 656 47 674 48
rect 656 45 670 47
rect 672 45 674 47
rect 656 44 674 45
rect 647 31 653 33
rect 647 29 650 31
rect 652 29 653 31
rect 647 27 653 29
rect 637 22 651 23
rect 637 20 647 22
rect 649 20 651 22
rect 637 19 651 20
rect 656 22 660 44
rect 678 41 682 60
rect 699 59 701 61
rect 703 59 705 61
rect 719 62 725 69
rect 719 60 721 62
rect 723 60 725 62
rect 758 67 759 69
rect 761 67 762 69
rect 719 59 725 60
rect 699 58 705 59
rect 730 58 734 60
rect 710 56 714 58
rect 710 55 711 56
rect 673 37 682 41
rect 686 54 711 55
rect 713 54 714 56
rect 730 56 731 58
rect 733 56 734 58
rect 686 51 714 54
rect 686 47 690 51
rect 686 45 687 47
rect 689 45 690 47
rect 673 34 677 37
rect 663 32 677 34
rect 686 33 690 45
rect 730 39 734 56
rect 712 38 734 39
rect 712 36 714 38
rect 716 36 734 38
rect 712 35 734 36
rect 663 30 664 32
rect 666 30 677 32
rect 663 28 677 30
rect 656 20 657 22
rect 659 20 660 22
rect 656 18 660 20
rect 666 22 670 24
rect 666 20 667 22
rect 669 20 670 22
rect 666 13 670 20
rect 673 23 677 28
rect 680 31 690 33
rect 680 29 681 31
rect 683 29 715 31
rect 680 27 711 29
rect 713 27 715 29
rect 709 26 715 27
rect 720 29 724 31
rect 720 27 721 29
rect 723 27 724 29
rect 673 22 688 23
rect 673 20 684 22
rect 686 20 688 22
rect 673 19 688 20
rect 699 22 705 23
rect 699 20 701 22
rect 703 20 705 22
rect 699 13 705 20
rect 720 13 724 27
rect 730 29 734 35
rect 730 27 731 29
rect 733 27 734 29
rect 730 25 734 27
rect 758 55 762 67
rect 758 53 759 55
rect 761 53 762 55
rect 776 57 780 69
rect 814 63 818 69
rect 814 61 815 63
rect 817 61 818 63
rect 814 59 818 61
rect 826 63 836 64
rect 826 61 832 63
rect 834 61 836 63
rect 826 60 836 61
rect 847 61 853 69
rect 776 55 777 57
rect 779 55 780 57
rect 776 53 780 55
rect 783 57 799 58
rect 783 55 795 57
rect 797 55 799 57
rect 783 54 799 55
rect 804 57 808 59
rect 804 55 805 57
rect 807 55 808 57
rect 758 51 762 53
rect 766 47 773 48
rect 766 45 769 47
rect 771 45 773 47
rect 766 44 773 45
rect 766 38 770 44
rect 783 39 787 54
rect 804 48 808 55
rect 790 47 799 48
rect 790 45 792 47
rect 794 45 799 47
rect 790 44 799 45
rect 754 37 770 38
rect 754 35 756 37
rect 758 35 770 37
rect 773 38 789 39
rect 773 36 775 38
rect 777 36 789 38
rect 773 35 789 36
rect 754 34 770 35
rect 766 29 770 34
rect 766 27 767 29
rect 769 27 770 29
rect 766 25 770 27
rect 777 22 781 24
rect 758 19 762 21
rect 758 17 759 19
rect 761 17 762 19
rect 758 13 762 17
rect 777 20 778 22
rect 780 20 781 22
rect 777 13 781 20
rect 785 23 789 35
rect 795 33 799 44
rect 804 47 822 48
rect 804 45 818 47
rect 820 45 822 47
rect 804 44 822 45
rect 795 31 801 33
rect 795 29 798 31
rect 800 29 801 31
rect 795 27 801 29
rect 785 22 799 23
rect 785 20 795 22
rect 797 20 799 22
rect 785 19 799 20
rect 804 22 808 44
rect 826 41 830 60
rect 847 59 849 61
rect 851 59 853 61
rect 867 62 873 69
rect 867 60 869 62
rect 871 60 873 62
rect 906 67 907 69
rect 909 67 910 69
rect 867 59 873 60
rect 847 58 853 59
rect 878 58 882 60
rect 858 56 862 58
rect 858 55 859 56
rect 821 37 830 41
rect 834 54 859 55
rect 861 54 862 56
rect 878 56 879 58
rect 881 56 882 58
rect 834 51 862 54
rect 834 47 838 51
rect 834 45 835 47
rect 837 45 838 47
rect 821 34 825 37
rect 811 32 825 34
rect 834 33 838 45
rect 878 39 882 56
rect 860 38 882 39
rect 860 36 862 38
rect 864 36 882 38
rect 860 35 882 36
rect 811 30 812 32
rect 814 30 825 32
rect 811 28 825 30
rect 804 20 805 22
rect 807 20 808 22
rect 804 18 808 20
rect 814 22 818 24
rect 814 20 815 22
rect 817 20 818 22
rect 814 13 818 20
rect 821 23 825 28
rect 828 31 838 33
rect 828 29 829 31
rect 831 29 863 31
rect 828 27 859 29
rect 861 27 863 29
rect 857 26 863 27
rect 868 29 872 31
rect 868 27 869 29
rect 871 27 872 29
rect 821 22 836 23
rect 821 20 832 22
rect 834 20 836 22
rect 821 19 836 20
rect 847 22 853 23
rect 847 20 849 22
rect 851 20 853 22
rect 847 13 853 20
rect 868 13 872 27
rect 878 29 882 35
rect 878 27 879 29
rect 881 27 882 29
rect 878 25 882 27
rect 906 55 910 67
rect 906 53 907 55
rect 909 53 910 55
rect 924 57 928 69
rect 962 63 966 69
rect 962 61 963 63
rect 965 61 966 63
rect 962 59 966 61
rect 974 63 984 64
rect 974 61 980 63
rect 982 61 984 63
rect 974 60 984 61
rect 995 61 1001 69
rect 924 55 925 57
rect 927 55 928 57
rect 924 53 928 55
rect 931 57 947 58
rect 931 55 943 57
rect 945 55 947 57
rect 931 54 947 55
rect 952 57 956 59
rect 952 55 953 57
rect 955 55 956 57
rect 906 51 910 53
rect 914 47 921 48
rect 914 45 917 47
rect 919 45 921 47
rect 914 44 921 45
rect 914 38 918 44
rect 931 39 935 54
rect 952 48 956 55
rect 938 47 947 48
rect 938 45 940 47
rect 942 45 947 47
rect 938 44 947 45
rect 902 37 918 38
rect 902 35 904 37
rect 906 35 918 37
rect 921 38 937 39
rect 921 36 923 38
rect 925 36 937 38
rect 921 35 937 36
rect 902 34 918 35
rect 914 29 918 34
rect 914 27 915 29
rect 917 27 918 29
rect 914 25 918 27
rect 925 22 929 24
rect 906 19 910 21
rect 906 17 907 19
rect 909 17 910 19
rect 906 13 910 17
rect 925 20 926 22
rect 928 20 929 22
rect 925 13 929 20
rect 933 23 937 35
rect 943 33 947 44
rect 952 47 970 48
rect 952 45 966 47
rect 968 45 970 47
rect 952 44 970 45
rect 943 31 949 33
rect 943 29 946 31
rect 948 29 949 31
rect 943 27 949 29
rect 933 22 947 23
rect 933 20 943 22
rect 945 20 947 22
rect 933 19 947 20
rect 952 22 956 44
rect 974 41 978 60
rect 995 59 997 61
rect 999 59 1001 61
rect 1015 62 1021 69
rect 1015 60 1017 62
rect 1019 60 1021 62
rect 1054 67 1055 69
rect 1057 67 1058 69
rect 1015 59 1021 60
rect 995 58 1001 59
rect 1026 58 1030 60
rect 1006 56 1010 58
rect 1006 55 1007 56
rect 969 37 978 41
rect 982 54 1007 55
rect 1009 54 1010 56
rect 1026 56 1027 58
rect 1029 56 1030 58
rect 982 51 1010 54
rect 982 47 986 51
rect 982 45 983 47
rect 985 45 986 47
rect 969 34 973 37
rect 959 32 973 34
rect 982 33 986 45
rect 1026 39 1030 56
rect 1008 38 1030 39
rect 1008 36 1010 38
rect 1012 36 1030 38
rect 1008 35 1030 36
rect 959 30 960 32
rect 962 30 973 32
rect 959 28 973 30
rect 952 20 953 22
rect 955 20 956 22
rect 952 18 956 20
rect 962 22 966 24
rect 962 20 963 22
rect 965 20 966 22
rect 962 13 966 20
rect 969 23 973 28
rect 976 31 986 33
rect 976 29 977 31
rect 979 29 1011 31
rect 976 27 1007 29
rect 1009 27 1011 29
rect 1005 26 1011 27
rect 1016 29 1020 31
rect 1016 27 1017 29
rect 1019 27 1020 29
rect 969 22 984 23
rect 969 20 980 22
rect 982 20 984 22
rect 969 19 984 20
rect 995 22 1001 23
rect 995 20 997 22
rect 999 20 1001 22
rect 995 13 1001 20
rect 1016 13 1020 27
rect 1026 29 1030 35
rect 1026 27 1027 29
rect 1029 27 1030 29
rect 1026 25 1030 27
rect 1054 55 1058 67
rect 1054 53 1055 55
rect 1057 53 1058 55
rect 1072 57 1076 69
rect 1110 63 1114 69
rect 1110 61 1111 63
rect 1113 61 1114 63
rect 1110 59 1114 61
rect 1122 63 1132 64
rect 1122 61 1128 63
rect 1130 61 1132 63
rect 1122 60 1132 61
rect 1143 61 1149 69
rect 1072 55 1073 57
rect 1075 55 1076 57
rect 1072 53 1076 55
rect 1079 57 1095 58
rect 1079 55 1091 57
rect 1093 55 1095 57
rect 1079 54 1095 55
rect 1100 57 1104 59
rect 1100 55 1101 57
rect 1103 55 1104 57
rect 1054 51 1058 53
rect 1062 47 1069 48
rect 1062 45 1065 47
rect 1067 45 1069 47
rect 1062 44 1069 45
rect 1062 38 1066 44
rect 1079 39 1083 54
rect 1100 48 1104 55
rect 1086 47 1095 48
rect 1086 45 1088 47
rect 1090 45 1095 47
rect 1086 44 1095 45
rect 1050 37 1066 38
rect 1050 35 1052 37
rect 1054 35 1066 37
rect 1069 38 1085 39
rect 1069 36 1071 38
rect 1073 36 1085 38
rect 1069 35 1085 36
rect 1050 34 1066 35
rect 1062 29 1066 34
rect 1062 27 1063 29
rect 1065 27 1066 29
rect 1062 25 1066 27
rect 1073 22 1077 24
rect 1054 19 1058 21
rect 1054 17 1055 19
rect 1057 17 1058 19
rect 1054 13 1058 17
rect 1073 20 1074 22
rect 1076 20 1077 22
rect 1073 13 1077 20
rect 1081 23 1085 35
rect 1091 33 1095 44
rect 1100 47 1118 48
rect 1100 45 1114 47
rect 1116 45 1118 47
rect 1100 44 1118 45
rect 1091 31 1097 33
rect 1091 29 1094 31
rect 1096 29 1097 31
rect 1091 27 1097 29
rect 1081 22 1095 23
rect 1081 20 1091 22
rect 1093 20 1095 22
rect 1081 19 1095 20
rect 1100 22 1104 44
rect 1122 41 1126 60
rect 1143 59 1145 61
rect 1147 59 1149 61
rect 1163 62 1169 69
rect 1163 60 1165 62
rect 1167 60 1169 62
rect 1163 59 1169 60
rect 1143 58 1149 59
rect 1174 58 1178 60
rect 1154 56 1158 58
rect 1154 55 1155 56
rect 1117 37 1126 41
rect 1130 54 1155 55
rect 1157 54 1158 56
rect 1174 56 1175 58
rect 1177 56 1178 58
rect 1130 51 1158 54
rect 1130 47 1134 51
rect 1130 45 1131 47
rect 1133 45 1134 47
rect 1117 34 1121 37
rect 1107 32 1121 34
rect 1130 33 1134 45
rect 1174 39 1178 56
rect 1156 38 1178 39
rect 1156 36 1158 38
rect 1160 36 1178 38
rect 1156 35 1178 36
rect 1107 30 1108 32
rect 1110 30 1121 32
rect 1107 28 1121 30
rect 1100 20 1101 22
rect 1103 20 1104 22
rect 1100 18 1104 20
rect 1110 22 1114 24
rect 1110 20 1111 22
rect 1113 20 1114 22
rect 1110 13 1114 20
rect 1117 23 1121 28
rect 1124 31 1134 33
rect 1124 29 1125 31
rect 1127 29 1159 31
rect 1124 27 1155 29
rect 1157 27 1159 29
rect 1153 26 1159 27
rect 1164 29 1168 31
rect 1164 27 1165 29
rect 1167 27 1168 29
rect 1117 22 1132 23
rect 1117 20 1128 22
rect 1130 20 1132 22
rect 1117 19 1132 20
rect 1143 22 1149 23
rect 1143 20 1145 22
rect 1147 20 1149 22
rect 1143 13 1149 20
rect 1164 13 1168 27
rect 1174 29 1178 35
rect 1174 27 1175 29
rect 1177 27 1178 29
rect 1174 25 1178 27
rect 12 -17 16 -15
rect 12 -19 13 -17
rect 15 -19 16 -17
rect 12 -25 16 -19
rect 22 -17 26 -3
rect 41 -10 47 -3
rect 41 -12 43 -10
rect 45 -12 47 -10
rect 41 -13 47 -12
rect 58 -10 73 -9
rect 58 -12 60 -10
rect 62 -12 73 -10
rect 58 -13 73 -12
rect 22 -19 23 -17
rect 25 -19 26 -17
rect 22 -21 26 -19
rect 31 -17 37 -16
rect 31 -19 33 -17
rect 35 -19 66 -17
rect 31 -21 63 -19
rect 65 -21 66 -19
rect 56 -23 66 -21
rect 69 -18 73 -13
rect 76 -10 80 -3
rect 76 -12 77 -10
rect 79 -12 80 -10
rect 76 -14 80 -12
rect 86 -10 90 -8
rect 86 -12 87 -10
rect 89 -12 90 -10
rect 69 -20 83 -18
rect 69 -22 80 -20
rect 82 -22 83 -20
rect 12 -26 34 -25
rect 12 -28 30 -26
rect 32 -28 34 -26
rect 12 -29 34 -28
rect 12 -46 16 -29
rect 56 -35 60 -23
rect 69 -24 83 -22
rect 69 -27 73 -24
rect 56 -37 57 -35
rect 59 -37 60 -35
rect 56 -41 60 -37
rect 32 -44 60 -41
rect 12 -48 13 -46
rect 15 -48 16 -46
rect 32 -46 33 -44
rect 35 -45 60 -44
rect 64 -31 73 -27
rect 35 -46 36 -45
rect 32 -48 36 -46
rect 12 -50 16 -48
rect 41 -49 47 -48
rect 21 -50 27 -49
rect 21 -52 23 -50
rect 25 -52 27 -50
rect 21 -59 27 -52
rect 41 -51 43 -49
rect 45 -51 47 -49
rect 64 -50 68 -31
rect 86 -34 90 -12
rect 95 -10 109 -9
rect 95 -12 97 -10
rect 99 -12 109 -10
rect 95 -13 109 -12
rect 93 -19 99 -17
rect 93 -21 94 -19
rect 96 -21 99 -19
rect 93 -23 99 -21
rect 72 -35 90 -34
rect 72 -37 74 -35
rect 76 -37 90 -35
rect 72 -38 90 -37
rect 95 -34 99 -23
rect 105 -25 109 -13
rect 113 -10 117 -3
rect 113 -12 114 -10
rect 116 -12 117 -10
rect 132 -7 136 -3
rect 132 -9 133 -7
rect 135 -9 136 -7
rect 132 -11 136 -9
rect 113 -14 117 -12
rect 124 -17 128 -15
rect 124 -19 125 -17
rect 127 -19 128 -17
rect 124 -24 128 -19
rect 124 -25 140 -24
rect 105 -26 121 -25
rect 105 -28 117 -26
rect 119 -28 121 -26
rect 105 -29 121 -28
rect 124 -27 136 -25
rect 138 -27 140 -25
rect 124 -28 140 -27
rect 95 -35 104 -34
rect 95 -37 100 -35
rect 102 -37 104 -35
rect 95 -38 104 -37
rect 86 -45 90 -38
rect 107 -44 111 -29
rect 124 -34 128 -28
rect 121 -35 128 -34
rect 121 -37 123 -35
rect 125 -37 128 -35
rect 121 -38 128 -37
rect 132 -43 136 -41
rect 86 -47 87 -45
rect 89 -47 90 -45
rect 86 -49 90 -47
rect 95 -45 111 -44
rect 95 -47 97 -45
rect 99 -47 111 -45
rect 95 -48 111 -47
rect 114 -45 118 -43
rect 114 -47 115 -45
rect 117 -47 118 -45
rect 41 -59 47 -51
rect 58 -51 68 -50
rect 58 -53 60 -51
rect 62 -53 68 -51
rect 58 -54 68 -53
rect 76 -51 80 -49
rect 76 -53 77 -51
rect 79 -53 80 -51
rect 76 -59 80 -53
rect 114 -59 118 -47
rect 132 -45 133 -43
rect 135 -45 136 -43
rect 132 -57 136 -45
rect 160 -17 164 -15
rect 160 -19 161 -17
rect 163 -19 164 -17
rect 160 -25 164 -19
rect 170 -17 174 -3
rect 189 -10 195 -3
rect 189 -12 191 -10
rect 193 -12 195 -10
rect 189 -13 195 -12
rect 206 -10 221 -9
rect 206 -12 208 -10
rect 210 -12 221 -10
rect 206 -13 221 -12
rect 170 -19 171 -17
rect 173 -19 174 -17
rect 170 -21 174 -19
rect 179 -17 185 -16
rect 179 -19 181 -17
rect 183 -19 214 -17
rect 179 -21 211 -19
rect 213 -21 214 -19
rect 204 -23 214 -21
rect 217 -18 221 -13
rect 224 -10 228 -3
rect 224 -12 225 -10
rect 227 -12 228 -10
rect 224 -14 228 -12
rect 234 -10 238 -8
rect 234 -12 235 -10
rect 237 -12 238 -10
rect 217 -20 231 -18
rect 217 -22 228 -20
rect 230 -22 231 -20
rect 160 -26 182 -25
rect 160 -28 178 -26
rect 180 -28 182 -26
rect 160 -29 182 -28
rect 160 -46 164 -29
rect 204 -35 208 -23
rect 217 -24 231 -22
rect 217 -27 221 -24
rect 204 -37 205 -35
rect 207 -37 208 -35
rect 204 -41 208 -37
rect 180 -44 208 -41
rect 160 -48 161 -46
rect 163 -48 164 -46
rect 180 -46 181 -44
rect 183 -45 208 -44
rect 212 -31 221 -27
rect 183 -46 184 -45
rect 180 -48 184 -46
rect 160 -50 164 -48
rect 189 -49 195 -48
rect 169 -50 175 -49
rect 132 -59 133 -57
rect 135 -59 136 -57
rect 169 -52 171 -50
rect 173 -52 175 -50
rect 169 -59 175 -52
rect 189 -51 191 -49
rect 193 -51 195 -49
rect 212 -50 216 -31
rect 234 -34 238 -12
rect 243 -10 257 -9
rect 243 -12 245 -10
rect 247 -12 257 -10
rect 243 -13 257 -12
rect 241 -19 247 -17
rect 241 -21 242 -19
rect 244 -21 247 -19
rect 241 -23 247 -21
rect 220 -35 238 -34
rect 220 -37 222 -35
rect 224 -37 238 -35
rect 220 -38 238 -37
rect 243 -34 247 -23
rect 253 -25 257 -13
rect 261 -10 265 -3
rect 261 -12 262 -10
rect 264 -12 265 -10
rect 280 -7 284 -3
rect 280 -9 281 -7
rect 283 -9 284 -7
rect 280 -11 284 -9
rect 261 -14 265 -12
rect 272 -17 276 -15
rect 272 -19 273 -17
rect 275 -19 276 -17
rect 272 -24 276 -19
rect 272 -25 288 -24
rect 253 -26 269 -25
rect 253 -28 265 -26
rect 267 -28 269 -26
rect 253 -29 269 -28
rect 272 -27 284 -25
rect 286 -27 288 -25
rect 272 -28 288 -27
rect 243 -35 252 -34
rect 243 -37 248 -35
rect 250 -37 252 -35
rect 243 -38 252 -37
rect 234 -45 238 -38
rect 255 -44 259 -29
rect 272 -34 276 -28
rect 269 -35 276 -34
rect 269 -37 271 -35
rect 273 -37 276 -35
rect 269 -38 276 -37
rect 280 -43 284 -41
rect 234 -47 235 -45
rect 237 -47 238 -45
rect 234 -49 238 -47
rect 243 -45 259 -44
rect 243 -47 245 -45
rect 247 -47 259 -45
rect 243 -48 259 -47
rect 262 -45 266 -43
rect 262 -47 263 -45
rect 265 -47 266 -45
rect 189 -59 195 -51
rect 206 -51 216 -50
rect 206 -53 208 -51
rect 210 -53 216 -51
rect 206 -54 216 -53
rect 224 -51 228 -49
rect 224 -53 225 -51
rect 227 -53 228 -51
rect 224 -59 228 -53
rect 262 -59 266 -47
rect 280 -45 281 -43
rect 283 -45 284 -43
rect 280 -57 284 -45
rect 308 -17 312 -15
rect 308 -19 309 -17
rect 311 -19 312 -17
rect 308 -25 312 -19
rect 318 -17 322 -3
rect 337 -10 343 -3
rect 337 -12 339 -10
rect 341 -12 343 -10
rect 337 -13 343 -12
rect 354 -10 369 -9
rect 354 -12 356 -10
rect 358 -12 369 -10
rect 354 -13 369 -12
rect 318 -19 319 -17
rect 321 -19 322 -17
rect 318 -21 322 -19
rect 327 -17 333 -16
rect 327 -19 329 -17
rect 331 -19 362 -17
rect 327 -21 359 -19
rect 361 -21 362 -19
rect 352 -23 362 -21
rect 365 -18 369 -13
rect 372 -10 376 -3
rect 372 -12 373 -10
rect 375 -12 376 -10
rect 372 -14 376 -12
rect 382 -10 386 -8
rect 382 -12 383 -10
rect 385 -12 386 -10
rect 365 -20 379 -18
rect 365 -22 376 -20
rect 378 -22 379 -20
rect 308 -26 330 -25
rect 308 -28 326 -26
rect 328 -28 330 -26
rect 308 -29 330 -28
rect 308 -46 312 -29
rect 352 -35 356 -23
rect 365 -24 379 -22
rect 365 -27 369 -24
rect 352 -37 353 -35
rect 355 -37 356 -35
rect 352 -41 356 -37
rect 328 -44 356 -41
rect 308 -48 309 -46
rect 311 -48 312 -46
rect 328 -46 329 -44
rect 331 -45 356 -44
rect 360 -31 369 -27
rect 331 -46 332 -45
rect 328 -48 332 -46
rect 308 -50 312 -48
rect 337 -49 343 -48
rect 317 -50 323 -49
rect 280 -59 281 -57
rect 283 -59 284 -57
rect 317 -52 319 -50
rect 321 -52 323 -50
rect 317 -59 323 -52
rect 337 -51 339 -49
rect 341 -51 343 -49
rect 360 -50 364 -31
rect 382 -34 386 -12
rect 391 -10 405 -9
rect 391 -12 393 -10
rect 395 -12 405 -10
rect 391 -13 405 -12
rect 389 -19 395 -17
rect 389 -21 390 -19
rect 392 -21 395 -19
rect 389 -23 395 -21
rect 368 -35 386 -34
rect 368 -37 370 -35
rect 372 -37 386 -35
rect 368 -38 386 -37
rect 391 -34 395 -23
rect 401 -25 405 -13
rect 409 -10 413 -3
rect 409 -12 410 -10
rect 412 -12 413 -10
rect 428 -7 432 -3
rect 428 -9 429 -7
rect 431 -9 432 -7
rect 428 -11 432 -9
rect 409 -14 413 -12
rect 420 -17 424 -15
rect 420 -19 421 -17
rect 423 -19 424 -17
rect 420 -24 424 -19
rect 420 -25 436 -24
rect 401 -26 417 -25
rect 401 -28 413 -26
rect 415 -28 417 -26
rect 401 -29 417 -28
rect 420 -27 432 -25
rect 434 -27 436 -25
rect 420 -28 436 -27
rect 391 -35 400 -34
rect 391 -37 396 -35
rect 398 -37 400 -35
rect 391 -38 400 -37
rect 382 -45 386 -38
rect 403 -44 407 -29
rect 420 -34 424 -28
rect 417 -35 424 -34
rect 417 -37 419 -35
rect 421 -37 424 -35
rect 417 -38 424 -37
rect 428 -43 432 -41
rect 382 -47 383 -45
rect 385 -47 386 -45
rect 382 -49 386 -47
rect 391 -45 407 -44
rect 391 -47 393 -45
rect 395 -47 407 -45
rect 391 -48 407 -47
rect 410 -45 414 -43
rect 410 -47 411 -45
rect 413 -47 414 -45
rect 337 -59 343 -51
rect 354 -51 364 -50
rect 354 -53 356 -51
rect 358 -53 364 -51
rect 354 -54 364 -53
rect 372 -51 376 -49
rect 372 -53 373 -51
rect 375 -53 376 -51
rect 372 -59 376 -53
rect 410 -59 414 -47
rect 428 -45 429 -43
rect 431 -45 432 -43
rect 428 -57 432 -45
rect 456 -17 460 -15
rect 456 -19 457 -17
rect 459 -19 460 -17
rect 456 -25 460 -19
rect 466 -17 470 -3
rect 485 -10 491 -3
rect 485 -12 487 -10
rect 489 -12 491 -10
rect 485 -13 491 -12
rect 502 -10 517 -9
rect 502 -12 504 -10
rect 506 -12 517 -10
rect 502 -13 517 -12
rect 466 -19 467 -17
rect 469 -19 470 -17
rect 466 -21 470 -19
rect 475 -17 481 -16
rect 475 -19 477 -17
rect 479 -19 510 -17
rect 475 -21 507 -19
rect 509 -21 510 -19
rect 500 -23 510 -21
rect 513 -18 517 -13
rect 520 -10 524 -3
rect 520 -12 521 -10
rect 523 -12 524 -10
rect 520 -14 524 -12
rect 530 -10 534 -8
rect 530 -12 531 -10
rect 533 -12 534 -10
rect 513 -20 527 -18
rect 513 -22 524 -20
rect 526 -22 527 -20
rect 456 -26 478 -25
rect 456 -28 474 -26
rect 476 -28 478 -26
rect 456 -29 478 -28
rect 456 -46 460 -29
rect 500 -35 504 -23
rect 513 -24 527 -22
rect 513 -27 517 -24
rect 500 -37 501 -35
rect 503 -37 504 -35
rect 500 -41 504 -37
rect 476 -44 504 -41
rect 456 -48 457 -46
rect 459 -48 460 -46
rect 476 -46 477 -44
rect 479 -45 504 -44
rect 508 -31 517 -27
rect 479 -46 480 -45
rect 476 -48 480 -46
rect 456 -50 460 -48
rect 485 -49 491 -48
rect 465 -50 471 -49
rect 428 -59 429 -57
rect 431 -59 432 -57
rect 465 -52 467 -50
rect 469 -52 471 -50
rect 465 -59 471 -52
rect 485 -51 487 -49
rect 489 -51 491 -49
rect 508 -50 512 -31
rect 530 -34 534 -12
rect 539 -10 553 -9
rect 539 -12 541 -10
rect 543 -12 553 -10
rect 539 -13 553 -12
rect 537 -19 543 -17
rect 537 -21 538 -19
rect 540 -21 543 -19
rect 537 -23 543 -21
rect 516 -35 534 -34
rect 516 -37 518 -35
rect 520 -37 534 -35
rect 516 -38 534 -37
rect 539 -34 543 -23
rect 549 -25 553 -13
rect 557 -10 561 -3
rect 557 -12 558 -10
rect 560 -12 561 -10
rect 576 -7 580 -3
rect 576 -9 577 -7
rect 579 -9 580 -7
rect 576 -11 580 -9
rect 557 -14 561 -12
rect 568 -17 572 -15
rect 568 -19 569 -17
rect 571 -19 572 -17
rect 568 -24 572 -19
rect 568 -25 584 -24
rect 549 -26 565 -25
rect 549 -28 561 -26
rect 563 -28 565 -26
rect 549 -29 565 -28
rect 568 -27 580 -25
rect 582 -27 584 -25
rect 568 -28 584 -27
rect 539 -35 548 -34
rect 539 -37 544 -35
rect 546 -37 548 -35
rect 539 -38 548 -37
rect 530 -45 534 -38
rect 551 -44 555 -29
rect 568 -34 572 -28
rect 565 -35 572 -34
rect 565 -37 567 -35
rect 569 -37 572 -35
rect 565 -38 572 -37
rect 576 -43 580 -41
rect 530 -47 531 -45
rect 533 -47 534 -45
rect 530 -49 534 -47
rect 539 -45 555 -44
rect 539 -47 541 -45
rect 543 -47 555 -45
rect 539 -48 555 -47
rect 558 -45 562 -43
rect 558 -47 559 -45
rect 561 -47 562 -45
rect 485 -59 491 -51
rect 502 -51 512 -50
rect 502 -53 504 -51
rect 506 -53 512 -51
rect 502 -54 512 -53
rect 520 -51 524 -49
rect 520 -53 521 -51
rect 523 -53 524 -51
rect 520 -59 524 -53
rect 558 -59 562 -47
rect 576 -45 577 -43
rect 579 -45 580 -43
rect 576 -57 580 -45
rect 604 -17 608 -15
rect 604 -19 605 -17
rect 607 -19 608 -17
rect 604 -25 608 -19
rect 614 -17 618 -3
rect 633 -10 639 -3
rect 633 -12 635 -10
rect 637 -12 639 -10
rect 633 -13 639 -12
rect 650 -10 665 -9
rect 650 -12 652 -10
rect 654 -12 665 -10
rect 650 -13 665 -12
rect 614 -19 615 -17
rect 617 -19 618 -17
rect 614 -21 618 -19
rect 623 -17 629 -16
rect 623 -19 625 -17
rect 627 -19 658 -17
rect 623 -21 655 -19
rect 657 -21 658 -19
rect 648 -23 658 -21
rect 661 -18 665 -13
rect 668 -10 672 -3
rect 668 -12 669 -10
rect 671 -12 672 -10
rect 668 -14 672 -12
rect 678 -10 682 -8
rect 678 -12 679 -10
rect 681 -12 682 -10
rect 661 -20 675 -18
rect 661 -22 672 -20
rect 674 -22 675 -20
rect 604 -26 626 -25
rect 604 -28 622 -26
rect 624 -28 626 -26
rect 604 -29 626 -28
rect 604 -46 608 -29
rect 648 -35 652 -23
rect 661 -24 675 -22
rect 661 -27 665 -24
rect 648 -37 649 -35
rect 651 -37 652 -35
rect 648 -41 652 -37
rect 624 -44 652 -41
rect 604 -48 605 -46
rect 607 -48 608 -46
rect 624 -46 625 -44
rect 627 -45 652 -44
rect 656 -31 665 -27
rect 627 -46 628 -45
rect 624 -48 628 -46
rect 604 -50 608 -48
rect 633 -49 639 -48
rect 613 -50 619 -49
rect 576 -59 577 -57
rect 579 -59 580 -57
rect 613 -52 615 -50
rect 617 -52 619 -50
rect 613 -59 619 -52
rect 633 -51 635 -49
rect 637 -51 639 -49
rect 656 -50 660 -31
rect 678 -34 682 -12
rect 687 -10 701 -9
rect 687 -12 689 -10
rect 691 -12 701 -10
rect 687 -13 701 -12
rect 685 -19 691 -17
rect 685 -21 686 -19
rect 688 -21 691 -19
rect 685 -23 691 -21
rect 664 -35 682 -34
rect 664 -37 666 -35
rect 668 -37 682 -35
rect 664 -38 682 -37
rect 687 -34 691 -23
rect 697 -25 701 -13
rect 705 -10 709 -3
rect 705 -12 706 -10
rect 708 -12 709 -10
rect 724 -7 728 -3
rect 724 -9 725 -7
rect 727 -9 728 -7
rect 724 -11 728 -9
rect 705 -14 709 -12
rect 716 -17 720 -15
rect 716 -19 717 -17
rect 719 -19 720 -17
rect 716 -24 720 -19
rect 716 -25 732 -24
rect 697 -26 713 -25
rect 697 -28 709 -26
rect 711 -28 713 -26
rect 697 -29 713 -28
rect 716 -27 728 -25
rect 730 -27 732 -25
rect 716 -28 732 -27
rect 687 -35 696 -34
rect 687 -37 692 -35
rect 694 -37 696 -35
rect 687 -38 696 -37
rect 678 -45 682 -38
rect 699 -44 703 -29
rect 716 -34 720 -28
rect 713 -35 720 -34
rect 713 -37 715 -35
rect 717 -37 720 -35
rect 713 -38 720 -37
rect 724 -43 728 -41
rect 678 -47 679 -45
rect 681 -47 682 -45
rect 678 -49 682 -47
rect 687 -45 703 -44
rect 687 -47 689 -45
rect 691 -47 703 -45
rect 687 -48 703 -47
rect 706 -45 710 -43
rect 706 -47 707 -45
rect 709 -47 710 -45
rect 633 -59 639 -51
rect 650 -51 660 -50
rect 650 -53 652 -51
rect 654 -53 660 -51
rect 650 -54 660 -53
rect 668 -51 672 -49
rect 668 -53 669 -51
rect 671 -53 672 -51
rect 668 -59 672 -53
rect 706 -59 710 -47
rect 724 -45 725 -43
rect 727 -45 728 -43
rect 724 -57 728 -45
rect 752 -17 756 -15
rect 752 -19 753 -17
rect 755 -19 756 -17
rect 752 -25 756 -19
rect 762 -17 766 -3
rect 781 -10 787 -3
rect 781 -12 783 -10
rect 785 -12 787 -10
rect 781 -13 787 -12
rect 798 -10 813 -9
rect 798 -12 800 -10
rect 802 -12 813 -10
rect 798 -13 813 -12
rect 762 -19 763 -17
rect 765 -19 766 -17
rect 762 -21 766 -19
rect 771 -17 777 -16
rect 771 -19 773 -17
rect 775 -19 806 -17
rect 771 -21 803 -19
rect 805 -21 806 -19
rect 796 -23 806 -21
rect 809 -18 813 -13
rect 816 -10 820 -3
rect 816 -12 817 -10
rect 819 -12 820 -10
rect 816 -14 820 -12
rect 826 -10 830 -8
rect 826 -12 827 -10
rect 829 -12 830 -10
rect 809 -20 823 -18
rect 809 -22 820 -20
rect 822 -22 823 -20
rect 752 -26 774 -25
rect 752 -28 770 -26
rect 772 -28 774 -26
rect 752 -29 774 -28
rect 752 -46 756 -29
rect 796 -35 800 -23
rect 809 -24 823 -22
rect 809 -27 813 -24
rect 796 -37 797 -35
rect 799 -37 800 -35
rect 796 -41 800 -37
rect 772 -44 800 -41
rect 752 -48 753 -46
rect 755 -48 756 -46
rect 772 -46 773 -44
rect 775 -45 800 -44
rect 804 -31 813 -27
rect 775 -46 776 -45
rect 772 -48 776 -46
rect 752 -50 756 -48
rect 781 -49 787 -48
rect 761 -50 767 -49
rect 724 -59 725 -57
rect 727 -59 728 -57
rect 761 -52 763 -50
rect 765 -52 767 -50
rect 761 -59 767 -52
rect 781 -51 783 -49
rect 785 -51 787 -49
rect 804 -50 808 -31
rect 826 -34 830 -12
rect 835 -10 849 -9
rect 835 -12 837 -10
rect 839 -12 849 -10
rect 835 -13 849 -12
rect 833 -19 839 -17
rect 833 -21 834 -19
rect 836 -21 839 -19
rect 833 -23 839 -21
rect 812 -35 830 -34
rect 812 -37 814 -35
rect 816 -37 830 -35
rect 812 -38 830 -37
rect 835 -34 839 -23
rect 845 -25 849 -13
rect 853 -10 857 -3
rect 853 -12 854 -10
rect 856 -12 857 -10
rect 872 -7 876 -3
rect 872 -9 873 -7
rect 875 -9 876 -7
rect 872 -11 876 -9
rect 853 -14 857 -12
rect 864 -17 868 -15
rect 864 -19 865 -17
rect 867 -19 868 -17
rect 864 -24 868 -19
rect 864 -25 880 -24
rect 845 -26 861 -25
rect 845 -28 857 -26
rect 859 -28 861 -26
rect 845 -29 861 -28
rect 864 -27 876 -25
rect 878 -27 880 -25
rect 864 -28 880 -27
rect 835 -35 844 -34
rect 835 -37 840 -35
rect 842 -37 844 -35
rect 835 -38 844 -37
rect 826 -45 830 -38
rect 847 -44 851 -29
rect 864 -34 868 -28
rect 861 -35 868 -34
rect 861 -37 863 -35
rect 865 -37 868 -35
rect 861 -38 868 -37
rect 872 -43 876 -41
rect 826 -47 827 -45
rect 829 -47 830 -45
rect 826 -49 830 -47
rect 835 -45 851 -44
rect 835 -47 837 -45
rect 839 -47 851 -45
rect 835 -48 851 -47
rect 854 -45 858 -43
rect 854 -47 855 -45
rect 857 -47 858 -45
rect 781 -59 787 -51
rect 798 -51 808 -50
rect 798 -53 800 -51
rect 802 -53 808 -51
rect 798 -54 808 -53
rect 816 -51 820 -49
rect 816 -53 817 -51
rect 819 -53 820 -51
rect 816 -59 820 -53
rect 854 -59 858 -47
rect 872 -45 873 -43
rect 875 -45 876 -43
rect 872 -57 876 -45
rect 900 -17 904 -15
rect 900 -19 901 -17
rect 903 -19 904 -17
rect 900 -25 904 -19
rect 910 -17 914 -3
rect 929 -10 935 -3
rect 929 -12 931 -10
rect 933 -12 935 -10
rect 929 -13 935 -12
rect 946 -10 961 -9
rect 946 -12 948 -10
rect 950 -12 961 -10
rect 946 -13 961 -12
rect 910 -19 911 -17
rect 913 -19 914 -17
rect 910 -21 914 -19
rect 919 -17 925 -16
rect 919 -19 921 -17
rect 923 -19 954 -17
rect 919 -21 951 -19
rect 953 -21 954 -19
rect 944 -23 954 -21
rect 957 -18 961 -13
rect 964 -10 968 -3
rect 964 -12 965 -10
rect 967 -12 968 -10
rect 964 -14 968 -12
rect 974 -10 978 -8
rect 974 -12 975 -10
rect 977 -12 978 -10
rect 957 -20 971 -18
rect 957 -22 968 -20
rect 970 -22 971 -20
rect 900 -26 922 -25
rect 900 -28 918 -26
rect 920 -28 922 -26
rect 900 -29 922 -28
rect 900 -46 904 -29
rect 944 -35 948 -23
rect 957 -24 971 -22
rect 957 -27 961 -24
rect 944 -37 945 -35
rect 947 -37 948 -35
rect 944 -41 948 -37
rect 920 -44 948 -41
rect 900 -48 901 -46
rect 903 -48 904 -46
rect 920 -46 921 -44
rect 923 -45 948 -44
rect 952 -31 961 -27
rect 923 -46 924 -45
rect 920 -48 924 -46
rect 900 -50 904 -48
rect 929 -49 935 -48
rect 909 -50 915 -49
rect 872 -59 873 -57
rect 875 -59 876 -57
rect 909 -52 911 -50
rect 913 -52 915 -50
rect 909 -59 915 -52
rect 929 -51 931 -49
rect 933 -51 935 -49
rect 952 -50 956 -31
rect 974 -34 978 -12
rect 983 -10 997 -9
rect 983 -12 985 -10
rect 987 -12 997 -10
rect 983 -13 997 -12
rect 981 -19 987 -17
rect 981 -21 982 -19
rect 984 -21 987 -19
rect 981 -23 987 -21
rect 960 -35 978 -34
rect 960 -37 962 -35
rect 964 -37 978 -35
rect 960 -38 978 -37
rect 983 -34 987 -23
rect 993 -25 997 -13
rect 1001 -10 1005 -3
rect 1001 -12 1002 -10
rect 1004 -12 1005 -10
rect 1020 -7 1024 -3
rect 1020 -9 1021 -7
rect 1023 -9 1024 -7
rect 1020 -11 1024 -9
rect 1001 -14 1005 -12
rect 1012 -17 1016 -15
rect 1012 -19 1013 -17
rect 1015 -19 1016 -17
rect 1012 -24 1016 -19
rect 1012 -25 1028 -24
rect 993 -26 1009 -25
rect 993 -28 1005 -26
rect 1007 -28 1009 -26
rect 993 -29 1009 -28
rect 1012 -27 1024 -25
rect 1026 -27 1028 -25
rect 1012 -28 1028 -27
rect 983 -35 992 -34
rect 983 -37 988 -35
rect 990 -37 992 -35
rect 983 -38 992 -37
rect 974 -45 978 -38
rect 995 -44 999 -29
rect 1012 -34 1016 -28
rect 1009 -35 1016 -34
rect 1009 -37 1011 -35
rect 1013 -37 1016 -35
rect 1009 -38 1016 -37
rect 1020 -43 1024 -41
rect 974 -47 975 -45
rect 977 -47 978 -45
rect 974 -49 978 -47
rect 983 -45 999 -44
rect 983 -47 985 -45
rect 987 -47 999 -45
rect 983 -48 999 -47
rect 1002 -45 1006 -43
rect 1002 -47 1003 -45
rect 1005 -47 1006 -45
rect 929 -59 935 -51
rect 946 -51 956 -50
rect 946 -53 948 -51
rect 950 -53 956 -51
rect 946 -54 956 -53
rect 964 -51 968 -49
rect 964 -53 965 -51
rect 967 -53 968 -51
rect 964 -59 968 -53
rect 1002 -59 1006 -47
rect 1020 -45 1021 -43
rect 1023 -45 1024 -43
rect 1020 -57 1024 -45
rect 1048 -17 1052 -15
rect 1048 -19 1049 -17
rect 1051 -19 1052 -17
rect 1048 -25 1052 -19
rect 1058 -17 1062 -3
rect 1077 -10 1083 -3
rect 1077 -12 1079 -10
rect 1081 -12 1083 -10
rect 1077 -13 1083 -12
rect 1094 -10 1109 -9
rect 1094 -12 1096 -10
rect 1098 -12 1109 -10
rect 1094 -13 1109 -12
rect 1058 -19 1059 -17
rect 1061 -19 1062 -17
rect 1058 -21 1062 -19
rect 1067 -17 1073 -16
rect 1067 -19 1069 -17
rect 1071 -19 1102 -17
rect 1067 -21 1099 -19
rect 1101 -21 1102 -19
rect 1092 -23 1102 -21
rect 1105 -18 1109 -13
rect 1112 -10 1116 -3
rect 1112 -12 1113 -10
rect 1115 -12 1116 -10
rect 1112 -14 1116 -12
rect 1122 -10 1126 -8
rect 1122 -12 1123 -10
rect 1125 -12 1126 -10
rect 1105 -20 1119 -18
rect 1105 -22 1116 -20
rect 1118 -22 1119 -20
rect 1048 -26 1070 -25
rect 1048 -28 1066 -26
rect 1068 -28 1070 -26
rect 1048 -29 1070 -28
rect 1048 -46 1052 -29
rect 1092 -35 1096 -23
rect 1105 -24 1119 -22
rect 1105 -27 1109 -24
rect 1092 -37 1093 -35
rect 1095 -37 1096 -35
rect 1092 -41 1096 -37
rect 1068 -44 1096 -41
rect 1048 -48 1049 -46
rect 1051 -48 1052 -46
rect 1068 -46 1069 -44
rect 1071 -45 1096 -44
rect 1100 -31 1109 -27
rect 1071 -46 1072 -45
rect 1068 -48 1072 -46
rect 1048 -50 1052 -48
rect 1077 -49 1083 -48
rect 1057 -50 1063 -49
rect 1020 -59 1021 -57
rect 1023 -59 1024 -57
rect 1057 -52 1059 -50
rect 1061 -52 1063 -50
rect 1057 -59 1063 -52
rect 1077 -51 1079 -49
rect 1081 -51 1083 -49
rect 1100 -50 1104 -31
rect 1122 -34 1126 -12
rect 1131 -10 1145 -9
rect 1131 -12 1133 -10
rect 1135 -12 1145 -10
rect 1131 -13 1145 -12
rect 1129 -19 1135 -17
rect 1129 -21 1130 -19
rect 1132 -21 1135 -19
rect 1129 -23 1135 -21
rect 1108 -35 1126 -34
rect 1108 -37 1110 -35
rect 1112 -37 1126 -35
rect 1108 -38 1126 -37
rect 1131 -34 1135 -23
rect 1141 -25 1145 -13
rect 1149 -10 1153 -3
rect 1149 -12 1150 -10
rect 1152 -12 1153 -10
rect 1168 -7 1172 -3
rect 1168 -9 1169 -7
rect 1171 -9 1172 -7
rect 1168 -11 1172 -9
rect 1149 -14 1153 -12
rect 1160 -17 1164 -15
rect 1160 -19 1161 -17
rect 1163 -19 1164 -17
rect 1160 -24 1164 -19
rect 1160 -25 1176 -24
rect 1141 -26 1157 -25
rect 1141 -28 1153 -26
rect 1155 -28 1157 -26
rect 1141 -29 1157 -28
rect 1160 -27 1172 -25
rect 1174 -27 1176 -25
rect 1160 -28 1176 -27
rect 1131 -35 1140 -34
rect 1131 -37 1136 -35
rect 1138 -37 1140 -35
rect 1131 -38 1140 -37
rect 1122 -45 1126 -38
rect 1143 -44 1147 -29
rect 1160 -34 1164 -28
rect 1157 -35 1164 -34
rect 1157 -37 1159 -35
rect 1161 -37 1164 -35
rect 1157 -38 1164 -37
rect 1168 -43 1172 -41
rect 1122 -47 1123 -45
rect 1125 -47 1126 -45
rect 1122 -49 1126 -47
rect 1131 -45 1147 -44
rect 1131 -47 1133 -45
rect 1135 -47 1147 -45
rect 1131 -48 1147 -47
rect 1150 -45 1154 -43
rect 1150 -47 1151 -45
rect 1153 -47 1154 -45
rect 1077 -59 1083 -51
rect 1094 -51 1104 -50
rect 1094 -53 1096 -51
rect 1098 -53 1104 -51
rect 1094 -54 1104 -53
rect 1112 -51 1116 -49
rect 1112 -53 1113 -51
rect 1115 -53 1116 -51
rect 1112 -59 1116 -53
rect 1150 -59 1154 -47
rect 1168 -45 1169 -43
rect 1171 -45 1172 -43
rect 1168 -57 1172 -45
rect 1168 -59 1169 -57
rect 1171 -59 1172 -57
rect 137 -82 143 -75
rect 137 -84 139 -82
rect 141 -84 143 -82
rect 137 -85 143 -84
rect 130 -101 131 -94
rect 130 -119 131 -113
rect 141 -118 145 -116
rect 141 -120 142 -118
rect 144 -120 145 -118
rect 141 -131 145 -120
<< via1 >>
rect 143 -40 145 -38
rect 141 -109 143 -107
<< labels >>
rlabel alu0 58 30 58 30 6 ci
rlabel alu0 54 46 54 46 6 ci
rlabel alu0 96 41 96 41 6 ci
rlabel alu0 105 29 105 29 6 ci
rlabel alu0 131 37 131 37 6 cn
rlabel alu0 120 54 120 54 6 ci
rlabel alu0 140 42 140 42 6 cn
rlabel alu1 77 9 77 9 6 vss
rlabel alu1 77 73 77 73 6 vdd
rlabel alu1 121 45 121 45 6 cp
rlabel alu1 129 49 129 49 6 cp
rlabel alu1 9 41 9 41 1 a7
rlabel alu1 17 45 17 45 1 a7
rlabel alu1 113 37 113 37 1 ain7
rlabel alu1 105 41 105 41 1 ain7
rlabel alu0 22 36 22 36 1 zna7
rlabel alu0 28 36 28 36 1 zna7
rlabel alu0 41 37 41 37 1 n4a7
rlabel alu0 52 21 52 21 1 n4a7
rlabel alu0 51 56 51 56 1 n4a7
rlabel alu0 66 38 66 38 1 n2a7
rlabel alu0 73 46 73 46 1 n2a7
rlabel alu0 78 31 78 31 1 n1a7
rlabel alu0 88 21 88 21 1 n1a7
rlabel alu0 91 62 91 62 1 n1a7
rlabel alu0 206 30 206 30 6 ci
rlabel alu0 202 46 202 46 6 ci
rlabel alu0 244 41 244 41 6 ci
rlabel alu0 253 29 253 29 6 ci
rlabel alu0 279 37 279 37 6 cn
rlabel alu0 268 54 268 54 6 ci
rlabel alu0 288 42 288 42 6 cn
rlabel alu1 225 9 225 9 6 vss
rlabel alu1 225 73 225 73 6 vdd
rlabel alu1 269 45 269 45 6 cp
rlabel alu1 277 49 277 49 6 cp
rlabel alu1 157 41 157 41 1 a6
rlabel alu1 165 45 165 45 1 a6
rlabel alu0 170 36 170 36 1 zna6
rlabel alu0 176 36 176 36 1 zna6
rlabel alu0 189 37 189 37 1 n4a6
rlabel alu0 200 21 200 21 1 n4a6
rlabel alu0 199 56 199 56 1 n4a6
rlabel alu0 214 38 214 38 1 n2a6
rlabel alu0 221 46 221 46 1 n2a6
rlabel alu0 226 31 226 31 1 n1a6
rlabel alu0 236 21 236 21 1 n1a6
rlabel alu0 239 62 239 62 1 n1a6
rlabel alu1 253 41 253 41 1 ain6
rlabel alu1 261 37 261 37 1 ain6
rlabel alu0 354 30 354 30 6 ci
rlabel alu0 350 46 350 46 6 ci
rlabel alu0 392 41 392 41 6 ci
rlabel alu0 401 29 401 29 6 ci
rlabel alu0 427 37 427 37 6 cn
rlabel alu0 416 54 416 54 6 ci
rlabel alu0 436 42 436 42 6 cn
rlabel alu1 373 9 373 9 6 vss
rlabel alu1 373 73 373 73 6 vdd
rlabel alu1 417 45 417 45 6 cp
rlabel alu1 425 49 425 49 6 cp
rlabel alu1 305 41 305 41 1 a5
rlabel alu1 313 45 313 45 1 a5
rlabel alu0 318 36 318 36 1 zna5
rlabel alu0 324 36 324 36 1 zna5
rlabel alu0 337 37 337 37 1 n4a5
rlabel alu0 347 56 347 56 1 n4a5
rlabel alu0 348 21 348 21 1 n4a5
rlabel alu0 362 38 362 38 1 n2a5
rlabel alu0 369 46 369 46 1 n2a5
rlabel alu0 374 31 374 31 1 n1a5
rlabel alu0 387 62 387 62 1 n1a5
rlabel alu0 384 21 384 21 1 n1a5
rlabel alu1 401 41 401 41 1 ain5
rlabel alu1 409 37 409 37 1 ain5
rlabel alu0 502 30 502 30 6 ci
rlabel alu0 498 46 498 46 6 ci
rlabel alu0 540 41 540 41 6 ci
rlabel alu0 549 29 549 29 6 ci
rlabel alu0 575 37 575 37 6 cn
rlabel alu0 564 54 564 54 6 ci
rlabel alu0 584 42 584 42 6 cn
rlabel alu1 521 9 521 9 6 vss
rlabel alu1 521 73 521 73 6 vdd
rlabel alu1 565 45 565 45 6 cp
rlabel alu1 573 49 573 49 6 cp
rlabel alu1 453 41 453 41 1 a4
rlabel alu1 461 45 461 45 1 a4
rlabel alu0 466 36 466 36 1 zna4
rlabel alu0 472 36 472 36 1 zna4
rlabel alu0 485 37 485 37 1 n4a4
rlabel alu0 496 21 496 21 1 n4a4
rlabel alu0 495 56 495 56 1 n4a4
rlabel alu0 510 38 510 38 1 n2a4
rlabel alu0 517 46 517 46 1 n2a4
rlabel alu0 522 31 522 31 1 n1a4
rlabel alu0 532 21 532 21 1 n1a4
rlabel alu0 535 62 535 62 1 n1a4
rlabel alu1 549 41 549 41 1 ain4
rlabel alu1 557 37 557 37 1 ain4
rlabel alu0 650 30 650 30 6 ci
rlabel alu0 646 46 646 46 6 ci
rlabel alu0 688 41 688 41 6 ci
rlabel alu0 697 29 697 29 6 ci
rlabel alu0 723 37 723 37 6 cn
rlabel alu0 712 54 712 54 6 ci
rlabel alu0 732 42 732 42 6 cn
rlabel alu1 669 9 669 9 6 vss
rlabel alu1 669 73 669 73 6 vdd
rlabel alu1 713 45 713 45 6 cp
rlabel alu1 721 49 721 49 6 cp
rlabel alu1 601 41 601 41 1 a3
rlabel alu1 609 45 609 45 1 a3
rlabel alu0 614 36 614 36 1 zna3
rlabel alu0 620 36 620 36 1 zna3
rlabel alu0 633 37 633 37 1 n4a3
rlabel alu0 644 21 644 21 1 n4a3
rlabel alu0 643 56 643 56 1 n4a3
rlabel alu0 658 38 658 38 1 n2a3
rlabel alu0 665 46 665 46 1 n2a3
rlabel alu0 670 31 670 31 1 n1a3
rlabel alu0 680 21 680 21 1 n1a3
rlabel alu0 683 62 683 62 1 n1a3
rlabel alu1 697 41 697 41 1 ain3
rlabel alu1 705 37 705 37 1 ain3
rlabel alu0 798 30 798 30 6 ci
rlabel alu0 794 46 794 46 6 ci
rlabel alu0 836 41 836 41 6 ci
rlabel alu0 845 29 845 29 6 ci
rlabel alu0 871 37 871 37 6 cn
rlabel alu0 860 54 860 54 6 ci
rlabel alu0 880 42 880 42 6 cn
rlabel alu1 817 9 817 9 6 vss
rlabel alu1 817 73 817 73 6 vdd
rlabel alu1 861 45 861 45 6 cp
rlabel alu1 869 49 869 49 6 cp
rlabel alu1 749 41 749 41 1 a2
rlabel alu1 757 45 757 45 1 a2
rlabel alu0 762 36 762 36 1 zna2
rlabel alu0 768 36 768 36 1 zna2
rlabel alu0 781 37 781 37 1 n4a2
rlabel alu0 792 21 792 21 1 n4a2
rlabel alu0 791 56 791 56 1 n4a2
rlabel alu0 806 38 806 38 1 n2a2
rlabel alu0 813 46 813 46 1 n2a2
rlabel alu0 818 31 818 31 1 n1a2
rlabel alu0 828 21 828 21 1 n1a2
rlabel alu0 831 62 831 62 1 n1a2
rlabel alu1 845 41 845 41 1 ain2
rlabel alu1 853 37 853 37 1 ain2
rlabel alu0 946 30 946 30 6 ci
rlabel alu0 942 46 942 46 6 ci
rlabel alu0 984 41 984 41 6 ci
rlabel alu0 993 29 993 29 6 ci
rlabel alu0 1019 37 1019 37 6 cn
rlabel alu0 1008 54 1008 54 6 ci
rlabel alu0 1028 42 1028 42 6 cn
rlabel alu1 965 9 965 9 6 vss
rlabel alu1 965 73 965 73 6 vdd
rlabel alu1 1009 45 1009 45 6 cp
rlabel alu1 1017 49 1017 49 6 cp
rlabel alu1 897 41 897 41 1 a1
rlabel alu1 905 45 905 45 1 a1
rlabel alu0 910 36 910 36 1 zna1
rlabel alu0 916 36 916 36 1 zna1
rlabel alu0 929 37 929 37 1 n4a1
rlabel alu0 940 21 940 21 1 n4a1
rlabel alu0 939 56 939 56 1 n4a1
rlabel alu0 954 38 954 38 1 n2a1
rlabel alu0 961 46 961 46 1 n2a1
rlabel alu0 966 31 966 31 1 n1a1
rlabel alu0 976 21 976 21 1 n1a1
rlabel alu0 979 62 979 62 1 n1a1
rlabel alu1 993 41 993 41 1 ain1
rlabel alu1 1001 37 1001 37 1 ain1
rlabel alu0 1094 30 1094 30 6 ci
rlabel alu0 1090 46 1090 46 6 ci
rlabel alu0 1141 29 1141 29 6 ci
rlabel alu0 1167 37 1167 37 6 cn
rlabel alu0 1156 54 1156 54 6 ci
rlabel alu1 1113 9 1113 9 6 vss
rlabel alu1 1113 73 1113 73 6 vdd
rlabel alu1 1157 45 1157 45 6 cp
rlabel alu1 1165 49 1165 49 6 cp
rlabel alu1 1045 41 1045 41 1 a0
rlabel alu1 1053 45 1053 45 1 a0
rlabel alu0 1058 36 1058 36 1 zna0
rlabel alu0 1064 36 1064 36 1 zna0
rlabel alu0 1077 37 1077 37 1 n4a0
rlabel alu0 1088 21 1088 21 1 n4a0
rlabel alu0 1087 56 1087 56 1 n4a0
rlabel alu0 1102 38 1102 38 1 n2a0
rlabel alu0 1109 46 1109 46 1 n2a0
rlabel alu0 1114 31 1114 31 1 n1a0
rlabel alu0 1124 21 1124 21 1 n1a0
rlabel alu0 1127 62 1127 62 1 n1a0
rlabel alu1 1141 41 1141 41 1 ain0
rlabel alu1 1149 37 1149 37 1 ain0
rlabel alu0 96 -20 96 -20 2 ci
rlabel alu0 100 -36 100 -36 2 ci
rlabel alu0 58 -31 58 -31 2 ci
rlabel alu0 49 -19 49 -19 2 ci
rlabel alu0 23 -27 23 -27 2 cn
rlabel alu0 34 -44 34 -44 2 ci
rlabel alu0 14 -32 14 -32 2 cn
rlabel alu1 77 1 77 1 2 vss
rlabel alu1 77 -63 77 -63 2 vdd
rlabel alu1 33 -35 33 -35 2 cp
rlabel alu1 25 -39 25 -39 2 cp
rlabel alu1 145 -31 145 -31 1 b7
rlabel alu1 137 -35 137 -35 1 b7
rlabel alu0 132 -26 132 -26 1 znb7
rlabel alu0 126 -26 126 -26 1 znb7
rlabel alu0 113 -27 113 -27 1 n4b7
rlabel alu0 102 -11 102 -11 1 n4b7
rlabel alu0 103 -46 103 -46 1 n4b7
rlabel alu0 88 -28 88 -28 1 n2b7
rlabel alu0 81 -36 81 -36 1 n2b7
rlabel alu0 76 -21 76 -21 1 n1b7
rlabel alu0 66 -11 66 -11 1 n1b7
rlabel alu0 63 -52 63 -52 1 n1b7
rlabel alu1 49 -31 49 -31 1 bin7
rlabel alu1 41 -27 41 -27 1 bin7
rlabel alu0 244 -20 244 -20 2 ci
rlabel alu0 248 -36 248 -36 2 ci
rlabel alu0 206 -31 206 -31 2 ci
rlabel alu0 197 -19 197 -19 2 ci
rlabel alu0 171 -27 171 -27 2 cn
rlabel alu0 182 -44 182 -44 2 ci
rlabel alu0 162 -32 162 -32 2 cn
rlabel alu1 225 1 225 1 2 vss
rlabel alu1 225 -63 225 -63 2 vdd
rlabel alu1 181 -35 181 -35 2 cp
rlabel alu1 173 -39 173 -39 2 cp
rlabel alu1 189 -27 189 -27 1 bin6
rlabel alu1 197 -31 197 -31 1 bin6
rlabel alu0 211 -52 211 -52 1 n1b6
rlabel alu0 224 -21 224 -21 1 n1b6
rlabel alu0 214 -11 214 -11 1 n1b6
rlabel alu0 236 -28 236 -28 1 n2b6
rlabel alu0 229 -36 229 -36 1 n2b6
rlabel alu0 250 -11 250 -11 1 n4b6
rlabel alu0 251 -46 251 -46 1 n4b6
rlabel alu0 261 -27 261 -27 1 n4b6
rlabel alu0 274 -26 274 -26 1 znb6
rlabel alu0 280 -26 280 -26 1 znb6
rlabel alu1 293 -31 293 -31 1 b6
rlabel alu1 285 -35 285 -35 1 b6
rlabel alu0 392 -20 392 -20 2 ci
rlabel alu0 396 -36 396 -36 2 ci
rlabel alu0 354 -31 354 -31 2 ci
rlabel alu0 345 -19 345 -19 2 ci
rlabel alu0 319 -27 319 -27 2 cn
rlabel alu0 330 -44 330 -44 2 ci
rlabel alu0 310 -32 310 -32 2 cn
rlabel alu1 373 1 373 1 2 vss
rlabel alu1 373 -63 373 -63 2 vdd
rlabel alu1 329 -35 329 -35 2 cp
rlabel alu1 321 -39 321 -39 2 cp
rlabel alu1 337 -27 337 -27 1 bin5
rlabel alu1 345 -31 345 -31 1 bin5
rlabel alu0 359 -52 359 -52 1 n1b5
rlabel alu0 372 -21 372 -21 1 n1b5
rlabel alu0 362 -11 362 -11 1 n1b5
rlabel alu0 377 -36 377 -36 1 n2b5
rlabel alu0 384 -28 384 -28 1 n2b5
rlabel alu0 399 -46 399 -46 1 n4b5
rlabel alu0 398 -11 398 -11 1 n4b5
rlabel alu0 409 -27 409 -27 1 n4b5
rlabel alu0 422 -26 422 -26 1 znb5
rlabel alu0 428 -26 428 -26 1 znb5
rlabel alu1 433 -35 433 -35 1 b5
rlabel alu1 441 -31 441 -31 1 b5
rlabel alu0 540 -20 540 -20 2 ci
rlabel alu0 544 -36 544 -36 2 ci
rlabel alu0 502 -31 502 -31 2 ci
rlabel alu0 493 -19 493 -19 2 ci
rlabel alu0 467 -27 467 -27 2 cn
rlabel alu0 478 -44 478 -44 2 ci
rlabel alu0 458 -32 458 -32 2 cn
rlabel alu1 521 1 521 1 2 vss
rlabel alu1 521 -63 521 -63 2 vdd
rlabel alu1 477 -35 477 -35 2 cp
rlabel alu1 469 -39 469 -39 2 cp
rlabel alu1 485 -27 485 -27 1 bin4
rlabel alu1 493 -31 493 -31 1 bin4
rlabel alu0 507 -52 507 -52 1 n1b4
rlabel alu0 520 -21 520 -21 1 n1b4
rlabel alu0 510 -11 510 -11 1 n1b4
rlabel alu0 525 -36 525 -36 1 n2b4
rlabel alu0 532 -28 532 -28 1 n2b4
rlabel alu0 547 -46 547 -46 1 n4b4
rlabel alu0 557 -27 557 -27 1 n4b4
rlabel alu0 546 -11 546 -11 1 n4b4
rlabel alu0 570 -26 570 -26 1 znb4
rlabel alu0 576 -26 576 -26 1 znb4
rlabel alu1 581 -35 581 -35 1 b4
rlabel alu1 589 -31 589 -31 1 b4
rlabel alu0 688 -20 688 -20 2 ci
rlabel alu0 692 -36 692 -36 2 ci
rlabel alu0 650 -31 650 -31 2 ci
rlabel alu0 641 -19 641 -19 2 ci
rlabel alu0 615 -27 615 -27 2 cn
rlabel alu0 626 -44 626 -44 2 ci
rlabel alu0 606 -32 606 -32 2 cn
rlabel alu1 669 1 669 1 2 vss
rlabel alu1 669 -63 669 -63 2 vdd
rlabel alu1 625 -35 625 -35 2 cp
rlabel alu1 617 -39 617 -39 2 cp
rlabel alu1 633 -27 633 -27 1 bin3
rlabel alu1 641 -31 641 -31 1 bin3
rlabel alu0 658 -11 658 -11 1 n1b3
rlabel alu0 655 -52 655 -52 1 n1b3
rlabel alu0 668 -21 668 -21 1 n1b3
rlabel alu0 673 -36 673 -36 1 n2b3
rlabel alu0 680 -28 680 -28 1 n2b3
rlabel alu0 695 -46 695 -46 1 n4b3
rlabel alu0 705 -27 705 -27 1 n4b3
rlabel alu0 694 -11 694 -11 1 n4b3
rlabel alu0 718 -26 718 -26 1 znb3
rlabel alu0 724 -26 724 -26 1 znb3
rlabel alu1 729 -35 729 -35 1 b3
rlabel alu1 737 -31 737 -31 1 b3
rlabel alu0 836 -20 836 -20 2 ci
rlabel alu0 840 -36 840 -36 2 ci
rlabel alu0 798 -31 798 -31 2 ci
rlabel alu0 789 -19 789 -19 2 ci
rlabel alu0 763 -27 763 -27 2 cn
rlabel alu0 774 -44 774 -44 2 ci
rlabel alu0 754 -32 754 -32 2 cn
rlabel alu1 817 1 817 1 2 vss
rlabel alu1 817 -63 817 -63 2 vdd
rlabel alu1 773 -35 773 -35 2 cp
rlabel alu1 765 -39 765 -39 2 cp
rlabel alu1 781 -27 781 -27 1 bin2
rlabel alu1 789 -31 789 -31 1 bin2
rlabel alu0 803 -52 803 -52 1 n1b2
rlabel alu0 806 -11 806 -11 1 n1b2
rlabel alu0 816 -21 816 -21 1 n1b2
rlabel alu0 821 -36 821 -36 1 n2b2
rlabel alu0 828 -28 828 -28 1 n2b2
rlabel alu0 843 -46 843 -46 1 n4b2
rlabel alu0 853 -27 853 -27 1 n4b2
rlabel alu0 842 -11 842 -11 1 n4b2
rlabel alu0 866 -26 866 -26 1 znb2
rlabel alu0 872 -26 872 -26 1 znb2
rlabel alu1 877 -35 877 -35 1 b2
rlabel alu1 885 -31 885 -31 1 b2
rlabel alu0 984 -20 984 -20 2 ci
rlabel alu0 988 -36 988 -36 2 ci
rlabel alu0 946 -31 946 -31 2 ci
rlabel alu0 937 -19 937 -19 2 ci
rlabel alu0 911 -27 911 -27 2 cn
rlabel alu0 922 -44 922 -44 2 ci
rlabel alu0 902 -32 902 -32 2 cn
rlabel alu1 965 1 965 1 2 vss
rlabel alu1 965 -63 965 -63 2 vdd
rlabel alu1 921 -35 921 -35 2 cp
rlabel alu1 913 -39 913 -39 2 cp
rlabel alu1 929 -27 929 -27 1 bin1
rlabel alu1 937 -31 937 -31 1 bin1
rlabel alu0 954 -11 954 -11 1 n1b1
rlabel alu0 951 -52 951 -52 1 n1b1
rlabel alu0 964 -21 964 -21 1 n1b1
rlabel alu0 969 -36 969 -36 1 n2b1
rlabel alu0 976 -28 976 -28 1 n2b1
rlabel alu0 991 -46 991 -46 1 n4b1
rlabel alu0 990 -11 990 -11 1 n4b1
rlabel alu0 1001 -27 1001 -27 1 n4b1
rlabel alu0 1014 -26 1014 -26 1 znb1
rlabel alu0 1020 -26 1020 -26 1 znb1
rlabel alu1 1025 -35 1025 -35 1 b1
rlabel alu1 1033 -31 1033 -31 1 b1
rlabel alu0 1176 42 1176 42 6 cn
rlabel alu0 1132 41 1132 41 6 ci
rlabel alu0 1132 -20 1132 -20 2 ci
rlabel alu0 1136 -36 1136 -36 2 ci
rlabel alu0 1094 -31 1094 -31 2 ci
rlabel alu0 1085 -19 1085 -19 2 ci
rlabel alu0 1059 -27 1059 -27 2 cn
rlabel alu0 1070 -44 1070 -44 2 ci
rlabel alu0 1050 -32 1050 -32 2 cn
rlabel alu1 1113 1 1113 1 2 vss
rlabel alu1 1113 -63 1113 -63 2 vdd
rlabel alu1 1069 -35 1069 -35 2 cp
rlabel alu1 1061 -39 1061 -39 2 cp
rlabel alu1 1077 -27 1077 -27 1 bin0
rlabel alu1 1085 -31 1085 -31 1 bin0
rlabel alu0 1099 -52 1099 -52 1 n1b0
rlabel alu0 1112 -21 1112 -21 1 n1b0
rlabel alu0 1102 -11 1102 -11 1 n1b0
rlabel alu0 1117 -36 1117 -36 1 n2b0
rlabel alu0 1124 -28 1124 -28 1 n2b0
rlabel alu0 1139 -46 1139 -46 1 n4b0
rlabel alu0 1149 -27 1149 -27 1 n4b0
rlabel alu0 1138 -11 1138 -11 1 n4b0
rlabel alu0 1162 -26 1162 -26 1 znb0
rlabel alu0 1168 -26 1168 -26 1 znb0
rlabel alu1 1173 -35 1173 -35 1 b0
rlabel alu1 1181 -31 1181 -31 1 b0
rlabel alu1 136 -135 136 -135 6 vss
rlabel alu1 136 -71 136 -71 6 vdd
rlabel alu1 128 -107 128 -107 1 binv7
rlabel alu1 136 -91 136 -91 1 binv7
rlabel alu1 136 -111 136 -111 1 b7
rlabel alu1 144 -107 144 -107 1 b7
<< end >>
