magic
tech scmos
timestamp 1199973029
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -5 40 69 97
<< pwell >>
rect -5 -9 69 40
<< poly >>
rect 2 81 11 83
rect 2 79 7 81
rect 9 79 11 81
rect 2 77 11 79
rect 9 74 11 77
rect 21 77 30 83
rect 34 81 43 83
rect 34 79 39 81
rect 41 79 43 81
rect 34 77 43 79
rect 21 74 23 77
rect 41 74 43 77
rect 53 81 62 83
rect 53 79 55 81
rect 57 79 62 81
rect 53 77 62 79
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 37 14 43
rect 18 41 30 43
rect 18 39 23 41
rect 25 39 30 41
rect 18 37 30 39
rect 34 41 46 43
rect 34 39 36 41
rect 38 39 46 41
rect 34 37 46 39
rect 50 37 62 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndif >>
rect 2 14 9 34
rect 11 25 21 34
rect 11 23 15 25
rect 17 23 21 25
rect 11 18 21 23
rect 11 16 15 18
rect 17 16 21 18
rect 11 14 21 16
rect 23 28 30 34
rect 23 26 26 28
rect 28 26 30 28
rect 23 21 30 26
rect 23 19 26 21
rect 28 19 30 21
rect 23 14 30 19
rect 34 18 41 34
rect 34 16 36 18
rect 38 16 41 18
rect 34 14 41 16
rect 43 29 53 34
rect 43 27 47 29
rect 49 27 53 29
rect 43 21 53 27
rect 43 19 47 21
rect 49 19 53 21
rect 43 14 53 19
rect 55 25 62 34
rect 55 23 58 25
rect 60 23 62 25
rect 55 18 62 23
rect 55 16 58 18
rect 60 16 62 18
rect 55 14 62 16
rect 13 2 19 14
rect 45 2 51 14
<< pdif >>
rect 13 74 19 86
rect 45 74 51 86
rect 2 46 9 74
rect 11 72 21 74
rect 11 70 15 72
rect 17 70 21 72
rect 11 65 21 70
rect 11 63 15 65
rect 17 63 21 65
rect 11 46 21 63
rect 23 61 30 74
rect 23 59 26 61
rect 28 59 30 61
rect 23 54 30 59
rect 23 52 26 54
rect 28 52 30 54
rect 23 46 30 52
rect 34 72 41 74
rect 34 70 36 72
rect 38 70 41 72
rect 34 65 41 70
rect 34 63 36 65
rect 38 63 41 65
rect 34 46 41 63
rect 43 61 53 74
rect 43 59 47 61
rect 49 59 53 61
rect 43 53 53 59
rect 43 51 47 53
rect 49 51 53 53
rect 43 46 53 51
rect 55 71 62 74
rect 55 69 58 71
rect 60 69 62 71
rect 55 64 62 69
rect 55 62 58 64
rect 60 62 62 64
rect 55 46 62 62
<< alu1 >>
rect -2 89 66 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 66 89
rect -2 86 66 87
rect 6 81 10 86
rect 6 79 7 81
rect 9 79 10 81
rect 6 77 10 79
rect 14 81 18 86
rect 14 79 15 81
rect 17 79 18 81
rect 14 73 18 79
rect 14 72 61 73
rect 14 70 15 72
rect 17 70 36 72
rect 38 71 61 72
rect 38 70 58 71
rect 14 69 58 70
rect 60 69 61 71
rect 14 65 18 69
rect 14 63 15 65
rect 17 63 18 65
rect 35 65 39 69
rect 35 63 36 65
rect 38 63 39 65
rect 57 64 61 69
rect 14 61 18 63
rect 22 61 29 63
rect 35 61 39 63
rect 46 61 50 63
rect 22 59 26 61
rect 28 59 29 61
rect 22 57 29 59
rect 14 38 18 55
rect 25 54 29 57
rect 46 59 47 61
rect 49 59 50 61
rect 57 62 58 64
rect 60 62 61 64
rect 57 60 61 62
rect 46 54 50 59
rect 25 52 26 54
rect 28 53 50 54
rect 28 52 47 53
rect 25 51 47 52
rect 49 51 50 53
rect 25 50 50 51
rect 22 41 26 43
rect 22 39 23 41
rect 25 39 26 41
rect 22 38 26 39
rect 35 41 39 43
rect 35 39 36 41
rect 38 39 39 41
rect 35 38 39 39
rect 14 34 39 38
rect 14 33 18 34
rect 46 30 50 50
rect 25 29 50 30
rect 25 28 47 29
rect 14 25 18 27
rect 14 23 15 25
rect 17 23 18 25
rect 25 26 26 28
rect 28 27 47 28
rect 49 27 50 29
rect 28 26 50 27
rect 25 23 29 26
rect 14 18 18 23
rect 14 16 15 18
rect 17 16 18 18
rect 22 21 29 23
rect 22 19 26 21
rect 28 19 29 21
rect 46 21 50 26
rect 22 17 29 19
rect 35 18 39 20
rect 14 9 18 16
rect 14 7 15 9
rect 17 7 18 9
rect 14 2 18 7
rect 35 16 36 18
rect 38 16 39 18
rect 46 19 47 21
rect 49 19 50 21
rect 46 17 50 19
rect 57 25 61 27
rect 57 23 58 25
rect 60 23 61 25
rect 57 18 61 23
rect 35 9 39 16
rect 35 7 36 9
rect 38 7 39 9
rect 35 2 39 7
rect 57 16 58 18
rect 60 16 61 18
rect 57 9 61 16
rect 57 7 58 9
rect 60 7 61 9
rect 57 2 61 7
rect -2 1 66 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< alu2 >>
rect -2 89 66 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 66 89
rect -2 81 66 87
rect -2 79 15 81
rect 17 79 66 81
rect -2 76 66 79
rect -2 9 66 12
rect -2 7 15 9
rect 17 7 36 9
rect 38 7 58 9
rect 60 7 66 9
rect -2 1 66 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 64 3
rect 57 -1 59 1
rect 61 -1 64 1
rect 57 -3 64 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 64 91
rect 57 87 59 89
rect 61 87 64 89
rect 57 85 64 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< polyct0 >>
rect 39 79 41 81
rect 55 79 57 81
<< polyct1 >>
rect 7 79 9 81
rect 23 39 25 41
rect 36 39 38 41
<< ndifct1 >>
rect 15 23 17 25
rect 15 16 17 18
rect 26 26 28 28
rect 26 19 28 21
rect 36 16 38 18
rect 47 27 49 29
rect 47 19 49 21
rect 58 23 60 25
rect 58 16 60 18
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
<< pdifct1 >>
rect 15 70 17 72
rect 15 63 17 65
rect 26 59 28 61
rect 26 52 28 54
rect 36 70 38 72
rect 36 63 38 65
rect 47 59 49 61
rect 47 51 49 53
rect 58 69 60 71
rect 58 62 60 64
<< alu0 >>
rect 37 81 59 82
rect 37 79 39 81
rect 41 79 55 81
rect 57 79 59 81
rect 37 78 59 79
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 15 79 17 81
rect 15 7 17 9
rect 36 7 38 9
rect 58 7 60 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
<< labels >>
rlabel alu1 24 20 24 20 6 z
rlabel alu1 24 36 24 36 6 a
rlabel alu1 16 44 16 44 6 a
rlabel alu1 24 60 24 60 6 z
rlabel alu1 32 28 32 28 6 z
rlabel alu1 32 36 32 36 6 a
rlabel alu1 40 28 40 28 6 z
rlabel alu1 32 52 32 52 6 z
rlabel alu1 40 52 40 52 6 z
rlabel alu1 48 40 48 40 6 z
rlabel alu2 32 6 32 6 6 vss
rlabel alu2 32 82 32 82 6 vdd
<< end >>
