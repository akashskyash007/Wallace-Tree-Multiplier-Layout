magic
tech scmos
timestamp 1199202035
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 9 34 11 38
rect 19 34 21 38
rect 29 35 31 38
rect 9 32 22 34
rect 9 30 18 32
rect 20 30 22 32
rect 9 28 22 30
rect 26 33 32 35
rect 26 31 28 33
rect 30 31 32 33
rect 26 29 32 31
rect 9 25 11 28
rect 19 25 21 28
rect 29 25 31 29
rect 9 6 11 11
rect 19 6 21 11
rect 29 6 31 11
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 15 9 21
rect 2 13 4 15
rect 6 13 9 15
rect 2 11 9 13
rect 11 17 19 25
rect 11 15 14 17
rect 16 15 19 17
rect 11 11 19 15
rect 21 15 29 25
rect 21 13 24 15
rect 26 13 29 15
rect 21 11 29 13
rect 31 23 38 25
rect 31 21 34 23
rect 36 21 38 23
rect 31 16 38 21
rect 31 14 34 16
rect 36 14 38 16
rect 31 11 38 14
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 51 36 66
rect 31 49 38 51
rect 31 47 34 49
rect 36 47 38 49
rect 31 42 38 47
rect 31 40 34 42
rect 36 40 38 42
rect 31 38 38 40
<< alu1 >>
rect -2 64 42 72
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 50 17 55
rect 2 48 14 50
rect 16 48 17 50
rect 2 46 17 48
rect 2 33 6 46
rect 17 38 30 42
rect 26 35 30 38
rect 2 29 14 33
rect 10 19 14 29
rect 26 33 31 35
rect 26 31 28 33
rect 30 31 31 33
rect 26 29 31 31
rect 10 17 17 19
rect 10 15 14 17
rect 16 15 17 17
rect 10 13 17 15
rect -2 0 42 8
<< nmos >>
rect 9 11 11 25
rect 19 11 21 25
rect 29 11 31 25
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
<< polyct0 >>
rect 18 30 20 32
<< polyct1 >>
rect 28 31 30 33
<< ndifct0 >>
rect 4 21 6 23
rect 4 13 6 15
rect 24 13 26 15
rect 34 21 36 23
rect 34 14 36 16
<< ndifct1 >>
rect 14 15 16 17
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 24 62 26 64
rect 24 55 26 57
rect 34 47 36 49
rect 34 40 36 42
<< pdifct1 >>
rect 14 55 16 57
rect 14 48 16 50
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 22 57 28 62
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 33 49 38 51
rect 33 47 34 49
rect 36 47 38 49
rect 33 42 38 47
rect 33 40 34 42
rect 36 40 38 42
rect 33 38 38 40
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 15 7 21
rect 3 13 4 15
rect 6 13 7 15
rect 17 32 21 34
rect 17 30 18 32
rect 20 30 21 32
rect 17 26 21 30
rect 34 26 38 38
rect 17 23 38 26
rect 17 22 34 23
rect 32 21 34 22
rect 36 21 38 23
rect 23 15 27 17
rect 23 13 24 15
rect 26 13 27 15
rect 32 16 38 21
rect 32 14 34 16
rect 36 14 38 16
rect 32 13 38 14
rect 3 8 7 13
rect 23 8 27 13
<< labels >>
rlabel alu0 19 28 19 28 6 an
rlabel alu0 36 32 36 32 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 28 32 28 32 6 a
rlabel alu1 20 40 20 40 6 a
rlabel alu1 20 68 20 68 6 vdd
<< end >>
