magic
tech scmos
timestamp 1199203508
<< ab >>
rect 0 0 128 72
<< nwell >>
rect -5 32 133 77
<< pwell >>
rect -5 -5 133 32
<< poly >>
rect 37 65 39 70
rect 47 65 49 70
rect 54 65 56 70
rect 9 57 11 61
rect 19 57 21 61
rect 85 61 87 66
rect 97 61 99 66
rect 107 61 109 66
rect 117 61 119 66
rect 9 35 11 38
rect 19 35 21 38
rect 37 35 39 46
rect 47 35 49 46
rect 54 43 56 46
rect 72 44 78 46
rect 53 41 59 43
rect 53 39 55 41
rect 57 39 59 41
rect 72 42 74 44
rect 76 42 78 44
rect 85 42 87 45
rect 72 40 87 42
rect 53 37 59 39
rect 9 33 15 35
rect 19 33 39 35
rect 43 33 49 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 25 31 27 33
rect 29 31 35 33
rect 25 29 35 31
rect 43 31 45 33
rect 47 31 49 33
rect 43 29 49 31
rect 13 21 15 29
rect 33 26 35 29
rect 45 26 47 29
rect 57 26 59 37
rect 97 36 99 45
rect 63 34 99 36
rect 107 35 109 45
rect 117 36 119 45
rect 63 32 65 34
rect 67 32 69 34
rect 63 30 69 32
rect 73 28 79 30
rect 73 26 75 28
rect 77 26 79 28
rect 73 24 79 26
rect 77 21 79 24
rect 33 12 35 17
rect 45 12 47 17
rect 57 12 59 17
rect 89 19 91 34
rect 103 33 109 35
rect 103 31 105 33
rect 107 31 109 33
rect 103 29 109 31
rect 113 34 119 36
rect 113 32 115 34
rect 117 32 119 34
rect 113 30 119 32
rect 107 25 109 29
rect 99 19 101 24
rect 107 22 111 25
rect 109 19 111 22
rect 116 19 118 30
rect 13 7 15 12
rect 77 4 79 14
rect 89 8 91 12
rect 99 4 101 12
rect 109 7 111 12
rect 116 7 118 12
rect 77 2 101 4
<< ndif >>
rect 17 21 33 26
rect 8 18 13 21
rect 6 16 13 18
rect 6 14 8 16
rect 10 14 13 16
rect 6 12 13 14
rect 15 17 33 21
rect 35 24 45 26
rect 35 22 38 24
rect 40 22 45 24
rect 35 17 45 22
rect 47 24 57 26
rect 47 22 52 24
rect 54 22 57 24
rect 47 17 57 22
rect 59 23 64 26
rect 59 21 66 23
rect 59 19 62 21
rect 64 19 66 21
rect 59 17 66 19
rect 70 19 77 21
rect 70 17 72 19
rect 74 17 77 19
rect 15 12 31 17
rect 70 14 77 17
rect 79 19 87 21
rect 79 14 89 19
rect 17 7 31 12
rect 17 5 19 7
rect 21 5 27 7
rect 29 5 31 7
rect 17 3 31 5
rect 81 12 89 14
rect 91 17 99 19
rect 91 15 94 17
rect 96 15 99 17
rect 91 12 99 15
rect 101 17 109 19
rect 101 15 104 17
rect 106 15 109 17
rect 101 12 109 15
rect 111 12 116 19
rect 118 12 126 19
rect 81 11 87 12
rect 81 9 83 11
rect 85 9 87 11
rect 81 7 87 9
rect 120 7 126 12
rect 120 5 122 7
rect 124 5 126 7
rect 120 3 126 5
<< pdif >>
rect 13 67 19 69
rect 13 65 15 67
rect 17 65 19 67
rect 89 67 95 69
rect 13 63 19 65
rect 13 57 17 63
rect 32 60 37 65
rect 30 58 37 60
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 48 9 53
rect 2 46 4 48
rect 6 46 9 48
rect 2 44 9 46
rect 4 38 9 44
rect 11 38 19 57
rect 21 50 26 57
rect 30 56 32 58
rect 34 56 37 58
rect 30 54 37 56
rect 21 48 28 50
rect 21 46 24 48
rect 26 46 28 48
rect 32 46 37 54
rect 39 57 47 65
rect 39 55 42 57
rect 44 55 47 57
rect 39 46 47 55
rect 49 46 54 65
rect 56 63 64 65
rect 56 61 59 63
rect 61 61 64 63
rect 56 56 64 61
rect 56 54 59 56
rect 61 54 64 56
rect 56 46 64 54
rect 89 65 91 67
rect 93 65 95 67
rect 89 61 95 65
rect 78 58 85 61
rect 78 56 80 58
rect 82 56 85 58
rect 78 54 85 56
rect 21 44 28 46
rect 21 38 26 44
rect 80 45 85 54
rect 87 45 97 61
rect 99 49 107 61
rect 99 47 102 49
rect 104 47 107 49
rect 99 45 107 47
rect 109 50 117 61
rect 109 48 112 50
rect 114 48 117 50
rect 109 45 117 48
rect 119 58 126 61
rect 119 56 122 58
rect 124 56 126 58
rect 119 54 126 56
rect 119 45 124 54
<< alu1 >>
rect -2 67 130 72
rect -2 65 5 67
rect 7 65 15 67
rect 17 65 70 67
rect 72 65 91 67
rect 93 65 130 67
rect -2 64 130 65
rect 74 46 87 50
rect 10 38 23 42
rect 10 33 14 38
rect 10 31 11 33
rect 13 31 14 33
rect 10 21 14 31
rect 25 33 31 34
rect 25 31 27 33
rect 29 31 31 33
rect 25 27 31 31
rect 18 21 31 27
rect 74 44 78 46
rect 76 42 78 44
rect 74 28 78 42
rect 110 50 126 51
rect 110 48 112 50
rect 114 48 126 50
rect 110 46 126 48
rect 74 26 75 28
rect 77 26 78 28
rect 74 24 78 26
rect 122 18 126 46
rect 102 17 126 18
rect 102 15 104 17
rect 106 15 126 17
rect 102 14 126 15
rect -2 7 130 8
rect -2 5 19 7
rect 21 5 27 7
rect 29 5 53 7
rect 55 5 61 7
rect 63 5 122 7
rect 124 5 130 7
rect -2 0 130 5
<< ptie >>
rect 51 7 65 9
rect 51 5 53 7
rect 55 5 61 7
rect 63 5 65 7
rect 51 3 65 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
rect 68 67 74 69
rect 68 65 70 67
rect 72 65 74 67
rect 68 49 74 65
<< nmos >>
rect 13 12 15 21
rect 33 17 35 26
rect 45 17 47 26
rect 57 17 59 26
rect 77 14 79 21
rect 89 12 91 19
rect 99 12 101 19
rect 109 12 111 19
rect 116 12 118 19
<< pmos >>
rect 9 38 11 57
rect 19 38 21 57
rect 37 46 39 65
rect 47 46 49 65
rect 54 46 56 65
rect 85 45 87 61
rect 97 45 99 61
rect 107 45 109 61
rect 117 45 119 61
<< polyct0 >>
rect 55 39 57 41
rect 45 31 47 33
rect 65 32 67 34
rect 105 31 107 33
rect 115 32 117 34
<< polyct1 >>
rect 74 42 76 44
rect 11 31 13 33
rect 27 31 29 33
rect 75 26 77 28
<< ndifct0 >>
rect 8 14 10 16
rect 38 22 40 24
rect 52 22 54 24
rect 62 19 64 21
rect 72 17 74 19
rect 94 15 96 17
rect 83 9 85 11
<< ndifct1 >>
rect 19 5 21 7
rect 27 5 29 7
rect 104 15 106 17
rect 122 5 124 7
<< ntiect1 >>
rect 5 65 7 67
rect 70 65 72 67
<< ptiect1 >>
rect 53 5 55 7
rect 61 5 63 7
<< pdifct0 >>
rect 4 53 6 55
rect 4 46 6 48
rect 32 56 34 58
rect 24 46 26 48
rect 42 55 44 57
rect 59 61 61 63
rect 59 54 61 56
rect 80 56 82 58
rect 102 47 104 49
rect 122 56 124 58
<< pdifct1 >>
rect 15 65 17 67
rect 91 65 93 67
rect 112 48 114 50
<< alu0 >>
rect 57 63 63 64
rect 57 61 59 63
rect 61 61 63 63
rect 2 58 36 59
rect 2 56 32 58
rect 34 56 36 58
rect 2 55 36 56
rect 40 57 51 58
rect 40 55 42 57
rect 44 55 51 57
rect 2 53 4 55
rect 6 53 7 55
rect 40 54 51 55
rect 2 48 7 53
rect 47 50 51 54
rect 57 56 63 61
rect 57 54 59 56
rect 61 54 63 56
rect 78 58 126 59
rect 78 56 80 58
rect 82 56 122 58
rect 124 56 126 58
rect 78 55 126 56
rect 57 53 63 54
rect 2 46 4 48
rect 6 46 7 48
rect 2 44 7 46
rect 22 48 41 49
rect 22 46 24 48
rect 26 46 41 48
rect 47 46 68 50
rect 22 45 41 46
rect 2 17 6 44
rect 37 42 41 45
rect 37 41 59 42
rect 37 39 55 41
rect 57 39 59 41
rect 37 38 59 39
rect 37 24 41 38
rect 37 22 38 24
rect 40 22 41 24
rect 37 20 41 22
rect 44 33 48 35
rect 44 31 45 33
rect 47 31 48 33
rect 64 34 68 46
rect 73 40 74 46
rect 64 32 65 34
rect 67 32 68 34
rect 44 17 48 31
rect 51 28 68 32
rect 92 34 96 55
rect 101 49 105 51
rect 101 47 102 49
rect 104 47 105 49
rect 101 42 105 47
rect 101 38 118 42
rect 114 34 118 38
rect 51 24 55 28
rect 84 33 109 34
rect 84 31 105 33
rect 107 31 109 33
rect 84 30 109 31
rect 114 32 115 34
rect 117 32 118 34
rect 51 22 52 24
rect 54 22 55 24
rect 51 20 55 22
rect 61 21 65 23
rect 61 19 62 21
rect 64 19 65 21
rect 84 20 88 30
rect 114 26 118 32
rect 61 17 65 19
rect 2 16 65 17
rect 70 19 88 20
rect 70 17 72 19
rect 74 17 88 19
rect 70 16 88 17
rect 93 22 118 26
rect 93 17 97 22
rect 2 14 8 16
rect 10 14 65 16
rect 2 13 65 14
rect 93 15 94 17
rect 96 15 97 17
rect 93 13 97 15
rect 81 11 87 12
rect 81 9 83 11
rect 85 9 87 11
rect 81 8 87 9
<< labels >>
rlabel alu0 4 51 4 51 6 an
rlabel alu0 53 26 53 26 6 iz
rlabel alu0 46 24 46 24 6 an
rlabel alu0 48 40 48 40 6 bn
rlabel alu0 39 34 39 34 6 bn
rlabel alu0 31 47 31 47 6 bn
rlabel alu0 45 56 45 56 6 iz
rlabel alu0 19 57 19 57 6 an
rlabel alu0 33 15 33 15 6 an
rlabel alu0 79 18 79 18 6 cn
rlabel alu0 63 18 63 18 6 an
rlabel alu0 66 39 66 39 6 iz
rlabel alu0 95 19 95 19 6 zn
rlabel alu0 96 32 96 32 6 cn
rlabel alu0 103 44 103 44 6 zn
rlabel alu0 116 32 116 32 6 zn
rlabel alu0 102 57 102 57 6 cn
rlabel alu1 28 28 28 28 6 b
rlabel alu1 20 24 20 24 6 b
rlabel alu1 12 28 12 28 6 a
rlabel alu1 20 40 20 40 6 a
rlabel alu1 64 4 64 4 6 vss
rlabel alu1 76 36 76 36 6 c
rlabel alu1 84 48 84 48 6 c
rlabel alu1 64 68 64 68 6 vdd
rlabel alu1 116 16 116 16 6 z
rlabel alu1 108 16 108 16 6 z
rlabel alu1 124 36 124 36 6 z
rlabel alu1 116 48 116 48 6 z
<< end >>
