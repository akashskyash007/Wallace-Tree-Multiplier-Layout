magic
tech scmos
timestamp 1199201757
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 20 65 22 70
rect 30 65 32 70
rect 42 65 44 70
rect 52 65 54 70
rect 9 61 11 65
rect 9 39 11 43
rect 20 39 22 52
rect 30 49 32 52
rect 30 47 37 49
rect 30 45 33 47
rect 35 45 37 47
rect 30 43 37 45
rect 42 47 44 52
rect 42 45 48 47
rect 42 43 44 45
rect 46 43 48 45
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 20 37 26 39
rect 20 35 22 37
rect 24 35 26 37
rect 20 33 26 35
rect 9 28 11 33
rect 24 28 26 33
rect 31 28 33 43
rect 42 41 48 43
rect 42 39 44 41
rect 38 37 44 39
rect 52 39 54 52
rect 52 37 58 39
rect 38 28 40 37
rect 52 35 54 37
rect 56 35 58 37
rect 52 33 58 35
rect 45 31 58 33
rect 45 28 47 31
rect 9 15 11 19
rect 24 7 26 12
rect 31 7 33 12
rect 38 7 40 12
rect 45 7 47 12
<< ndif >>
rect 4 25 9 28
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 19 24 28
rect 13 12 24 19
rect 26 12 31 28
rect 33 12 38 28
rect 40 12 45 28
rect 47 22 52 28
rect 47 20 54 22
rect 47 18 50 20
rect 52 18 54 20
rect 47 16 54 18
rect 47 12 52 16
rect 13 11 22 12
rect 13 9 16 11
rect 18 9 22 11
rect 13 7 22 9
<< pdif >>
rect 34 71 40 73
rect 34 69 36 71
rect 38 69 40 71
rect 34 65 40 69
rect 13 62 20 65
rect 13 61 15 62
rect 4 56 9 61
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 60 15 61
rect 17 60 20 62
rect 11 52 20 60
rect 22 62 30 65
rect 22 60 25 62
rect 27 60 30 62
rect 22 52 30 60
rect 32 52 42 65
rect 44 62 52 65
rect 44 60 47 62
rect 49 60 52 62
rect 44 52 52 60
rect 54 63 61 65
rect 54 61 57 63
rect 59 61 61 63
rect 54 56 61 61
rect 54 54 57 56
rect 59 54 61 56
rect 54 52 61 54
rect 11 43 18 52
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 36 71
rect 38 69 66 71
rect -2 68 66 69
rect 2 54 7 63
rect 2 52 4 54
rect 6 52 7 54
rect 2 47 7 52
rect 2 45 4 47
rect 6 45 7 47
rect 2 43 7 45
rect 2 23 6 43
rect 34 47 38 55
rect 25 45 33 46
rect 35 45 38 47
rect 25 42 38 45
rect 42 46 46 55
rect 42 45 55 46
rect 42 43 44 45
rect 46 43 55 45
rect 42 42 55 43
rect 20 37 31 38
rect 20 35 22 37
rect 24 35 31 37
rect 20 34 31 35
rect 41 37 62 38
rect 41 35 54 37
rect 56 35 62 37
rect 41 34 62 35
rect 27 30 31 34
rect 27 26 47 30
rect 2 21 4 23
rect 6 21 15 22
rect 2 17 15 21
rect 58 17 62 34
rect -2 11 66 12
rect -2 9 16 11
rect 18 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 19 11 28
rect 24 12 26 28
rect 31 12 33 28
rect 38 12 40 28
rect 45 12 47 28
<< pmos >>
rect 9 43 11 61
rect 20 52 22 65
rect 30 52 32 65
rect 42 52 44 65
rect 52 52 54 65
<< polyct0 >>
rect 33 46 34 47
rect 11 35 13 37
<< polyct1 >>
rect 34 46 35 47
rect 33 45 35 46
rect 44 43 46 45
rect 22 35 24 37
rect 54 35 56 37
<< ndifct0 >>
rect 50 18 52 20
<< ndifct1 >>
rect 4 21 6 23
rect 16 9 18 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 15 60 17 62
rect 25 60 27 62
rect 47 60 49 62
rect 57 61 59 63
rect 57 54 59 56
<< pdifct1 >>
rect 36 69 38 71
rect 4 52 6 54
rect 4 45 6 47
<< alu0 >>
rect 14 62 18 68
rect 56 63 60 68
rect 14 60 15 62
rect 17 60 18 62
rect 14 58 18 60
rect 22 62 51 63
rect 22 60 25 62
rect 27 60 47 62
rect 49 60 51 62
rect 22 59 51 60
rect 56 61 57 63
rect 59 61 60 63
rect 22 54 26 59
rect 56 56 60 61
rect 12 50 26 54
rect 12 39 16 50
rect 32 47 34 48
rect 32 46 33 47
rect 56 54 57 56
rect 59 54 60 56
rect 56 52 60 54
rect 10 37 16 39
rect 10 35 11 37
rect 13 35 16 37
rect 10 33 16 35
rect 12 30 16 33
rect 12 26 23 30
rect 6 22 7 25
rect 19 21 23 26
rect 19 20 54 21
rect 19 18 50 20
rect 52 18 54 20
rect 19 17 54 18
<< labels >>
rlabel alu0 14 40 14 40 6 zn
rlabel alu0 36 19 36 19 6 zn
rlabel alu0 36 61 36 61 6 zn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 36 28 36 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 36 44 36 6 d
rlabel alu1 36 52 36 52 6 b
rlabel alu1 44 52 44 52 6 c
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 36 52 36 6 d
rlabel alu1 60 24 60 24 6 d
rlabel alu1 52 44 52 44 6 c
<< end >>
