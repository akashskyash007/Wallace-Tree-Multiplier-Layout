magic
tech scmos
timestamp 1199973067
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -5 40 69 97
<< pwell >>
rect -5 -9 69 40
<< poly >>
rect 2 81 11 83
rect 2 79 7 81
rect 9 79 11 81
rect 2 77 11 79
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 37 14 43
rect 18 41 30 43
rect 18 39 20 41
rect 22 39 30 41
rect 18 37 30 39
rect 34 41 46 43
rect 34 39 39 41
rect 41 39 46 41
rect 34 37 46 39
rect 50 41 62 43
rect 50 39 55 41
rect 57 39 62 41
rect 50 37 62 39
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndif >>
rect 2 14 9 34
rect 11 25 21 34
rect 11 23 15 25
rect 17 23 21 25
rect 11 18 21 23
rect 11 16 15 18
rect 17 16 21 18
rect 11 14 21 16
rect 23 28 30 34
rect 23 26 26 28
rect 28 26 30 28
rect 23 21 30 26
rect 23 19 26 21
rect 28 19 30 21
rect 23 14 30 19
rect 34 20 41 34
rect 34 18 36 20
rect 38 18 41 20
rect 34 14 41 18
rect 43 14 53 34
rect 55 27 62 34
rect 55 25 58 27
rect 60 25 62 27
rect 55 20 62 25
rect 55 18 58 20
rect 60 18 62 20
rect 55 14 62 18
rect 13 2 19 14
rect 45 2 51 14
<< pdif >>
rect 13 74 19 86
rect 45 74 51 86
rect 2 46 9 74
rect 11 72 21 74
rect 11 70 14 72
rect 16 70 21 72
rect 11 65 21 70
rect 11 63 14 65
rect 16 63 21 65
rect 11 46 21 63
rect 23 61 30 74
rect 23 59 26 61
rect 28 59 30 61
rect 23 54 30 59
rect 23 52 26 54
rect 28 52 30 54
rect 23 46 30 52
rect 34 72 41 74
rect 34 70 36 72
rect 38 70 41 72
rect 34 46 41 70
rect 43 58 53 74
rect 43 56 47 58
rect 49 56 53 58
rect 43 50 53 56
rect 43 48 47 50
rect 49 48 53 50
rect 43 46 53 48
rect 55 72 62 74
rect 55 70 58 72
rect 60 70 62 72
rect 55 65 62 70
rect 55 63 58 65
rect 60 63 62 65
rect 55 46 62 63
<< alu1 >>
rect -2 89 66 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 66 89
rect -2 86 66 87
rect 13 81 17 86
rect 13 79 14 81
rect 16 79 17 81
rect 13 72 17 79
rect 13 70 14 72
rect 16 70 17 72
rect 13 65 17 70
rect 35 81 39 86
rect 35 79 36 81
rect 38 79 39 81
rect 35 72 39 79
rect 35 70 36 72
rect 38 70 39 72
rect 35 68 39 70
rect 57 81 61 86
rect 57 79 58 81
rect 60 79 61 81
rect 57 72 61 79
rect 57 70 58 72
rect 60 70 61 72
rect 13 63 14 65
rect 16 63 17 65
rect 57 65 61 70
rect 57 63 58 65
rect 60 63 61 65
rect 13 61 17 63
rect 21 61 50 63
rect 57 61 61 63
rect 21 59 26 61
rect 28 59 50 61
rect 21 58 50 59
rect 25 54 29 58
rect 13 42 19 54
rect 25 52 26 54
rect 28 52 29 54
rect 25 50 29 52
rect 46 56 47 58
rect 49 56 50 58
rect 46 50 50 56
rect 46 48 47 50
rect 49 48 50 50
rect 13 41 24 42
rect 13 39 20 41
rect 22 39 24 41
rect 13 38 24 39
rect 38 41 42 47
rect 38 39 39 41
rect 41 39 42 41
rect 13 34 19 38
rect 14 25 18 27
rect 14 23 15 25
rect 17 23 18 25
rect 14 18 18 23
rect 14 16 15 18
rect 17 16 18 18
rect 38 25 42 39
rect 46 29 50 48
rect 54 41 58 55
rect 54 39 55 41
rect 57 39 58 41
rect 54 33 58 39
rect 46 27 61 29
rect 46 25 58 27
rect 60 25 61 27
rect 54 20 61 25
rect 54 18 58 20
rect 60 18 61 20
rect 54 16 61 18
rect 14 9 18 16
rect 14 7 15 9
rect 17 7 18 9
rect 14 2 18 7
rect -2 1 66 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< alu2 >>
rect -2 89 66 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 66 89
rect -2 81 66 87
rect -2 79 14 81
rect 16 79 36 81
rect 38 79 58 81
rect 60 79 66 81
rect -2 76 66 79
rect -2 9 66 12
rect -2 7 15 9
rect 17 7 66 9
rect -2 1 66 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 64 3
rect 57 -1 59 1
rect 61 -1 64 1
rect 57 -3 64 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 64 91
rect 57 87 59 89
rect 61 87 64 89
rect 57 85 64 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< polyct0 >>
rect 7 79 9 81
<< polyct1 >>
rect 20 39 22 41
rect 39 39 41 41
rect 55 39 57 41
<< ndifct0 >>
rect 26 26 28 28
rect 26 19 28 21
rect 36 18 38 20
<< ndifct1 >>
rect 15 23 17 25
rect 15 16 17 18
rect 58 25 60 27
rect 58 18 60 20
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
<< pdifct1 >>
rect 14 70 16 72
rect 14 63 16 65
rect 26 59 28 61
rect 26 52 28 54
rect 36 70 38 72
rect 47 56 49 58
rect 47 48 49 50
rect 58 70 60 72
rect 58 63 60 65
<< alu0 >>
rect 5 81 13 82
rect 5 79 7 81
rect 9 79 13 81
rect 5 78 13 79
rect 25 28 29 30
rect 25 26 26 28
rect 28 26 29 28
rect 25 21 29 26
rect 25 19 26 21
rect 28 20 40 21
rect 28 19 36 20
rect 25 18 36 19
rect 38 18 40 20
rect 25 17 40 18
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 14 79 16 81
rect 36 79 38 81
rect 58 79 60 81
rect 15 7 17 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
<< labels >>
rlabel alu1 16 44 16 44 6 a
rlabel alu1 24 60 24 60 6 z
rlabel alu1 40 36 40 36 6 b
rlabel alu1 32 60 32 60 6 z
rlabel alu1 40 60 40 60 6 z
rlabel alu1 56 20 56 20 6 z
rlabel alu1 56 44 56 44 6 c
rlabel alu1 48 44 48 44 6 z
rlabel alu2 32 6 32 6 6 vss
rlabel alu2 32 82 32 82 6 vdd
<< end >>
