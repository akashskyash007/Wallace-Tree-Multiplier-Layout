magic
tech scmos
timestamp 1199201862
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 41 66 43 70
rect 9 29 11 39
rect 19 36 21 39
rect 19 34 25 36
rect 19 32 21 34
rect 23 32 25 34
rect 19 30 25 32
rect 29 35 31 39
rect 29 33 35 35
rect 29 31 31 33
rect 33 31 35 33
rect 9 27 15 29
rect 9 25 11 27
rect 13 25 15 27
rect 9 23 15 25
rect 12 19 14 23
rect 20 19 22 30
rect 29 29 35 31
rect 30 19 32 29
rect 41 28 43 39
rect 41 26 47 28
rect 41 24 43 26
rect 45 24 47 26
rect 38 22 47 24
rect 38 19 40 22
rect 12 2 14 7
rect 20 2 22 7
rect 30 2 32 7
rect 38 2 40 7
<< ndif >>
rect 3 7 12 19
rect 14 7 20 19
rect 22 16 30 19
rect 22 14 25 16
rect 27 14 30 16
rect 22 7 30 14
rect 32 7 38 19
rect 40 11 48 19
rect 40 9 43 11
rect 45 9 48 11
rect 40 7 48 9
rect 3 5 6 7
rect 8 5 10 7
rect 3 3 10 5
<< pdif >>
rect 4 59 9 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 53 9 55
rect 4 39 9 53
rect 11 50 19 66
rect 11 48 14 50
rect 16 48 19 50
rect 11 39 19 48
rect 21 57 29 66
rect 21 55 24 57
rect 26 55 29 57
rect 21 39 29 55
rect 31 64 41 66
rect 31 62 35 64
rect 37 62 41 64
rect 31 39 41 62
rect 43 59 48 66
rect 43 57 50 59
rect 43 55 46 57
rect 48 55 50 57
rect 43 53 50 55
rect 43 39 48 53
<< alu1 >>
rect -2 64 58 72
rect 2 50 18 51
rect 2 48 14 50
rect 16 48 18 50
rect 2 47 18 48
rect 2 19 6 47
rect 26 43 30 51
rect 10 27 14 43
rect 18 37 30 43
rect 34 46 47 50
rect 34 29 38 46
rect 10 25 11 27
rect 13 25 22 27
rect 10 23 22 25
rect 18 21 22 23
rect 26 25 30 27
rect 42 26 46 35
rect 42 25 43 26
rect 26 24 43 25
rect 45 24 46 26
rect 26 21 46 24
rect 2 13 14 19
rect 34 13 38 21
rect -2 7 58 8
rect -2 5 6 7
rect 8 5 58 7
rect -2 0 58 5
<< nmos >>
rect 12 7 14 19
rect 20 7 22 19
rect 30 7 32 19
rect 38 7 40 19
<< pmos >>
rect 9 39 11 66
rect 19 39 21 66
rect 29 39 31 66
rect 41 39 43 66
<< polyct0 >>
rect 21 32 23 34
rect 31 31 33 33
<< polyct1 >>
rect 11 25 13 27
rect 43 24 45 26
<< ndifct0 >>
rect 25 14 27 16
rect 43 9 45 11
<< ndifct1 >>
rect 6 5 8 7
<< pdifct0 >>
rect 4 55 6 57
rect 24 55 26 57
rect 35 62 37 64
rect 46 55 48 57
<< pdifct1 >>
rect 14 48 16 50
<< alu0 >>
rect 33 62 35 64
rect 37 62 39 64
rect 33 61 39 62
rect 2 57 50 58
rect 2 55 4 57
rect 6 55 24 57
rect 26 55 46 57
rect 48 55 50 57
rect 2 54 50 55
rect 20 34 24 37
rect 20 32 21 34
rect 23 32 24 34
rect 20 30 24 32
rect 29 33 34 34
rect 29 31 31 33
rect 33 31 34 33
rect 29 30 34 31
rect 14 16 29 17
rect 14 14 25 16
rect 27 14 29 16
rect 14 13 29 14
rect 42 11 46 13
rect 42 9 43 11
rect 45 9 46 11
rect 42 8 46 9
<< labels >>
rlabel alu0 26 56 26 56 6 n3
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 24 20 24 6 b1
rlabel alu1 20 40 20 40 6 b2
rlabel alu1 12 36 12 36 6 b1
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 16 36 16 6 a1
rlabel alu1 28 24 28 24 6 a1
rlabel alu1 36 36 36 36 6 a2
rlabel alu1 28 44 28 44 6 b2
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 28 44 28 6 a1
rlabel alu1 44 48 44 48 6 a2
<< end >>
