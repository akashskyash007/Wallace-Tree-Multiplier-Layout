magic
tech scmos
timestamp 1199202985
<< ab >>
rect 0 0 152 80
<< nwell >>
rect -5 36 157 88
<< pwell >>
rect -5 -8 157 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 84 70 86 74
rect 94 70 96 74
rect 101 70 103 74
rect 111 63 113 68
rect 118 63 120 68
rect 128 58 130 63
rect 135 58 137 63
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 16 37 29 39
rect 23 35 25 37
rect 27 35 29 37
rect 23 33 29 35
rect 33 37 45 39
rect 49 37 62 39
rect 67 39 69 42
rect 77 39 79 42
rect 84 39 86 42
rect 94 39 96 42
rect 67 37 80 39
rect 84 37 96 39
rect 33 35 35 37
rect 37 35 39 37
rect 33 33 39 35
rect 49 35 51 37
rect 53 35 62 37
rect 49 33 62 35
rect 73 35 75 37
rect 77 35 80 37
rect 73 33 80 35
rect 9 31 16 33
rect 9 29 12 31
rect 14 29 16 31
rect 27 30 29 33
rect 37 30 39 33
rect 50 30 52 33
rect 60 30 62 33
rect 78 30 80 33
rect 88 35 91 37
rect 93 35 96 37
rect 88 33 96 35
rect 101 39 103 42
rect 111 39 113 42
rect 101 37 113 39
rect 101 35 107 37
rect 109 35 113 37
rect 101 33 113 35
rect 118 39 120 42
rect 128 39 130 42
rect 118 37 130 39
rect 118 35 123 37
rect 125 35 130 37
rect 118 33 130 35
rect 135 39 137 42
rect 135 37 143 39
rect 135 35 139 37
rect 141 35 143 37
rect 135 33 143 35
rect 88 30 90 33
rect 101 30 103 33
rect 111 30 113 33
rect 125 30 127 33
rect 135 30 137 33
rect 9 27 16 29
rect 27 6 29 10
rect 37 6 39 10
rect 50 6 52 10
rect 60 6 62 10
rect 78 6 80 10
rect 88 6 90 10
rect 101 6 103 10
rect 111 6 113 10
rect 125 6 127 10
rect 135 6 137 10
<< ndif >>
rect 19 11 27 30
rect 19 9 21 11
rect 23 10 27 11
rect 29 21 37 30
rect 29 19 32 21
rect 34 19 37 21
rect 29 10 37 19
rect 39 11 50 30
rect 39 10 43 11
rect 23 9 25 10
rect 19 7 25 9
rect 41 9 43 10
rect 45 10 50 11
rect 52 21 60 30
rect 52 19 55 21
rect 57 19 60 21
rect 52 10 60 19
rect 62 11 78 30
rect 62 10 69 11
rect 45 9 48 10
rect 41 7 48 9
rect 64 9 69 10
rect 71 10 78 11
rect 80 21 88 30
rect 80 19 83 21
rect 85 19 88 21
rect 80 10 88 19
rect 90 11 101 30
rect 90 10 94 11
rect 71 9 76 10
rect 64 7 76 9
rect 92 9 94 10
rect 96 10 101 11
rect 103 21 111 30
rect 103 19 106 21
rect 108 19 111 21
rect 103 10 111 19
rect 113 11 125 30
rect 113 10 118 11
rect 96 9 99 10
rect 92 7 99 9
rect 115 9 118 10
rect 120 10 125 11
rect 127 21 135 30
rect 127 19 130 21
rect 132 19 135 21
rect 127 10 135 19
rect 137 21 146 30
rect 137 19 141 21
rect 143 19 146 21
rect 137 14 146 19
rect 137 12 141 14
rect 143 12 146 14
rect 137 10 146 12
rect 120 9 123 10
rect 115 7 123 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 42 16 70
rect 18 61 26 70
rect 18 59 21 61
rect 23 59 26 61
rect 18 53 26 59
rect 18 51 21 53
rect 23 51 26 53
rect 18 42 26 51
rect 28 42 33 70
rect 35 68 43 70
rect 35 66 38 68
rect 40 66 43 68
rect 35 61 43 66
rect 35 59 38 61
rect 40 59 43 61
rect 35 42 43 59
rect 45 42 50 70
rect 52 60 60 70
rect 52 58 55 60
rect 57 58 60 60
rect 52 53 60 58
rect 52 51 55 53
rect 57 51 60 53
rect 52 42 60 51
rect 62 42 67 70
rect 69 68 77 70
rect 69 66 72 68
rect 74 66 77 68
rect 69 61 77 66
rect 69 59 72 61
rect 74 59 77 61
rect 69 42 77 59
rect 79 42 84 70
rect 86 61 94 70
rect 86 59 89 61
rect 91 59 94 61
rect 86 53 94 59
rect 86 51 89 53
rect 91 51 94 53
rect 86 42 94 51
rect 96 42 101 70
rect 103 63 109 70
rect 103 61 111 63
rect 103 59 106 61
rect 108 59 111 61
rect 103 42 111 59
rect 113 42 118 63
rect 120 58 125 63
rect 120 53 128 58
rect 120 51 123 53
rect 125 51 128 53
rect 120 42 128 51
rect 130 42 135 58
rect 137 56 145 58
rect 137 54 140 56
rect 142 54 145 56
rect 137 42 145 54
<< alu1 >>
rect -2 81 154 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 154 81
rect -2 68 154 79
rect 18 61 24 63
rect 18 59 21 61
rect 23 59 24 61
rect 18 54 24 59
rect 54 60 58 62
rect 54 58 55 60
rect 57 58 58 60
rect 88 61 94 63
rect 88 59 89 61
rect 91 59 94 61
rect 54 54 58 58
rect 88 54 94 59
rect 2 53 127 54
rect 2 51 21 53
rect 23 51 55 53
rect 57 51 89 53
rect 91 51 123 53
rect 125 51 127 53
rect 2 50 127 51
rect 2 22 6 50
rect 23 42 127 46
rect 23 37 29 42
rect 23 35 25 37
rect 27 35 29 37
rect 23 34 29 35
rect 33 37 39 38
rect 33 35 35 37
rect 37 35 39 37
rect 11 31 15 33
rect 11 29 12 31
rect 14 30 15 31
rect 33 30 39 35
rect 49 37 55 42
rect 49 35 51 37
rect 53 35 55 37
rect 49 34 55 35
rect 73 37 79 38
rect 73 35 75 37
rect 77 35 79 37
rect 73 30 79 35
rect 89 37 95 42
rect 89 35 91 37
rect 93 35 95 37
rect 89 34 95 35
rect 105 37 111 38
rect 105 35 107 37
rect 109 35 111 37
rect 105 30 111 35
rect 121 37 127 42
rect 121 35 123 37
rect 125 35 127 37
rect 121 34 127 35
rect 137 37 143 38
rect 137 35 139 37
rect 141 35 143 37
rect 137 30 143 35
rect 14 29 143 30
rect 11 26 143 29
rect 2 21 135 22
rect 2 19 32 21
rect 34 19 55 21
rect 57 19 83 21
rect 85 19 106 21
rect 108 19 130 21
rect 132 19 135 21
rect 2 18 135 19
rect -2 11 154 12
rect -2 9 21 11
rect 23 9 43 11
rect 45 9 69 11
rect 71 9 94 11
rect 96 9 118 11
rect 120 9 154 11
rect -2 1 154 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 154 1
rect -2 -2 154 -1
<< ptie >>
rect 0 1 152 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 152 1
rect 0 -3 152 -1
<< ntie >>
rect 0 81 152 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 152 81
rect 0 77 152 79
<< nmos >>
rect 27 10 29 30
rect 37 10 39 30
rect 50 10 52 30
rect 60 10 62 30
rect 78 10 80 30
rect 88 10 90 30
rect 101 10 103 30
rect 111 10 113 30
rect 125 10 127 30
rect 135 10 137 30
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 84 42 86 70
rect 94 42 96 70
rect 101 42 103 70
rect 111 42 113 63
rect 118 42 120 63
rect 128 42 130 58
rect 135 42 137 58
<< polyct1 >>
rect 25 35 27 37
rect 35 35 37 37
rect 51 35 53 37
rect 75 35 77 37
rect 12 29 14 31
rect 91 35 93 37
rect 107 35 109 37
rect 123 35 125 37
rect 139 35 141 37
<< ndifct0 >>
rect 141 19 143 21
rect 141 12 143 14
<< ndifct1 >>
rect 21 9 23 11
rect 32 19 34 21
rect 43 9 45 11
rect 55 19 57 21
rect 69 9 71 11
rect 83 19 85 21
rect 94 9 96 11
rect 106 19 108 21
rect 118 9 120 11
rect 130 19 132 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 38 66 40 68
rect 38 59 40 61
rect 72 66 74 68
rect 72 59 74 61
rect 106 59 108 61
rect 140 54 142 56
<< pdifct1 >>
rect 21 59 23 61
rect 21 51 23 53
rect 55 58 57 60
rect 55 51 57 53
rect 89 59 91 61
rect 89 51 91 53
rect 123 51 125 53
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 36 66 38 68
rect 40 66 42 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 36 61 42 66
rect 70 66 72 68
rect 74 66 76 68
rect 36 59 38 61
rect 40 59 42 61
rect 36 58 42 59
rect 70 61 76 66
rect 70 59 72 61
rect 74 59 76 61
rect 70 58 76 59
rect 104 61 110 68
rect 104 59 106 61
rect 108 59 110 61
rect 104 58 110 59
rect 139 56 143 68
rect 139 54 140 56
rect 142 54 143 56
rect 139 52 143 54
rect 139 21 145 22
rect 139 19 141 21
rect 143 19 145 21
rect 139 14 145 19
rect 139 12 141 14
rect 143 12 145 14
<< labels >>
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 52 28 52 28 6 a
rlabel alu1 52 20 52 20 6 z
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 32 36 32 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 52 40 52 40 6 b
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 76 6 76 6 6 vss
rlabel alu1 60 20 60 20 6 z
rlabel alu1 60 28 60 28 6 a
rlabel alu1 84 28 84 28 6 a
rlabel ndifct1 84 20 84 20 6 z
rlabel alu1 76 20 76 20 6 z
rlabel alu1 68 28 68 28 6 a
rlabel alu1 68 20 68 20 6 z
rlabel alu1 76 32 76 32 6 a
rlabel alu1 60 44 60 44 6 b
rlabel alu1 76 44 76 44 6 b
rlabel alu1 84 44 84 44 6 b
rlabel alu1 68 44 68 44 6 b
rlabel alu1 68 52 68 52 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 76 74 76 74 6 vdd
rlabel alu1 92 20 92 20 6 z
rlabel alu1 92 28 92 28 6 a
rlabel alu1 116 28 116 28 6 a
rlabel alu1 116 20 116 20 6 z
rlabel alu1 108 20 108 20 6 z
rlabel alu1 100 28 100 28 6 a
rlabel alu1 100 20 100 20 6 z
rlabel alu1 108 32 108 32 6 a
rlabel alu1 92 40 92 40 6 b
rlabel alu1 108 44 108 44 6 b
rlabel alu1 116 44 116 44 6 b
rlabel alu1 100 44 100 44 6 b
rlabel alu1 100 52 100 52 6 z
rlabel alu1 108 52 108 52 6 z
rlabel alu1 116 52 116 52 6 z
rlabel alu1 92 56 92 56 6 z
rlabel alu1 124 20 124 20 6 z
rlabel alu1 124 28 124 28 6 a
rlabel alu1 132 28 132 28 6 a
rlabel alu1 132 20 132 20 6 z
rlabel alu1 140 32 140 32 6 a
rlabel alu1 124 40 124 40 6 b
rlabel pdifct1 124 52 124 52 6 z
<< end >>
