magic
tech scmos
timestamp 1199203432
<< ab >>
rect 0 0 144 72
<< nwell >>
rect -5 32 149 77
<< pwell >>
rect -5 -5 149 32
<< poly >>
rect 18 65 20 70
rect 28 65 30 70
rect 38 68 50 70
rect 38 65 40 68
rect 48 65 50 68
rect 69 66 71 70
rect 79 66 81 70
rect 91 66 93 70
rect 101 66 103 70
rect 118 66 120 70
rect 128 66 130 70
rect 2 35 8 37
rect 18 35 20 38
rect 28 35 30 38
rect 38 35 40 38
rect 2 33 4 35
rect 6 33 8 35
rect 16 33 31 35
rect 2 31 11 33
rect 9 26 11 31
rect 16 26 18 33
rect 25 31 27 33
rect 29 31 31 33
rect 25 29 31 31
rect 35 33 41 35
rect 48 34 50 38
rect 69 35 71 38
rect 79 35 81 38
rect 91 35 93 38
rect 101 35 103 38
rect 69 33 87 35
rect 35 31 37 33
rect 39 31 41 33
rect 81 31 83 33
rect 85 31 87 33
rect 35 29 41 31
rect 28 26 30 29
rect 35 26 37 29
rect 45 26 47 30
rect 55 26 57 31
rect 81 29 87 31
rect 91 33 104 35
rect 91 31 99 33
rect 101 31 104 33
rect 91 29 104 31
rect 108 33 114 35
rect 108 31 110 33
rect 112 31 114 33
rect 118 34 120 38
rect 128 35 130 38
rect 118 31 121 34
rect 108 29 114 31
rect 85 26 87 29
rect 92 26 94 29
rect 102 26 104 29
rect 109 26 111 29
rect 119 26 121 31
rect 128 33 135 35
rect 128 31 131 33
rect 133 31 135 33
rect 128 29 135 31
rect 129 26 131 29
rect 9 14 11 19
rect 16 14 18 19
rect 85 8 87 12
rect 92 8 94 12
rect 102 8 104 12
rect 109 8 111 12
rect 28 2 30 7
rect 35 2 37 7
rect 45 4 47 7
rect 55 4 57 7
rect 119 4 121 12
rect 129 4 131 12
rect 45 2 131 4
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 19 9 22
rect 11 19 16 26
rect 18 19 28 26
rect 20 9 28 19
rect 20 7 22 9
rect 24 7 28 9
rect 30 7 35 26
rect 37 17 45 26
rect 37 15 40 17
rect 42 15 45 17
rect 37 7 45 15
rect 47 24 55 26
rect 47 22 50 24
rect 52 22 55 24
rect 47 7 55 22
rect 57 19 62 26
rect 57 17 64 19
rect 57 15 60 17
rect 62 15 64 17
rect 57 13 64 15
rect 57 7 62 13
rect 78 16 85 26
rect 78 14 80 16
rect 82 14 85 16
rect 78 12 85 14
rect 87 12 92 26
rect 94 17 102 26
rect 94 15 97 17
rect 99 15 102 17
rect 94 12 102 15
rect 104 12 109 26
rect 111 16 119 26
rect 111 14 114 16
rect 116 14 119 16
rect 111 12 119 14
rect 121 24 129 26
rect 121 22 124 24
rect 126 22 129 24
rect 121 17 129 22
rect 121 15 124 17
rect 126 15 129 17
rect 121 12 129 15
rect 131 23 138 26
rect 131 21 134 23
rect 136 21 138 23
rect 131 16 138 21
rect 131 14 134 16
rect 136 14 138 16
rect 131 12 138 14
rect 20 5 26 7
<< pdif >>
rect 13 51 18 65
rect 11 49 18 51
rect 11 47 13 49
rect 15 47 18 49
rect 11 42 18 47
rect 11 40 13 42
rect 15 40 18 42
rect 11 38 18 40
rect 20 57 28 65
rect 20 55 23 57
rect 25 55 28 57
rect 20 38 28 55
rect 30 49 38 65
rect 30 47 33 49
rect 35 47 38 49
rect 30 38 38 47
rect 40 42 48 65
rect 40 40 43 42
rect 45 40 48 42
rect 40 38 48 40
rect 50 51 55 65
rect 62 64 69 66
rect 62 62 64 64
rect 66 62 69 64
rect 50 49 57 51
rect 50 47 53 49
rect 55 47 57 49
rect 50 42 57 47
rect 50 40 53 42
rect 55 40 57 42
rect 50 38 57 40
rect 62 38 69 62
rect 71 49 79 66
rect 71 47 74 49
rect 76 47 79 49
rect 71 42 79 47
rect 71 40 74 42
rect 76 40 79 42
rect 71 38 79 40
rect 81 64 91 66
rect 81 62 85 64
rect 87 62 91 64
rect 81 38 91 62
rect 93 49 101 66
rect 93 47 96 49
rect 98 47 101 49
rect 93 38 101 47
rect 103 64 118 66
rect 103 62 106 64
rect 108 62 113 64
rect 115 62 118 64
rect 103 57 118 62
rect 103 55 113 57
rect 115 55 118 57
rect 103 38 118 55
rect 120 42 128 66
rect 120 40 123 42
rect 125 40 128 42
rect 120 38 128 40
rect 130 64 138 66
rect 130 62 134 64
rect 136 62 138 64
rect 130 38 138 62
<< alu1 >>
rect -2 67 146 72
rect -2 65 5 67
rect 7 65 146 67
rect -2 64 146 65
rect 121 54 134 58
rect 10 49 57 50
rect 10 47 13 49
rect 15 47 33 49
rect 35 47 53 49
rect 55 47 57 49
rect 10 46 57 47
rect 10 42 16 46
rect 10 40 13 42
rect 15 40 16 42
rect 10 38 16 40
rect 52 42 57 46
rect 52 40 53 42
rect 55 40 57 42
rect 52 38 57 40
rect 10 27 14 38
rect 2 24 14 27
rect 2 22 4 24
rect 6 22 14 24
rect 81 38 119 42
rect 81 33 87 38
rect 81 31 83 33
rect 85 31 87 33
rect 81 30 87 31
rect 97 33 103 34
rect 97 31 99 33
rect 101 31 103 33
rect 97 26 103 31
rect 130 33 134 54
rect 130 31 131 33
rect 133 31 134 33
rect 130 29 134 31
rect 97 22 111 26
rect 2 21 14 22
rect 9 18 14 21
rect 9 17 64 18
rect 9 15 40 17
rect 42 15 60 17
rect 62 15 64 17
rect 9 14 64 15
rect -2 7 22 8
rect 24 7 146 8
rect -2 5 5 7
rect 7 5 12 7
rect 14 5 146 7
rect -2 0 146 5
<< ptie >>
rect 3 7 16 9
rect 3 5 5 7
rect 7 5 12 7
rect 14 5 16 7
rect 68 10 74 26
rect 68 8 70 10
rect 72 8 74 10
rect 3 3 16 5
rect 68 6 74 8
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 56 9 65
<< nmos >>
rect 9 19 11 26
rect 16 19 18 26
rect 28 7 30 26
rect 35 7 37 26
rect 45 7 47 26
rect 55 7 57 26
rect 85 12 87 26
rect 92 12 94 26
rect 102 12 104 26
rect 109 12 111 26
rect 119 12 121 26
rect 129 12 131 26
<< pmos >>
rect 18 38 20 65
rect 28 38 30 65
rect 38 38 40 65
rect 48 38 50 65
rect 69 38 71 66
rect 79 38 81 66
rect 91 38 93 66
rect 101 38 103 66
rect 118 38 120 66
rect 128 38 130 66
<< polyct0 >>
rect 4 33 6 35
rect 27 31 29 33
rect 37 31 39 33
rect 110 31 112 33
<< polyct1 >>
rect 83 31 85 33
rect 99 31 101 33
rect 131 31 133 33
<< ndifct0 >>
rect 22 8 24 9
rect 50 22 52 24
rect 80 14 82 16
rect 97 15 99 17
rect 114 14 116 16
rect 124 22 126 24
rect 124 15 126 17
rect 134 21 136 23
rect 134 14 136 16
<< ndifct1 >>
rect 4 22 6 24
rect 22 7 24 8
rect 40 15 42 17
rect 60 15 62 17
<< ntiect1 >>
rect 5 65 7 67
<< ptiect0 >>
rect 70 8 72 10
<< ptiect1 >>
rect 5 5 7 7
rect 12 5 14 7
<< pdifct0 >>
rect 23 55 25 57
rect 43 40 45 42
rect 64 62 66 64
rect 74 47 76 49
rect 74 40 76 42
rect 85 62 87 64
rect 96 47 98 49
rect 106 62 108 64
rect 113 62 115 64
rect 113 55 115 57
rect 123 40 125 42
rect 134 62 136 64
<< pdifct1 >>
rect 13 47 15 49
rect 13 40 15 42
rect 33 47 35 49
rect 53 47 55 49
rect 53 40 55 42
<< alu0 >>
rect 62 62 64 64
rect 66 62 68 64
rect 62 61 68 62
rect 83 62 85 64
rect 87 62 89 64
rect 83 61 89 62
rect 103 62 106 64
rect 108 62 113 64
rect 115 62 117 64
rect 103 61 117 62
rect 132 62 134 64
rect 136 62 138 64
rect 132 61 138 62
rect 2 57 107 58
rect 2 55 23 57
rect 25 55 107 57
rect 2 54 107 55
rect 111 57 117 61
rect 111 55 113 57
rect 115 55 117 57
rect 111 54 117 55
rect 2 37 6 54
rect 41 42 47 43
rect 26 40 43 42
rect 45 40 47 42
rect 26 38 47 40
rect 2 35 7 37
rect 2 33 4 35
rect 6 33 7 35
rect 2 31 7 33
rect 26 33 30 38
rect 61 34 65 54
rect 103 50 107 54
rect 26 31 27 33
rect 29 31 30 33
rect 26 26 30 31
rect 35 33 65 34
rect 35 31 37 33
rect 39 31 65 33
rect 35 30 65 31
rect 72 49 100 50
rect 72 47 74 49
rect 76 47 96 49
rect 98 47 100 49
rect 72 46 100 47
rect 103 46 126 50
rect 72 42 77 46
rect 122 42 126 46
rect 72 40 74 42
rect 76 40 77 42
rect 72 26 77 40
rect 122 40 123 42
rect 125 40 126 42
rect 108 33 114 38
rect 108 31 110 33
rect 112 31 114 33
rect 108 30 114 31
rect 122 26 126 40
rect 26 24 92 26
rect 26 22 50 24
rect 52 22 92 24
rect 122 24 127 26
rect 122 22 124 24
rect 126 22 127 24
rect 48 21 54 22
rect 88 18 92 22
rect 88 17 101 18
rect 78 16 84 17
rect 78 14 80 16
rect 82 14 84 16
rect 88 15 97 17
rect 99 15 101 17
rect 88 14 101 15
rect 113 16 117 18
rect 113 14 114 16
rect 116 14 117 16
rect 69 10 73 12
rect 20 9 26 10
rect 20 8 22 9
rect 24 8 26 9
rect 69 8 70 10
rect 72 8 73 10
rect 78 8 84 14
rect 113 8 117 14
rect 122 17 127 22
rect 122 15 124 17
rect 126 15 127 17
rect 122 13 127 15
rect 133 23 137 25
rect 133 21 134 23
rect 136 21 137 23
rect 133 16 137 21
rect 133 14 134 16
rect 136 14 137 16
rect 133 8 137 14
<< labels >>
rlabel polyct0 28 32 28 32 6 an
rlabel alu0 4 44 4 44 6 bn
rlabel alu0 50 32 50 32 6 bn
rlabel alu0 44 40 44 40 6 an
rlabel alu0 94 16 94 16 6 an
rlabel alu0 59 24 59 24 6 an
rlabel alu0 74 36 74 36 6 an
rlabel alu0 86 48 86 48 6 an
rlabel alu0 124 31 124 31 6 bn
rlabel alu0 54 56 54 56 6 bn
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 4 24 4 24 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 60 16 60 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 72 4 72 4 6 vss
rlabel alu1 100 28 100 28 6 a1
rlabel alu1 84 36 84 36 6 a2
rlabel alu1 100 40 100 40 6 a2
rlabel alu1 92 40 92 40 6 a2
rlabel alu1 72 68 72 68 6 vdd
rlabel alu1 108 24 108 24 6 a1
rlabel alu1 116 40 116 40 6 a2
rlabel alu1 132 40 132 40 6 b
rlabel alu1 108 40 108 40 6 a2
rlabel alu1 124 56 124 56 6 b
<< end >>
