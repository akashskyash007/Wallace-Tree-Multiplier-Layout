magic
tech scmos
timestamp 1199202097
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 25 72 110 74
rect 15 63 17 68
rect 25 64 27 72
rect 56 69 58 72
rect 35 64 37 68
rect 77 64 79 68
rect 87 64 89 72
rect 97 64 99 68
rect 56 44 58 47
rect 56 42 61 44
rect 15 39 17 42
rect 2 37 17 39
rect 25 39 27 42
rect 25 37 30 39
rect 2 35 4 37
rect 6 35 17 37
rect 2 33 17 35
rect 12 26 14 33
rect 28 31 30 37
rect 35 38 37 42
rect 59 40 61 42
rect 59 38 65 40
rect 77 39 79 42
rect 35 36 55 38
rect 43 34 51 36
rect 53 34 55 36
rect 43 32 55 34
rect 59 36 61 38
rect 63 36 65 38
rect 59 34 65 36
rect 73 37 79 39
rect 87 37 89 42
rect 97 39 99 42
rect 94 37 99 39
rect 73 35 75 37
rect 77 35 79 37
rect 22 26 24 31
rect 28 29 34 31
rect 32 26 34 29
rect 12 11 14 16
rect 22 8 24 16
rect 32 12 34 16
rect 43 8 45 32
rect 59 30 61 34
rect 73 33 79 35
rect 94 33 96 37
rect 108 33 110 72
rect 73 31 83 33
rect 81 28 83 31
rect 91 31 96 33
rect 101 31 110 33
rect 91 28 93 31
rect 101 28 103 31
rect 59 15 61 20
rect 81 13 83 18
rect 91 8 93 18
rect 101 13 103 18
rect 22 6 93 8
<< ndif >>
rect 3 20 12 26
rect 3 18 6 20
rect 8 18 12 20
rect 3 16 12 18
rect 14 24 22 26
rect 14 22 17 24
rect 19 22 22 24
rect 14 16 22 22
rect 24 24 32 26
rect 24 22 27 24
rect 29 22 32 24
rect 24 16 32 22
rect 34 23 39 26
rect 34 21 41 23
rect 34 19 37 21
rect 39 19 41 21
rect 34 16 41 19
rect 52 28 59 30
rect 52 26 54 28
rect 56 26 59 28
rect 52 24 59 26
rect 54 20 59 24
rect 61 28 66 30
rect 61 22 81 28
rect 61 20 72 22
rect 74 20 81 22
rect 63 18 81 20
rect 83 26 91 28
rect 83 24 86 26
rect 88 24 91 26
rect 83 18 91 24
rect 93 22 101 28
rect 93 20 96 22
rect 98 20 101 22
rect 93 18 101 20
rect 103 26 110 28
rect 103 24 106 26
rect 108 24 110 26
rect 103 22 110 24
rect 103 18 108 22
<< pdif >>
rect 20 63 25 64
rect 7 61 15 63
rect 7 59 10 61
rect 12 59 15 61
rect 7 54 15 59
rect 7 52 10 54
rect 12 52 15 54
rect 7 42 15 52
rect 17 53 25 63
rect 17 51 20 53
rect 22 51 25 53
rect 17 46 25 51
rect 17 44 20 46
rect 22 44 25 46
rect 17 42 25 44
rect 27 53 35 64
rect 27 51 30 53
rect 32 51 35 53
rect 27 46 35 51
rect 27 44 30 46
rect 32 44 35 46
rect 27 42 35 44
rect 37 55 42 64
rect 37 53 44 55
rect 51 53 56 69
rect 37 51 40 53
rect 42 51 44 53
rect 37 46 44 51
rect 49 51 56 53
rect 49 49 51 51
rect 53 49 56 51
rect 49 47 56 49
rect 58 67 75 69
rect 58 65 64 67
rect 66 65 75 67
rect 58 64 75 65
rect 58 47 77 64
rect 37 44 40 46
rect 42 44 44 46
rect 37 42 44 44
rect 67 42 77 47
rect 79 53 87 64
rect 79 51 82 53
rect 84 51 87 53
rect 79 46 87 51
rect 79 44 82 46
rect 84 44 87 46
rect 79 42 87 44
rect 89 53 97 64
rect 89 51 92 53
rect 94 51 97 53
rect 89 46 97 51
rect 89 44 92 46
rect 94 44 97 46
rect 89 42 97 44
rect 99 62 106 64
rect 99 60 102 62
rect 104 60 106 62
rect 99 55 106 60
rect 99 53 102 55
rect 104 53 106 55
rect 99 51 106 53
rect 99 42 104 51
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 68 114 79
rect 2 41 14 47
rect 2 37 7 41
rect 2 35 4 37
rect 6 35 7 37
rect 2 25 7 35
rect 26 53 33 55
rect 26 51 30 53
rect 32 51 33 53
rect 26 46 33 51
rect 26 44 30 46
rect 32 44 33 46
rect 26 42 33 44
rect 26 31 30 42
rect 65 50 78 54
rect 26 25 38 31
rect 26 24 30 25
rect 26 22 27 24
rect 29 22 30 24
rect 57 39 63 46
rect 57 38 70 39
rect 57 36 61 38
rect 63 36 70 38
rect 57 33 70 36
rect 74 37 78 50
rect 74 35 75 37
rect 77 35 78 37
rect 74 33 78 35
rect 90 53 95 55
rect 90 51 92 53
rect 94 51 95 53
rect 90 46 95 51
rect 90 44 92 46
rect 94 44 95 46
rect 90 39 95 44
rect 90 33 102 39
rect 26 17 30 22
rect 98 23 102 33
rect 94 22 102 23
rect 94 20 96 22
rect 98 20 102 22
rect 94 17 102 20
rect -2 1 114 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 12 16 14 26
rect 22 16 24 26
rect 32 16 34 26
rect 59 20 61 30
rect 81 18 83 28
rect 91 18 93 28
rect 101 18 103 28
<< pmos >>
rect 15 42 17 63
rect 25 42 27 64
rect 35 42 37 64
rect 56 47 58 69
rect 77 42 79 64
rect 87 42 89 64
rect 97 42 99 64
<< polyct0 >>
rect 51 34 53 36
<< polyct1 >>
rect 4 35 6 37
rect 61 36 63 38
rect 75 35 77 37
<< ndifct0 >>
rect 6 18 8 20
rect 17 22 19 24
rect 37 19 39 21
rect 54 26 56 28
rect 72 20 74 22
rect 86 24 88 26
rect 106 24 108 26
<< ndifct1 >>
rect 27 22 29 24
rect 96 20 98 22
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 10 59 12 61
rect 10 52 12 54
rect 20 51 22 53
rect 20 44 22 46
rect 40 51 42 53
rect 51 49 53 51
rect 64 65 66 67
rect 40 44 42 46
rect 82 51 84 53
rect 82 44 84 46
rect 102 60 104 62
rect 102 53 104 55
<< pdifct1 >>
rect 30 51 32 53
rect 30 44 32 46
rect 92 51 94 53
rect 92 44 94 46
<< alu0 >>
rect 9 61 13 68
rect 62 67 68 68
rect 62 65 64 67
rect 66 65 68 67
rect 62 64 68 65
rect 9 59 10 61
rect 12 59 13 61
rect 9 54 13 59
rect 9 52 10 54
rect 12 52 13 54
rect 9 50 13 52
rect 19 61 52 63
rect 72 62 106 63
rect 72 61 102 62
rect 19 60 102 61
rect 104 60 106 62
rect 19 59 106 60
rect 19 53 23 59
rect 48 57 76 59
rect 100 56 106 59
rect 100 55 109 56
rect 19 51 20 53
rect 22 51 23 53
rect 19 46 23 51
rect 19 44 20 46
rect 22 44 23 46
rect 19 38 23 44
rect 16 34 23 38
rect 39 53 43 55
rect 39 51 40 53
rect 42 51 43 53
rect 39 46 43 51
rect 39 44 40 46
rect 42 44 43 46
rect 16 24 20 34
rect 16 22 17 24
rect 19 22 20 24
rect 4 20 10 21
rect 16 20 20 22
rect 39 39 43 44
rect 50 51 54 53
rect 50 49 51 51
rect 53 49 54 51
rect 39 35 46 39
rect 42 22 46 35
rect 50 36 54 49
rect 50 34 51 36
rect 53 34 54 36
rect 50 29 54 34
rect 81 53 85 55
rect 81 51 82 53
rect 84 51 85 53
rect 81 46 85 51
rect 81 44 82 46
rect 84 44 85 46
rect 81 30 85 44
rect 100 53 102 55
rect 104 53 109 55
rect 100 52 109 53
rect 50 28 58 29
rect 50 26 54 28
rect 56 26 58 28
rect 50 25 58 26
rect 62 26 89 30
rect 62 22 66 26
rect 85 24 86 26
rect 88 24 89 26
rect 4 18 6 20
rect 8 18 10 20
rect 4 12 10 18
rect 35 21 66 22
rect 35 19 37 21
rect 39 19 66 21
rect 35 18 66 19
rect 70 22 76 23
rect 85 22 89 24
rect 105 26 109 52
rect 105 24 106 26
rect 108 24 109 26
rect 105 22 109 24
rect 70 20 72 22
rect 74 20 76 22
rect 47 12 53 15
rect 70 12 76 20
<< labels >>
rlabel alu0 18 29 18 29 6 a0n
rlabel alu0 21 48 21 48 6 a0n
rlabel alu0 52 39 52 39 6 sn
rlabel pdifct0 41 45 41 45 6 a1n
rlabel alu0 50 20 50 20 6 a1n
rlabel alu0 75 28 75 28 6 a1n
rlabel alu0 107 39 107 39 6 a0n
rlabel alu0 83 40 83 40 6 a1n
rlabel alu0 89 61 89 61 6 a0n
rlabel alu1 4 36 4 36 6 a0
rlabel alu1 12 44 12 44 6 a0
rlabel alu1 28 36 28 36 6 z0
rlabel alu1 36 28 36 28 6 z0
rlabel alu1 56 6 56 6 6 vss
rlabel alu1 68 36 68 36 6 s
rlabel alu1 76 40 76 40 6 a1
rlabel alu1 60 40 60 40 6 s
rlabel alu1 68 52 68 52 6 a1
rlabel alu1 56 74 56 74 6 vdd
rlabel alu1 100 28 100 28 6 z1
rlabel alu1 92 44 92 44 6 z1
<< end >>
