magic
tech scmos
timestamp 1199202677
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 14 69 16 74
rect 24 69 26 74
rect 35 61 37 66
rect 45 61 47 65
rect 14 39 16 42
rect 24 39 26 42
rect 35 39 37 42
rect 45 39 47 42
rect 9 37 26 39
rect 9 35 11 37
rect 13 35 26 37
rect 9 33 26 35
rect 24 30 26 33
rect 31 37 47 39
rect 31 35 43 37
rect 45 35 47 37
rect 31 33 47 35
rect 31 30 33 33
rect 24 6 26 11
rect 31 6 33 11
<< ndif >>
rect 17 28 24 30
rect 17 26 19 28
rect 21 26 24 28
rect 17 21 24 26
rect 17 19 19 21
rect 21 19 24 21
rect 17 17 24 19
rect 19 11 24 17
rect 26 11 31 30
rect 33 22 41 30
rect 33 20 36 22
rect 38 20 41 22
rect 33 15 41 20
rect 33 13 36 15
rect 38 13 41 15
rect 33 11 41 13
<< pdif >>
rect 6 67 14 69
rect 6 65 9 67
rect 11 65 14 67
rect 6 60 14 65
rect 6 58 9 60
rect 11 58 14 60
rect 6 42 14 58
rect 16 53 24 69
rect 16 51 19 53
rect 21 51 24 53
rect 16 46 24 51
rect 16 44 19 46
rect 21 44 24 46
rect 16 42 24 44
rect 26 67 33 69
rect 26 65 29 67
rect 31 65 33 67
rect 26 61 33 65
rect 26 60 35 61
rect 26 58 29 60
rect 31 58 35 60
rect 26 42 35 58
rect 37 53 45 61
rect 37 51 40 53
rect 42 51 45 53
rect 37 46 45 51
rect 37 44 40 46
rect 42 44 45 46
rect 37 42 45 44
rect 47 59 54 61
rect 47 57 50 59
rect 52 57 54 59
rect 47 52 54 57
rect 47 50 50 52
rect 52 50 54 52
rect 47 42 54 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 18 53 22 55
rect 18 51 19 53
rect 21 51 22 53
rect 2 39 6 47
rect 18 46 22 51
rect 39 53 43 55
rect 39 51 40 53
rect 42 51 43 53
rect 39 46 43 51
rect 18 44 19 46
rect 21 44 40 46
rect 42 44 43 46
rect 18 42 43 44
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 18 28 22 42
rect 41 37 54 38
rect 41 35 43 37
rect 45 35 54 37
rect 41 34 54 35
rect 18 26 19 28
rect 21 26 22 28
rect 18 21 22 26
rect 50 25 54 34
rect 18 19 19 21
rect 21 19 22 21
rect 18 17 22 19
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 24 11 26 30
rect 31 11 33 30
<< pmos >>
rect 14 42 16 69
rect 24 42 26 69
rect 35 42 37 61
rect 45 42 47 61
<< polyct1 >>
rect 11 35 13 37
rect 43 35 45 37
<< ndifct0 >>
rect 36 20 38 22
rect 36 13 38 15
<< ndifct1 >>
rect 19 26 21 28
rect 19 19 21 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 9 65 11 67
rect 9 58 11 60
rect 29 65 31 67
rect 29 58 31 60
rect 50 57 52 59
rect 50 50 52 52
<< pdifct1 >>
rect 19 51 21 53
rect 19 44 21 46
rect 40 51 42 53
rect 40 44 42 46
<< alu0 >>
rect 8 67 12 68
rect 8 65 9 67
rect 11 65 12 67
rect 8 60 12 65
rect 8 58 9 60
rect 11 58 12 60
rect 8 56 12 58
rect 28 67 32 68
rect 28 65 29 67
rect 31 65 32 67
rect 28 60 32 65
rect 28 58 29 60
rect 31 58 32 60
rect 28 56 32 58
rect 49 59 53 68
rect 49 57 50 59
rect 52 57 53 59
rect 49 52 53 57
rect 49 50 50 52
rect 52 50 53 52
rect 49 48 53 50
rect 35 22 39 24
rect 35 20 36 22
rect 38 20 39 22
rect 35 15 39 20
rect 35 13 36 15
rect 38 13 39 15
rect 35 12 39 13
<< labels >>
rlabel alu1 4 40 4 40 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 36 20 36 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 44 36 44 6 z
rlabel alu1 28 44 28 44 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 36 44 36 6 a
rlabel alu1 52 28 52 28 6 a
<< end >>
