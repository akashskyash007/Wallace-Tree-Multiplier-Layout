magic
tech scmos
timestamp 1199202639
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 9 67 11 72
rect 19 67 21 72
rect 9 30 11 50
rect 19 47 21 50
rect 19 45 31 47
rect 25 43 27 45
rect 29 43 31 45
rect 25 41 31 43
rect 26 35 28 41
rect 35 37 41 39
rect 35 36 37 37
rect 16 33 28 35
rect 16 30 18 33
rect 26 30 28 33
rect 33 35 37 36
rect 39 35 41 37
rect 33 33 41 35
rect 33 30 35 33
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
<< ndif >>
rect 2 27 9 30
rect 2 25 4 27
rect 6 25 9 27
rect 2 20 9 25
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 16 30
rect 18 28 26 30
rect 18 26 21 28
rect 23 26 26 28
rect 18 21 26 26
rect 18 19 21 21
rect 23 19 26 21
rect 18 16 26 19
rect 28 16 33 30
rect 35 27 43 30
rect 35 25 38 27
rect 40 25 43 27
rect 35 20 43 25
rect 35 18 38 20
rect 40 18 43 20
rect 35 16 43 18
<< pdif >>
rect 2 65 9 67
rect 2 63 4 65
rect 6 63 9 65
rect 2 58 9 63
rect 2 56 4 58
rect 6 56 9 58
rect 2 50 9 56
rect 11 54 19 67
rect 11 52 14 54
rect 16 52 19 54
rect 11 50 19 52
rect 21 65 29 67
rect 21 63 24 65
rect 26 63 29 65
rect 21 50 29 63
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 10 54 18 55
rect 10 52 14 54
rect 16 52 18 54
rect 10 51 18 52
rect 10 31 14 51
rect 26 49 38 55
rect 26 45 30 49
rect 26 43 27 45
rect 29 43 30 45
rect 26 41 30 43
rect 42 39 46 47
rect 34 37 46 39
rect 34 35 37 37
rect 39 35 46 37
rect 34 33 46 35
rect 10 28 24 31
rect 10 27 21 28
rect 18 26 21 27
rect 23 26 24 28
rect 18 21 24 26
rect 18 19 21 21
rect 23 19 24 21
rect 18 17 24 19
rect -2 1 50 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 9 16 11 30
rect 16 16 18 30
rect 26 16 28 30
rect 33 16 35 30
<< pmos >>
rect 9 50 11 67
rect 19 50 21 67
<< polyct1 >>
rect 27 43 29 45
rect 37 35 39 37
<< ndifct0 >>
rect 4 25 6 27
rect 4 18 6 20
rect 38 25 40 27
rect 38 18 40 20
<< ndifct1 >>
rect 21 26 23 28
rect 21 19 23 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 4 63 6 65
rect 4 56 6 58
rect 24 63 26 65
<< pdifct1 >>
rect 14 52 16 54
<< alu0 >>
rect 3 65 7 68
rect 3 63 4 65
rect 6 63 7 65
rect 3 58 7 63
rect 23 65 27 68
rect 23 63 24 65
rect 26 63 27 65
rect 23 61 27 63
rect 3 56 4 58
rect 6 56 7 58
rect 3 54 7 56
rect 3 27 7 29
rect 3 25 4 27
rect 6 25 7 27
rect 3 20 7 25
rect 3 18 4 20
rect 6 18 7 20
rect 3 12 7 18
rect 36 27 42 28
rect 36 25 38 27
rect 40 25 42 27
rect 36 20 42 25
rect 36 18 38 20
rect 40 18 42 20
rect 36 12 42 18
<< labels >>
rlabel alu1 20 24 20 24 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 48 28 48 6 b
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 36 36 36 36 6 a
rlabel alu1 44 40 44 40 6 a
rlabel alu1 36 52 36 52 6 b
<< end >>
