magic
tech scmos
timestamp 1199201675
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 9 66 11 70
rect 19 63 21 68
rect 29 63 31 68
rect 9 35 11 38
rect 19 35 21 46
rect 29 43 31 46
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 29 37 35 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 9 26 11 29
rect 22 26 24 29
rect 29 26 31 37
rect 9 7 11 12
rect 22 7 24 12
rect 29 7 31 12
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 16 9 22
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 12 22 26
rect 24 12 29 26
rect 31 18 36 26
rect 31 16 38 18
rect 31 14 34 16
rect 36 14 38 16
rect 31 12 38 14
rect 13 7 20 12
rect 13 5 15 7
rect 17 5 20 7
rect 13 3 20 5
<< pdif >>
rect 4 59 9 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 4 38 9 46
rect 11 63 17 66
rect 11 61 19 63
rect 11 59 14 61
rect 16 59 19 61
rect 11 46 19 59
rect 21 57 29 63
rect 21 55 24 57
rect 26 55 29 57
rect 21 50 29 55
rect 21 48 24 50
rect 26 48 29 50
rect 21 46 29 48
rect 31 61 38 63
rect 31 59 34 61
rect 36 59 38 61
rect 31 46 38 59
rect 11 38 17 46
<< alu1 >>
rect -2 64 42 72
rect 2 57 7 59
rect 2 55 4 57
rect 6 55 7 57
rect 2 50 7 55
rect 2 48 4 50
rect 6 48 7 50
rect 2 46 7 48
rect 2 24 6 46
rect 34 42 38 51
rect 25 41 38 42
rect 25 39 31 41
rect 33 39 38 41
rect 25 38 38 39
rect 17 33 31 34
rect 17 31 21 33
rect 23 31 31 33
rect 17 30 31 31
rect 2 22 4 24
rect 2 19 6 22
rect 2 16 14 19
rect 2 14 4 16
rect 6 14 14 16
rect 2 13 14 14
rect 26 21 31 30
rect -2 7 42 8
rect -2 5 15 7
rect 17 5 42 7
rect -2 0 42 5
<< nmos >>
rect 9 12 11 26
rect 22 12 24 26
rect 29 12 31 26
<< pmos >>
rect 9 38 11 66
rect 19 46 21 63
rect 29 46 31 63
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 31 39 33 41
rect 21 31 23 33
<< ndifct0 >>
rect 34 14 36 16
<< ndifct1 >>
rect 4 22 6 24
rect 4 14 6 16
rect 15 5 17 7
<< pdifct0 >>
rect 14 59 16 61
rect 24 55 26 57
rect 24 48 26 50
rect 34 59 36 61
<< pdifct1 >>
rect 4 55 6 57
rect 4 48 6 50
<< alu0 >>
rect 13 61 17 64
rect 13 59 14 61
rect 16 59 17 61
rect 33 61 37 64
rect 33 59 34 61
rect 36 59 37 61
rect 13 57 17 59
rect 23 57 27 59
rect 33 57 37 59
rect 23 55 24 57
rect 26 55 27 57
rect 23 50 27 55
rect 10 48 24 50
rect 26 48 27 50
rect 10 46 27 48
rect 10 33 14 46
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 6 19 7 26
rect 10 22 22 26
rect 18 17 22 22
rect 18 16 38 17
rect 18 14 34 16
rect 36 14 38 16
rect 18 13 38 14
<< labels >>
rlabel alu0 12 36 12 36 6 zn
rlabel alu0 28 15 28 15 6 zn
rlabel alu0 25 52 25 52 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 20 32 20 32 6 a
rlabel alu1 28 28 28 28 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 36 48 36 48 6 b
<< end >>
