magic
tech scmos
timestamp 1199202347
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 10 70 12 74
rect 20 61 22 65
rect 10 39 12 42
rect 20 39 22 42
rect 9 37 22 39
rect 9 35 18 37
rect 20 35 22 37
rect 9 33 22 35
rect 9 30 11 33
rect 9 13 11 18
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 18 9 24
rect 11 22 19 30
rect 11 20 14 22
rect 16 20 19 22
rect 11 18 19 20
<< pdif >>
rect 2 68 10 70
rect 2 66 5 68
rect 7 66 10 68
rect 2 61 10 66
rect 2 59 5 61
rect 7 59 10 61
rect 2 42 10 59
rect 12 61 17 70
rect 12 53 20 61
rect 12 51 15 53
rect 17 51 20 53
rect 12 46 20 51
rect 12 44 15 46
rect 17 44 20 46
rect 12 42 20 44
rect 22 59 30 61
rect 22 57 25 59
rect 27 57 30 59
rect 22 52 30 57
rect 22 50 25 52
rect 27 50 30 52
rect 22 42 30 50
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 46 16 47
rect 2 44 15 46
rect 17 44 23 46
rect 2 42 23 44
rect 2 30 6 42
rect 16 37 30 38
rect 16 35 18 37
rect 20 35 30 37
rect 16 34 30 35
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 24 7 26
rect 26 25 30 34
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 18 11 30
<< pmos >>
rect 10 42 12 70
rect 20 42 22 61
<< polyct1 >>
rect 18 35 20 37
<< ndifct0 >>
rect 14 20 16 22
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 5 66 7 68
rect 5 59 7 61
rect 15 51 17 53
rect 25 57 27 59
rect 25 50 27 52
<< pdifct1 >>
rect 15 44 17 46
<< alu0 >>
rect 3 66 5 68
rect 7 66 9 68
rect 3 61 9 66
rect 3 59 5 61
rect 7 59 9 61
rect 3 58 9 59
rect 23 59 29 68
rect 23 57 25 59
rect 27 57 29 59
rect 14 53 18 55
rect 14 51 15 53
rect 17 51 18 53
rect 14 47 18 51
rect 23 52 29 57
rect 23 50 25 52
rect 27 50 29 52
rect 23 49 29 50
rect 16 46 18 47
rect 13 22 17 24
rect 13 20 14 22
rect 16 20 17 22
rect 13 12 17 20
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 20 44 20 44 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 28 28 28 6 a
<< end >>
