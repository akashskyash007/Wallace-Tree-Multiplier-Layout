magic
tech scmos
timestamp 1199203429
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 47 70 49 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 40 31 43
rect 58 56 60 61
rect 68 56 70 61
rect 29 39 39 40
rect 47 39 49 42
rect 58 39 60 42
rect 68 39 70 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 29 38 42 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 36 37 42 38
rect 36 35 38 37
rect 40 35 42 37
rect 13 30 15 33
rect 20 30 22 33
rect 30 30 32 34
rect 36 33 42 35
rect 40 30 42 33
rect 47 37 54 39
rect 58 37 78 39
rect 47 35 50 37
rect 52 35 54 37
rect 47 33 54 35
rect 47 30 49 33
rect 63 30 65 37
rect 72 35 74 37
rect 76 35 78 37
rect 72 33 78 35
rect 13 12 15 17
rect 20 12 22 17
rect 40 12 42 16
rect 47 12 49 16
rect 30 8 32 11
rect 63 8 65 17
rect 30 6 65 8
<< ndif >>
rect 4 17 13 30
rect 15 17 20 30
rect 22 21 30 30
rect 22 19 25 21
rect 27 19 30 21
rect 22 17 30 19
rect 4 11 11 17
rect 25 11 30 17
rect 32 26 40 30
rect 32 24 35 26
rect 37 24 40 26
rect 32 16 40 24
rect 42 16 47 30
rect 49 21 63 30
rect 49 19 58 21
rect 60 19 63 21
rect 49 17 63 19
rect 65 28 72 30
rect 65 26 68 28
rect 70 26 72 28
rect 65 24 72 26
rect 65 17 70 24
rect 49 16 61 17
rect 32 11 37 16
rect 4 9 7 11
rect 9 9 11 11
rect 4 7 11 9
<< pdif >>
rect 72 71 78 73
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 57 9 59
rect 4 42 9 57
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 43 29 51
rect 31 68 38 70
rect 31 66 34 68
rect 36 66 38 68
rect 31 59 38 66
rect 31 43 36 59
rect 42 55 47 70
rect 40 53 47 55
rect 40 51 42 53
rect 44 51 47 53
rect 40 49 47 51
rect 21 42 26 43
rect 42 42 47 49
rect 49 68 56 70
rect 49 66 52 68
rect 54 66 56 68
rect 49 56 56 66
rect 72 69 74 71
rect 76 69 78 71
rect 72 56 78 69
rect 49 42 58 56
rect 60 53 68 56
rect 60 51 63 53
rect 65 51 68 53
rect 60 46 68 51
rect 60 44 63 46
rect 65 44 68 46
rect 60 42 68 44
rect 70 42 78 56
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 71 82 79
rect -2 69 74 71
rect 76 69 82 71
rect -2 68 82 69
rect 64 58 78 63
rect 2 53 17 55
rect 2 51 14 53
rect 16 51 17 53
rect 2 49 17 51
rect 2 22 6 49
rect 34 37 46 39
rect 34 35 38 37
rect 40 35 46 37
rect 34 33 46 35
rect 50 37 54 39
rect 52 35 54 37
rect 2 21 31 22
rect 2 19 25 21
rect 27 19 31 21
rect 2 18 31 19
rect 42 17 46 33
rect 50 30 54 35
rect 74 39 78 58
rect 73 37 78 39
rect 73 35 74 37
rect 76 35 78 37
rect 73 33 78 35
rect 50 26 63 30
rect 50 17 54 26
rect -2 11 82 12
rect -2 9 7 11
rect 9 9 82 11
rect -2 1 82 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 13 17 15 30
rect 20 17 22 30
rect 30 11 32 30
rect 40 16 42 30
rect 47 16 49 30
rect 63 17 65 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 43 31 70
rect 47 42 49 70
rect 58 42 60 56
rect 68 42 70 56
<< polyct0 >>
rect 11 35 13 37
rect 21 35 23 37
<< polyct1 >>
rect 38 35 40 37
rect 50 35 52 37
rect 74 35 76 37
<< ndifct0 >>
rect 35 24 37 26
rect 58 19 60 21
rect 68 26 70 28
<< ndifct1 >>
rect 25 19 27 21
rect 7 9 9 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 59 6 61
rect 24 51 26 53
rect 34 66 36 68
rect 42 51 44 53
rect 52 66 54 68
rect 63 51 65 53
rect 63 44 65 46
<< pdifct1 >>
rect 14 51 16 53
rect 74 69 76 71
<< alu0 >>
rect 32 66 34 68
rect 36 66 38 68
rect 32 65 38 66
rect 50 66 52 68
rect 54 66 56 68
rect 50 65 56 66
rect 2 61 54 62
rect 2 59 4 61
rect 6 59 54 61
rect 2 58 54 59
rect 20 53 46 54
rect 20 51 24 53
rect 26 51 42 53
rect 44 51 46 53
rect 20 50 46 51
rect 20 46 24 50
rect 50 47 54 58
rect 61 53 67 54
rect 61 51 63 53
rect 65 51 67 53
rect 61 47 67 51
rect 10 42 24 46
rect 27 46 70 47
rect 27 44 63 46
rect 65 44 70 46
rect 27 43 70 44
rect 10 37 14 42
rect 27 38 31 43
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 19 37 31 38
rect 19 35 21 37
rect 23 35 31 37
rect 19 34 31 35
rect 49 33 50 39
rect 10 26 38 30
rect 34 24 35 26
rect 37 24 38 26
rect 34 22 38 24
rect 66 30 70 43
rect 66 28 71 30
rect 66 26 68 28
rect 70 26 71 28
rect 66 24 71 26
rect 57 21 61 23
rect 57 19 58 21
rect 60 19 61 21
rect 57 12 61 19
<< labels >>
rlabel polyct0 12 36 12 36 6 an
rlabel alu0 24 28 24 28 6 an
rlabel alu0 25 36 25 36 6 bn
rlabel alu0 33 52 33 52 6 an
rlabel alu0 28 60 28 60 6 bn
rlabel alu0 68 35 68 35 6 bn
rlabel alu0 64 48 64 48 6 bn
rlabel alu0 48 45 48 45 6 bn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 36 36 36 36 6 a2
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 52 28 52 28 6 a1
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 28 60 28 6 a1
rlabel alu1 76 48 76 48 6 b
rlabel alu1 68 60 68 60 6 b
<< end >>
