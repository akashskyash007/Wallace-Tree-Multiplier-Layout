magic
tech scmos
timestamp 1199202497
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 9 62 11 67
rect 19 62 21 67
rect 26 62 28 67
rect 36 62 38 67
rect 43 62 45 67
rect 56 55 62 57
rect 56 53 58 55
rect 60 53 62 55
rect 9 31 11 50
rect 19 41 21 50
rect 16 39 22 41
rect 16 37 18 39
rect 20 37 22 39
rect 16 35 22 37
rect 26 37 28 50
rect 36 47 38 50
rect 33 45 39 47
rect 33 43 35 45
rect 37 43 39 45
rect 33 41 39 43
rect 43 39 45 50
rect 53 51 62 53
rect 53 48 55 51
rect 43 37 49 39
rect 26 35 38 37
rect 8 29 14 31
rect 8 27 10 29
rect 12 27 14 29
rect 8 25 14 27
rect 9 22 11 25
rect 19 22 21 35
rect 26 29 32 31
rect 26 27 28 29
rect 30 27 32 29
rect 26 25 32 27
rect 26 22 28 25
rect 36 22 38 35
rect 43 35 45 37
rect 47 35 49 37
rect 43 33 49 35
rect 43 22 45 33
rect 53 22 55 42
rect 9 11 11 16
rect 19 11 21 16
rect 26 11 28 16
rect 36 8 38 16
rect 43 12 45 16
rect 53 8 55 16
rect 36 6 55 8
<< ndif >>
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 20 19 22
rect 11 18 14 20
rect 16 18 19 20
rect 11 16 19 18
rect 21 16 26 22
rect 28 20 36 22
rect 28 18 31 20
rect 33 18 36 20
rect 28 16 36 18
rect 38 16 43 22
rect 45 20 53 22
rect 45 18 48 20
rect 50 18 53 20
rect 45 16 53 18
rect 55 20 62 22
rect 55 18 58 20
rect 60 18 62 20
rect 55 16 62 18
<< pdif >>
rect 4 56 9 62
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 11 60 19 62
rect 11 58 14 60
rect 16 58 19 60
rect 11 50 19 58
rect 21 50 26 62
rect 28 54 36 62
rect 28 52 31 54
rect 33 52 36 54
rect 28 50 36 52
rect 38 50 43 62
rect 45 60 52 62
rect 45 58 48 60
rect 50 58 52 60
rect 45 56 52 58
rect 45 50 51 56
rect 47 48 51 50
rect 47 42 53 48
rect 55 46 62 48
rect 55 44 58 46
rect 60 44 62 46
rect 55 42 62 44
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 57 55 62 63
rect 2 54 8 55
rect 57 54 58 55
rect 2 52 4 54
rect 6 52 15 54
rect 2 50 15 52
rect 49 53 58 54
rect 60 53 62 55
rect 49 50 62 53
rect 2 21 6 50
rect 25 40 31 46
rect 16 39 31 40
rect 16 37 18 39
rect 20 37 31 39
rect 16 34 31 37
rect 42 37 48 39
rect 42 35 45 37
rect 47 35 48 37
rect 42 31 48 35
rect 42 25 54 31
rect 2 20 8 21
rect 2 18 4 20
rect 6 18 8 20
rect 2 17 8 18
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 16 11 22
rect 19 16 21 22
rect 26 16 28 22
rect 36 16 38 22
rect 43 16 45 22
rect 53 16 55 22
<< pmos >>
rect 9 50 11 62
rect 19 50 21 62
rect 26 50 28 62
rect 36 50 38 62
rect 43 50 45 62
rect 53 42 55 48
<< polyct0 >>
rect 35 43 37 45
rect 10 27 12 29
rect 28 27 30 29
<< polyct1 >>
rect 58 53 60 55
rect 18 37 20 39
rect 45 35 47 37
<< ndifct0 >>
rect 14 18 16 20
rect 31 18 33 20
rect 48 18 50 20
rect 58 18 60 20
<< ndifct1 >>
rect 4 18 6 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 14 58 16 60
rect 31 52 33 54
rect 48 58 50 60
rect 58 44 60 46
<< pdifct1 >>
rect 4 52 6 54
<< alu0 >>
rect 12 60 18 68
rect 12 58 14 60
rect 16 58 18 60
rect 12 57 18 58
rect 46 60 52 68
rect 46 58 48 60
rect 50 58 52 60
rect 46 57 52 58
rect 29 54 35 55
rect 18 52 31 54
rect 33 52 35 54
rect 18 50 35 52
rect 18 47 22 50
rect 9 43 22 47
rect 34 46 62 47
rect 9 29 13 43
rect 34 45 58 46
rect 34 43 35 45
rect 37 44 58 45
rect 60 44 62 46
rect 37 43 62 44
rect 34 31 38 43
rect 27 29 38 31
rect 9 27 10 29
rect 12 27 24 29
rect 9 25 24 27
rect 27 27 28 29
rect 30 27 38 29
rect 27 25 38 27
rect 13 20 17 22
rect 13 18 14 20
rect 16 18 17 20
rect 13 12 17 18
rect 20 21 24 25
rect 58 21 62 43
rect 20 20 35 21
rect 20 18 31 20
rect 33 18 35 20
rect 20 17 35 18
rect 46 20 52 21
rect 46 18 48 20
rect 50 18 52 20
rect 46 12 52 18
rect 56 20 62 21
rect 56 18 58 20
rect 60 18 62 20
rect 56 17 62 18
<< labels >>
rlabel alu0 11 36 11 36 6 zn
rlabel alu0 27 19 27 19 6 zn
rlabel alu0 32 28 32 28 6 sn
rlabel alu0 36 36 36 36 6 sn
rlabel alu0 26 52 26 52 6 zn
rlabel alu0 60 32 60 32 6 sn
rlabel alu0 48 45 48 45 6 sn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 36 20 36 6 a0
rlabel alu1 28 40 28 40 6 a0
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 a1
rlabel alu1 52 52 52 52 6 s
rlabel alu1 60 60 60 60 6 s
<< end >>
