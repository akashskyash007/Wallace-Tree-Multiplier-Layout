magic
tech scmos
timestamp 1199203033
<< ab >>
rect 0 0 136 80
<< nwell >>
rect -5 36 141 88
<< pwell >>
rect -5 -8 141 36
<< poly >>
rect 39 70 41 74
rect 46 70 48 74
rect 53 70 55 74
rect 63 70 65 74
rect 70 70 72 74
rect 77 70 79 74
rect 87 70 89 74
rect 94 70 96 74
rect 101 70 103 74
rect 111 70 113 74
rect 118 70 120 74
rect 125 70 127 74
rect 15 62 17 67
rect 22 62 24 67
rect 29 62 31 67
rect 15 39 17 42
rect 9 37 17 39
rect 9 35 11 37
rect 13 35 17 37
rect 9 33 17 35
rect 9 22 11 33
rect 22 31 24 42
rect 29 39 31 42
rect 39 39 41 42
rect 29 37 41 39
rect 35 35 37 37
rect 39 35 41 37
rect 46 39 48 42
rect 53 39 55 42
rect 63 39 65 42
rect 46 36 49 39
rect 53 37 65 39
rect 35 33 41 35
rect 21 29 27 31
rect 21 28 23 29
rect 19 27 23 28
rect 25 27 27 29
rect 39 27 41 33
rect 47 31 49 36
rect 47 29 55 31
rect 47 27 50 29
rect 52 27 55 29
rect 19 25 27 27
rect 31 25 43 27
rect 47 25 55 27
rect 19 22 21 25
rect 31 22 33 25
rect 41 22 43 25
rect 53 22 55 25
rect 63 24 65 37
rect 70 31 72 42
rect 77 39 79 42
rect 87 39 89 42
rect 77 37 90 39
rect 84 35 86 37
rect 88 35 90 37
rect 84 33 90 35
rect 70 29 80 31
rect 74 27 76 29
rect 78 27 80 29
rect 74 25 80 27
rect 9 6 11 10
rect 19 6 21 10
rect 31 6 33 10
rect 41 6 43 10
rect 94 23 96 42
rect 90 21 96 23
rect 90 19 92 21
rect 94 19 96 21
rect 90 17 96 19
rect 101 39 103 42
rect 111 39 113 42
rect 101 37 113 39
rect 101 35 107 37
rect 109 35 113 37
rect 101 33 113 35
rect 53 6 55 10
rect 63 9 65 12
rect 101 9 103 33
rect 118 23 120 42
rect 125 31 127 42
rect 125 29 131 31
rect 125 27 127 29
rect 129 27 131 29
rect 125 25 131 27
rect 113 21 120 23
rect 113 19 115 21
rect 117 19 120 21
rect 113 17 120 19
rect 63 7 103 9
<< ndif >>
rect 58 22 63 24
rect 2 14 9 22
rect 2 12 4 14
rect 6 12 9 14
rect 2 10 9 12
rect 11 20 19 22
rect 11 18 14 20
rect 16 18 19 20
rect 11 10 19 18
rect 21 11 31 22
rect 21 10 25 11
rect 23 9 25 10
rect 27 10 31 11
rect 33 20 41 22
rect 33 18 36 20
rect 38 18 41 20
rect 33 10 41 18
rect 43 11 53 22
rect 43 10 47 11
rect 27 9 29 10
rect 23 7 29 9
rect 45 9 47 10
rect 49 10 53 11
rect 55 20 63 22
rect 55 18 58 20
rect 60 18 63 20
rect 55 12 63 18
rect 65 16 72 24
rect 65 14 68 16
rect 70 14 72 16
rect 65 12 72 14
rect 55 10 60 12
rect 49 9 51 10
rect 45 7 51 9
<< pdif >>
rect 33 62 39 70
rect 8 60 15 62
rect 8 58 10 60
rect 12 58 15 60
rect 8 53 15 58
rect 8 51 10 53
rect 12 51 15 53
rect 8 49 15 51
rect 10 42 15 49
rect 17 42 22 62
rect 24 42 29 62
rect 31 60 39 62
rect 31 58 34 60
rect 36 58 39 60
rect 31 42 39 58
rect 41 42 46 70
rect 48 42 53 70
rect 55 61 63 70
rect 55 59 58 61
rect 60 59 63 61
rect 55 53 63 59
rect 55 51 58 53
rect 60 51 63 53
rect 55 42 63 51
rect 65 42 70 70
rect 72 42 77 70
rect 79 68 87 70
rect 79 66 82 68
rect 84 66 87 68
rect 79 61 87 66
rect 79 59 82 61
rect 84 59 87 61
rect 79 42 87 59
rect 89 42 94 70
rect 96 42 101 70
rect 103 61 111 70
rect 103 59 106 61
rect 108 59 111 61
rect 103 53 111 59
rect 103 51 106 53
rect 108 51 111 53
rect 103 42 111 51
rect 113 42 118 70
rect 120 42 125 70
rect 127 68 134 70
rect 127 66 130 68
rect 132 66 134 68
rect 127 61 134 66
rect 127 59 130 61
rect 132 59 134 61
rect 127 42 134 59
<< alu1 >>
rect -2 81 138 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 138 81
rect -2 68 138 79
rect 9 60 14 63
rect 9 58 10 60
rect 12 58 14 60
rect 9 55 14 58
rect 57 61 62 63
rect 57 59 58 61
rect 60 59 62 61
rect 2 54 14 55
rect 57 54 62 59
rect 105 61 111 63
rect 105 59 106 61
rect 108 59 111 61
rect 105 54 111 59
rect 2 53 111 54
rect 2 51 10 53
rect 12 51 58 53
rect 60 51 106 53
rect 108 51 111 53
rect 2 50 111 51
rect 2 29 6 50
rect 10 42 111 46
rect 10 37 14 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 25 30 31 38
rect 35 37 98 38
rect 35 35 37 37
rect 39 35 86 37
rect 88 35 98 37
rect 35 34 98 35
rect 105 37 111 42
rect 105 35 107 37
rect 109 35 111 37
rect 105 34 111 35
rect 94 30 98 34
rect 21 29 87 30
rect 2 25 14 29
rect 21 27 23 29
rect 25 27 50 29
rect 52 27 76 29
rect 78 27 87 29
rect 21 26 87 27
rect 94 29 131 30
rect 94 27 127 29
rect 129 27 131 29
rect 94 26 131 27
rect 10 22 14 25
rect 81 22 87 26
rect 10 20 63 22
rect 10 18 14 20
rect 16 18 36 20
rect 38 18 58 20
rect 60 18 63 20
rect 81 21 119 22
rect 81 19 92 21
rect 94 19 115 21
rect 117 19 119 21
rect 81 18 119 19
rect 10 17 63 18
rect -2 11 138 12
rect -2 9 25 11
rect 27 9 47 11
rect 49 9 138 11
rect -2 1 138 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 138 1
rect -2 -2 138 -1
<< ptie >>
rect 0 1 136 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 136 1
rect 0 -3 136 -1
<< ntie >>
rect 0 81 136 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 136 81
rect 0 77 136 79
<< nmos >>
rect 9 10 11 22
rect 19 10 21 22
rect 31 10 33 22
rect 41 10 43 22
rect 53 10 55 22
rect 63 12 65 24
<< pmos >>
rect 15 42 17 62
rect 22 42 24 62
rect 29 42 31 62
rect 39 42 41 70
rect 46 42 48 70
rect 53 42 55 70
rect 63 42 65 70
rect 70 42 72 70
rect 77 42 79 70
rect 87 42 89 70
rect 94 42 96 70
rect 101 42 103 70
rect 111 42 113 70
rect 118 42 120 70
rect 125 42 127 70
<< polyct1 >>
rect 11 35 13 37
rect 37 35 39 37
rect 23 27 25 29
rect 50 27 52 29
rect 86 35 88 37
rect 76 27 78 29
rect 92 19 94 21
rect 107 35 109 37
rect 127 27 129 29
rect 115 19 117 21
<< ndifct0 >>
rect 4 12 6 14
rect 68 14 70 16
<< ndifct1 >>
rect 14 18 16 20
rect 25 9 27 11
rect 36 18 38 20
rect 47 9 49 11
rect 58 18 60 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
<< pdifct0 >>
rect 34 58 36 60
rect 82 66 84 68
rect 82 59 84 61
rect 130 66 132 68
rect 130 59 132 61
<< pdifct1 >>
rect 10 58 12 60
rect 10 51 12 53
rect 58 59 60 61
rect 58 51 60 53
rect 106 59 108 61
rect 106 51 108 53
<< alu0 >>
rect 32 60 38 68
rect 80 66 82 68
rect 84 66 86 68
rect 32 58 34 60
rect 36 58 38 60
rect 32 57 38 58
rect 80 61 86 66
rect 128 66 130 68
rect 132 66 134 68
rect 80 59 82 61
rect 84 59 86 61
rect 80 58 86 59
rect 128 61 134 66
rect 128 59 130 61
rect 132 59 134 61
rect 128 58 134 59
rect 67 16 71 18
rect 3 14 7 16
rect 3 12 4 14
rect 6 12 7 14
rect 67 14 68 16
rect 70 14 71 16
rect 67 12 71 14
<< labels >>
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 44 20 44 6 c
rlabel alu1 4 40 4 40 6 z
rlabel polyct1 12 36 12 36 6 c
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 44 28 44 28 6 b
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 28 36 28 6 b
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 32 28 32 6 b
rlabel alu1 28 44 28 44 6 c
rlabel alu1 44 44 44 44 6 c
rlabel alu1 44 36 44 36 6 a
rlabel alu1 36 44 36 44 6 c
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 68 6 68 6 6 vss
rlabel alu1 52 20 52 20 6 z
rlabel alu1 52 28 52 28 6 b
rlabel alu1 68 28 68 28 6 b
rlabel alu1 76 28 76 28 6 b
rlabel alu1 60 28 60 28 6 b
rlabel alu1 60 20 60 20 6 z
rlabel alu1 52 36 52 36 6 a
rlabel alu1 52 44 52 44 6 c
rlabel alu1 68 44 68 44 6 c
rlabel alu1 76 44 76 44 6 c
rlabel alu1 76 36 76 36 6 a
rlabel alu1 68 36 68 36 6 a
rlabel alu1 60 44 60 44 6 c
rlabel alu1 60 36 60 36 6 a
rlabel alu1 68 52 68 52 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 60 56 60 56 6 z
rlabel alu1 68 74 68 74 6 vdd
rlabel alu1 84 20 84 20 6 b
rlabel alu1 84 28 84 28 6 b
rlabel alu1 108 28 108 28 6 a
rlabel alu1 100 28 100 28 6 a
rlabel alu1 100 20 100 20 6 b
rlabel alu1 108 20 108 20 6 b
rlabel alu1 92 20 92 20 6 b
rlabel alu1 84 36 84 36 6 a
rlabel alu1 84 44 84 44 6 c
rlabel alu1 92 44 92 44 6 c
rlabel alu1 108 40 108 40 6 c
rlabel alu1 100 44 100 44 6 c
rlabel alu1 92 36 92 36 6 a
rlabel alu1 92 52 92 52 6 z
rlabel alu1 100 52 100 52 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 108 56 108 56 6 z
rlabel alu1 116 28 116 28 6 a
rlabel alu1 124 28 124 28 6 a
rlabel polyct1 116 20 116 20 6 b
<< end >>
