magic
tech scmos
timestamp 1199470207
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 15 94 17 98
rect 27 94 29 98
rect 35 94 37 98
rect 47 94 49 98
rect 55 94 57 98
rect 15 53 17 56
rect 15 51 23 53
rect 15 49 19 51
rect 21 49 23 51
rect 15 47 23 49
rect 27 47 29 56
rect 35 53 37 56
rect 47 53 49 56
rect 35 51 49 53
rect 55 53 57 56
rect 55 51 63 53
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 55 49 59 51
rect 61 49 63 51
rect 55 47 63 49
rect 15 38 17 47
rect 27 45 33 47
rect 27 43 29 45
rect 31 43 33 45
rect 27 41 33 43
rect 39 43 43 47
rect 39 41 53 43
rect 27 38 29 41
rect 39 38 41 41
rect 51 38 53 41
rect 39 17 41 22
rect 51 17 53 22
rect 15 2 17 6
rect 27 2 29 6
<< ndif >>
rect 7 36 15 38
rect 7 34 9 36
rect 11 34 15 36
rect 7 28 15 34
rect 7 26 9 28
rect 11 26 15 28
rect 7 24 15 26
rect 10 6 15 24
rect 17 31 27 38
rect 17 29 21 31
rect 23 29 27 31
rect 17 21 27 29
rect 17 19 21 21
rect 23 19 27 21
rect 17 6 27 19
rect 29 22 39 38
rect 41 31 51 38
rect 41 29 45 31
rect 47 29 51 31
rect 41 22 51 29
rect 53 31 62 38
rect 53 29 57 31
rect 59 29 62 31
rect 53 22 62 29
rect 29 21 37 22
rect 29 19 33 21
rect 35 19 37 21
rect 29 11 37 19
rect 29 9 33 11
rect 35 9 37 11
rect 29 6 37 9
<< pdif >>
rect 10 70 15 94
rect 7 68 15 70
rect 7 66 9 68
rect 11 66 15 68
rect 7 60 15 66
rect 7 58 9 60
rect 11 58 15 60
rect 7 56 15 58
rect 17 91 27 94
rect 17 89 21 91
rect 23 89 27 91
rect 17 81 27 89
rect 17 79 21 81
rect 23 79 27 81
rect 17 56 27 79
rect 29 56 35 94
rect 37 81 47 94
rect 37 79 41 81
rect 43 79 47 81
rect 37 71 47 79
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 49 56 55 94
rect 57 91 66 94
rect 57 89 61 91
rect 63 89 66 91
rect 57 81 66 89
rect 57 79 61 81
rect 63 79 66 81
rect 57 56 66 79
<< alu1 >>
rect -2 91 72 100
rect -2 89 21 91
rect 23 89 61 91
rect 63 89 72 91
rect -2 88 72 89
rect 20 81 24 88
rect 20 79 21 81
rect 23 79 24 81
rect 20 77 24 79
rect 38 81 44 83
rect 38 79 41 81
rect 43 79 44 81
rect 38 73 44 79
rect 60 81 64 88
rect 60 79 61 81
rect 63 79 64 81
rect 60 77 64 79
rect 8 71 44 73
rect 8 69 41 71
rect 43 69 44 71
rect 8 68 44 69
rect 8 66 9 68
rect 11 67 44 68
rect 11 66 12 67
rect 8 60 12 66
rect 48 63 52 73
rect 8 58 9 60
rect 11 58 12 60
rect 8 36 12 58
rect 18 58 33 63
rect 18 51 22 58
rect 18 49 19 51
rect 21 49 22 51
rect 18 37 22 49
rect 38 57 52 63
rect 38 51 42 57
rect 38 49 39 51
rect 41 49 42 51
rect 38 47 42 49
rect 58 51 63 63
rect 58 49 59 51
rect 61 49 63 51
rect 27 45 33 47
rect 27 43 29 45
rect 31 43 33 45
rect 27 42 33 43
rect 58 42 63 49
rect 27 38 63 42
rect 8 34 9 36
rect 11 34 12 36
rect 8 28 12 34
rect 8 26 9 28
rect 11 26 12 28
rect 8 24 12 26
rect 19 31 49 32
rect 19 29 21 31
rect 23 29 45 31
rect 47 29 49 31
rect 19 28 49 29
rect 56 31 60 33
rect 56 29 57 31
rect 59 29 60 31
rect 19 21 25 28
rect 19 19 21 21
rect 23 19 25 21
rect 19 18 25 19
rect 32 21 36 23
rect 32 19 33 21
rect 35 19 36 21
rect 32 12 36 19
rect 56 12 60 29
rect -2 11 72 12
rect -2 9 33 11
rect 35 9 72 11
rect -2 7 72 9
rect -2 5 49 7
rect 51 5 59 7
rect 61 5 72 7
rect -2 0 72 5
<< ptie >>
rect 47 7 63 9
rect 47 5 49 7
rect 51 5 59 7
rect 61 5 63 7
rect 47 3 63 5
<< nmos >>
rect 15 6 17 38
rect 27 6 29 38
rect 39 22 41 38
rect 51 22 53 38
<< pmos >>
rect 15 56 17 94
rect 27 56 29 94
rect 35 56 37 94
rect 47 56 49 94
rect 55 56 57 94
<< polyct1 >>
rect 19 49 21 51
rect 39 49 41 51
rect 59 49 61 51
rect 29 43 31 45
<< ndifct1 >>
rect 9 34 11 36
rect 9 26 11 28
rect 21 29 23 31
rect 21 19 23 21
rect 45 29 47 31
rect 57 29 59 31
rect 33 19 35 21
rect 33 9 35 11
<< ptiect1 >>
rect 49 5 51 7
rect 59 5 61 7
<< pdifct1 >>
rect 9 66 11 68
rect 9 58 11 60
rect 21 89 23 91
rect 21 79 23 81
rect 41 79 43 81
rect 41 69 43 71
rect 61 89 63 91
rect 61 79 63 81
<< labels >>
rlabel alu1 22 25 22 25 6 n3
rlabel alu1 10 50 10 50 6 z
rlabel polyct1 20 50 20 50 6 b
rlabel alu1 20 70 20 70 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 30 40 30 40 6 a1
rlabel alu1 30 60 30 60 6 b
rlabel alu1 30 70 30 70 6 z
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 34 30 34 30 6 n3
rlabel alu1 50 40 50 40 6 a1
rlabel alu1 40 40 40 40 6 a1
rlabel alu1 40 55 40 55 6 a2
rlabel alu1 40 75 40 75 6 z
rlabel alu1 50 65 50 65 6 a2
rlabel polyct1 60 50 60 50 6 a1
<< end >>
