magic
tech scmos
timestamp 1199542766
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 11 94 13 98
rect 19 94 21 98
rect 27 94 29 98
rect 43 94 45 98
rect 55 94 57 98
rect 11 33 13 56
rect 19 43 21 56
rect 27 53 29 56
rect 67 76 69 80
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 37 49
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 7 31 13 33
rect 7 29 9 31
rect 11 29 13 31
rect 7 27 13 29
rect 19 29 21 37
rect 19 27 25 29
rect 11 24 13 27
rect 23 24 25 27
rect 35 25 37 47
rect 43 43 45 55
rect 55 43 57 55
rect 67 53 69 56
rect 61 51 69 53
rect 61 49 63 51
rect 65 49 69 51
rect 61 47 69 49
rect 43 41 63 43
rect 43 39 59 41
rect 61 39 63 41
rect 43 37 63 39
rect 45 25 47 37
rect 57 25 59 37
rect 67 25 69 47
rect 11 10 13 14
rect 23 10 25 14
rect 35 11 37 15
rect 67 11 69 15
rect 45 2 47 6
rect 57 2 59 6
<< ndif >>
rect 30 24 35 25
rect 3 21 11 24
rect 3 19 5 21
rect 7 19 11 21
rect 3 14 11 19
rect 13 14 23 24
rect 25 21 35 24
rect 25 19 29 21
rect 31 19 35 21
rect 25 15 35 19
rect 37 15 45 25
rect 25 14 33 15
rect 15 11 21 14
rect 15 9 17 11
rect 19 9 21 11
rect 39 9 45 15
rect 15 7 21 9
rect 37 7 45 9
rect 37 5 39 7
rect 41 6 45 7
rect 47 21 57 25
rect 47 19 51 21
rect 53 19 57 21
rect 47 6 57 19
rect 59 15 67 25
rect 69 21 77 25
rect 69 19 73 21
rect 75 19 77 21
rect 69 15 77 19
rect 59 9 65 15
rect 59 7 67 9
rect 59 6 63 7
rect 41 5 43 6
rect 37 3 43 5
rect 61 5 63 6
rect 65 5 67 7
rect 61 3 67 5
<< pdif >>
rect 3 81 11 94
rect 3 79 5 81
rect 7 79 11 81
rect 3 56 11 79
rect 13 56 19 94
rect 21 56 27 94
rect 29 91 43 94
rect 29 89 37 91
rect 39 89 43 91
rect 29 56 43 89
rect 35 55 43 56
rect 45 71 55 94
rect 45 69 49 71
rect 51 69 55 71
rect 45 61 55 69
rect 45 59 49 61
rect 51 59 55 61
rect 45 55 55 59
rect 57 91 65 94
rect 57 89 61 91
rect 63 89 65 91
rect 57 76 65 89
rect 57 56 67 76
rect 69 61 77 76
rect 69 59 73 61
rect 75 59 77 61
rect 69 56 77 59
rect 57 55 62 56
<< alu1 >>
rect -2 95 82 100
rect -2 93 73 95
rect 75 93 82 95
rect -2 91 82 93
rect -2 89 37 91
rect 39 89 61 91
rect 63 89 82 91
rect -2 88 82 89
rect 3 81 66 82
rect 3 79 5 81
rect 7 79 66 81
rect 3 78 66 79
rect 8 31 12 73
rect 8 29 9 31
rect 11 29 12 31
rect 8 27 12 29
rect 18 41 22 73
rect 18 39 19 41
rect 21 39 22 41
rect 18 27 22 39
rect 28 51 32 73
rect 28 49 29 51
rect 31 49 32 51
rect 28 27 32 49
rect 38 22 42 78
rect 3 21 42 22
rect 3 19 5 21
rect 7 19 29 21
rect 31 19 42 21
rect 3 18 42 19
rect 48 71 52 73
rect 48 69 49 71
rect 51 69 52 71
rect 48 61 52 69
rect 48 59 49 61
rect 51 59 52 61
rect 48 22 52 59
rect 62 51 66 78
rect 62 49 63 51
rect 65 49 66 51
rect 62 47 66 49
rect 72 61 76 63
rect 72 59 73 61
rect 75 59 76 61
rect 72 42 76 59
rect 57 41 76 42
rect 57 39 59 41
rect 61 39 76 41
rect 57 38 76 39
rect 48 21 55 22
rect 48 19 51 21
rect 53 19 55 21
rect 48 18 55 19
rect 72 21 76 38
rect 72 19 73 21
rect 75 19 76 21
rect 48 17 52 18
rect 72 17 76 19
rect -2 11 82 12
rect -2 9 17 11
rect 19 9 82 11
rect -2 7 82 9
rect -2 5 39 7
rect 41 5 63 7
rect 65 5 82 7
rect -2 0 82 5
<< ntie >>
rect 71 95 77 97
rect 71 93 73 95
rect 75 93 77 95
rect 71 86 77 93
<< nmos >>
rect 11 14 13 24
rect 23 14 25 24
rect 35 15 37 25
rect 45 6 47 25
rect 57 6 59 25
rect 67 15 69 25
<< pmos >>
rect 11 56 13 94
rect 19 56 21 94
rect 27 56 29 94
rect 43 55 45 94
rect 55 55 57 94
rect 67 56 69 76
<< polyct1 >>
rect 29 49 31 51
rect 19 39 21 41
rect 9 29 11 31
rect 63 49 65 51
rect 59 39 61 41
<< ndifct1 >>
rect 5 19 7 21
rect 29 19 31 21
rect 17 9 19 11
rect 39 5 41 7
rect 51 19 53 21
rect 73 19 75 21
rect 63 5 65 7
<< ntiect1 >>
rect 73 93 75 95
<< pdifct1 >>
rect 5 79 7 81
rect 37 89 39 91
rect 49 69 51 71
rect 49 59 51 61
rect 61 89 63 91
rect 73 59 75 61
<< labels >>
rlabel alu1 10 50 10 50 6 i2
rlabel polyct1 30 50 30 50 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel ndifct1 40 6 40 6 6 vss
rlabel alu1 50 45 50 45 6 nq
rlabel alu1 40 94 40 94 6 vdd
<< end >>
