magic
tech scmos
timestamp 1199202466
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 20 72 55 74
rect 10 54 12 59
rect 20 54 22 72
rect 53 63 55 72
rect 30 61 36 63
rect 30 59 32 61
rect 34 59 36 61
rect 30 57 36 59
rect 30 54 32 57
rect 40 54 42 59
rect 53 46 55 57
rect 50 44 56 46
rect 50 42 52 44
rect 54 42 56 44
rect 10 39 12 42
rect 2 37 12 39
rect 20 38 22 42
rect 2 35 4 37
rect 6 35 12 37
rect 2 33 12 35
rect 30 34 32 42
rect 10 23 12 33
rect 20 32 32 34
rect 40 39 42 42
rect 50 40 56 42
rect 40 37 46 39
rect 40 35 42 37
rect 44 35 46 37
rect 40 33 46 35
rect 20 23 22 32
rect 30 23 32 28
rect 40 23 42 33
rect 53 27 55 40
rect 53 18 55 21
rect 10 12 12 17
rect 20 12 22 17
rect 30 9 32 17
rect 40 13 42 17
rect 51 15 55 18
rect 51 9 53 15
rect 30 7 53 9
<< ndif >>
rect 44 23 53 27
rect 2 21 10 23
rect 2 19 4 21
rect 6 19 10 21
rect 2 17 10 19
rect 12 21 20 23
rect 12 19 15 21
rect 17 19 20 21
rect 12 17 20 19
rect 22 21 30 23
rect 22 19 25 21
rect 27 19 30 21
rect 22 17 30 19
rect 32 21 40 23
rect 32 19 35 21
rect 37 19 40 21
rect 32 17 40 19
rect 42 21 53 23
rect 55 25 62 27
rect 55 23 58 25
rect 60 23 62 25
rect 55 21 62 23
rect 42 19 45 21
rect 47 19 49 21
rect 42 17 49 19
<< pdif >>
rect 2 62 8 64
rect 2 60 4 62
rect 6 60 8 62
rect 2 54 8 60
rect 44 68 50 70
rect 44 66 46 68
rect 48 66 50 68
rect 44 63 50 66
rect 44 57 53 63
rect 55 61 62 63
rect 55 59 58 61
rect 60 59 62 61
rect 55 57 62 59
rect 44 54 50 57
rect 2 42 10 54
rect 12 46 20 54
rect 12 44 15 46
rect 17 44 20 46
rect 12 42 20 44
rect 22 46 30 54
rect 22 44 25 46
rect 27 44 30 46
rect 22 42 30 44
rect 32 46 40 54
rect 32 44 35 46
rect 37 44 40 46
rect 32 42 40 44
rect 42 49 50 54
rect 42 42 48 49
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 50 15 54
rect 2 39 6 50
rect 26 48 30 55
rect 41 50 54 54
rect 2 37 7 39
rect 2 35 4 37
rect 6 35 7 37
rect 2 33 7 35
rect 24 46 30 48
rect 24 44 25 46
rect 27 44 30 46
rect 24 42 30 44
rect 26 23 30 42
rect 24 21 30 23
rect 24 19 25 21
rect 27 19 30 21
rect 24 17 30 19
rect 50 46 54 50
rect 50 44 55 46
rect 50 42 52 44
rect 54 42 55 44
rect 50 40 55 42
rect 41 37 46 39
rect 41 35 42 37
rect 44 35 46 37
rect 41 33 46 35
rect 42 31 46 33
rect 42 25 54 31
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 10 17 12 23
rect 20 17 22 23
rect 30 17 32 23
rect 40 17 42 23
rect 53 21 55 27
<< pmos >>
rect 53 57 55 63
rect 10 42 12 54
rect 20 42 22 54
rect 30 42 32 54
rect 40 42 42 54
<< polyct0 >>
rect 32 59 34 61
<< polyct1 >>
rect 52 42 54 44
rect 4 35 6 37
rect 42 35 44 37
<< ndifct0 >>
rect 4 19 6 21
rect 15 19 17 21
rect 35 19 37 21
rect 58 23 60 25
rect 45 19 47 21
<< ndifct1 >>
rect 25 19 27 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 4 60 6 62
rect 46 66 48 68
rect 58 59 60 61
rect 15 44 17 46
rect 35 44 37 46
<< pdifct1 >>
rect 25 44 27 46
<< alu0 >>
rect 3 62 7 68
rect 44 66 46 68
rect 48 66 50 68
rect 44 65 50 66
rect 3 60 4 62
rect 6 60 7 62
rect 3 58 7 60
rect 30 61 62 62
rect 30 59 32 61
rect 34 59 58 61
rect 60 59 62 61
rect 30 58 62 59
rect 13 46 20 47
rect 13 44 15 46
rect 17 44 20 46
rect 13 43 20 44
rect 3 21 7 23
rect 16 22 20 43
rect 3 19 4 21
rect 6 19 7 21
rect 3 12 7 19
rect 13 21 20 22
rect 13 19 15 21
rect 17 19 20 21
rect 13 18 20 19
rect 33 46 39 47
rect 33 44 35 46
rect 37 44 39 46
rect 33 43 39 44
rect 33 22 37 43
rect 58 27 62 58
rect 57 25 62 27
rect 57 23 58 25
rect 60 23 62 25
rect 33 21 39 22
rect 33 19 35 21
rect 37 19 39 21
rect 33 18 39 19
rect 43 21 49 22
rect 57 21 62 23
rect 43 19 45 21
rect 47 19 49 21
rect 43 12 49 19
<< labels >>
rlabel alu0 18 32 18 32 6 a0n
rlabel pdifct0 16 45 16 45 6 a0n
rlabel alu0 35 32 35 32 6 a1n
rlabel pdifct0 36 45 36 45 6 a1n
rlabel alu0 46 60 46 60 6 sn
rlabel alu0 60 41 60 41 6 sn
rlabel alu1 4 40 4 40 6 a0
rlabel alu1 12 52 12 52 6 a0
rlabel alu1 28 36 28 36 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 44 52 44 52 6 s
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 a1
rlabel alu1 52 44 52 44 6 s
<< end >>
