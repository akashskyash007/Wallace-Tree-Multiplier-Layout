magic
tech scmos
timestamp 1199203549
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 19 70 21 74
rect 29 70 31 74
rect 36 70 38 74
rect 9 63 11 68
rect 69 58 71 63
rect 52 52 58 54
rect 52 50 54 52
rect 56 50 58 52
rect 9 44 11 47
rect 9 42 15 44
rect 9 40 11 42
rect 13 40 15 42
rect 9 38 15 40
rect 19 39 21 47
rect 10 23 12 38
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 29 38 31 47
rect 36 44 38 47
rect 52 44 58 50
rect 36 42 58 44
rect 29 36 48 38
rect 19 33 25 35
rect 37 34 44 36
rect 46 34 48 36
rect 19 29 21 33
rect 17 26 21 29
rect 37 32 48 34
rect 56 35 58 42
rect 69 39 71 42
rect 65 37 71 39
rect 65 35 67 37
rect 69 35 71 37
rect 56 32 59 35
rect 65 33 71 35
rect 17 23 19 26
rect 27 23 29 28
rect 37 23 39 32
rect 57 29 59 32
rect 69 24 71 33
rect 57 18 59 22
rect 10 11 12 16
rect 17 11 19 16
rect 27 8 29 16
rect 37 12 39 16
rect 69 8 71 17
rect 27 6 71 8
<< ndif >>
rect 50 26 57 29
rect 50 24 52 26
rect 54 24 57 26
rect 2 16 10 23
rect 12 16 17 23
rect 19 21 27 23
rect 19 19 22 21
rect 24 19 27 21
rect 19 16 27 19
rect 29 21 37 23
rect 29 19 32 21
rect 34 19 37 21
rect 29 16 37 19
rect 39 20 46 23
rect 50 22 57 24
rect 59 24 67 29
rect 59 22 69 24
rect 39 18 42 20
rect 44 18 46 20
rect 61 21 69 22
rect 61 19 63 21
rect 65 19 69 21
rect 39 16 46 18
rect 61 17 69 19
rect 71 22 78 24
rect 71 20 74 22
rect 76 20 78 22
rect 71 17 78 20
rect 2 11 8 16
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
<< pdif >>
rect 61 71 67 73
rect 14 63 19 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 57 9 59
rect 4 47 9 57
rect 11 53 19 63
rect 11 51 14 53
rect 16 51 19 53
rect 11 47 19 51
rect 21 51 29 70
rect 21 49 24 51
rect 26 49 29 51
rect 21 47 29 49
rect 31 47 36 70
rect 38 68 47 70
rect 38 66 41 68
rect 43 66 47 68
rect 38 47 47 66
rect 61 69 63 71
rect 65 69 67 71
rect 61 58 67 69
rect 61 42 69 58
rect 71 55 76 58
rect 71 53 78 55
rect 71 51 74 53
rect 76 51 78 53
rect 71 46 78 51
rect 71 44 74 46
rect 76 44 78 46
rect 71 42 78 44
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 71 82 79
rect -2 69 63 71
rect 65 69 82 71
rect -2 68 82 69
rect 2 53 18 54
rect 2 51 14 53
rect 16 51 18 53
rect 2 50 18 51
rect 2 22 6 50
rect 42 39 46 55
rect 50 52 62 55
rect 50 50 54 52
rect 56 50 62 52
rect 50 49 62 50
rect 58 41 62 49
rect 42 36 54 39
rect 42 34 44 36
rect 46 34 54 36
rect 42 33 54 34
rect 66 37 70 47
rect 66 35 67 37
rect 69 35 70 37
rect 66 31 70 35
rect 2 21 26 22
rect 2 19 22 21
rect 24 19 26 21
rect 2 18 26 19
rect 58 25 70 31
rect -2 11 82 12
rect -2 9 4 11
rect 6 9 82 11
rect -2 1 82 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 10 16 12 23
rect 17 16 19 23
rect 27 16 29 23
rect 37 16 39 23
rect 57 22 59 29
rect 69 17 71 24
<< pmos >>
rect 9 47 11 63
rect 19 47 21 70
rect 29 47 31 70
rect 36 47 38 70
rect 69 42 71 58
<< polyct0 >>
rect 11 40 13 42
rect 21 35 23 37
<< polyct1 >>
rect 54 50 56 52
rect 44 34 46 36
rect 67 35 69 37
<< ndifct0 >>
rect 52 24 54 26
rect 32 19 34 21
rect 42 18 44 20
rect 63 19 65 21
rect 74 20 76 22
<< ndifct1 >>
rect 22 19 24 21
rect 4 9 6 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 59 6 61
rect 24 49 26 51
rect 41 66 43 68
rect 74 51 76 53
rect 74 44 76 46
<< pdifct1 >>
rect 14 51 16 53
rect 63 69 65 71
<< alu0 >>
rect 39 66 41 68
rect 43 66 45 68
rect 39 65 45 66
rect 2 61 77 62
rect 2 59 4 61
rect 6 59 77 61
rect 2 58 77 59
rect 23 51 27 53
rect 23 49 24 51
rect 26 49 27 51
rect 23 46 27 49
rect 10 42 27 46
rect 10 40 11 42
rect 13 40 14 42
rect 10 30 14 40
rect 31 38 35 58
rect 19 37 35 38
rect 19 35 21 37
rect 23 35 35 37
rect 19 34 35 35
rect 73 53 77 58
rect 73 51 74 53
rect 76 51 77 53
rect 10 29 35 30
rect 10 26 55 29
rect 31 25 52 26
rect 31 21 35 25
rect 51 24 52 25
rect 54 24 55 26
rect 73 46 77 51
rect 73 44 74 46
rect 76 44 77 46
rect 51 22 55 24
rect 73 22 77 44
rect 61 21 67 22
rect 31 19 32 21
rect 34 19 35 21
rect 31 17 35 19
rect 40 20 46 21
rect 40 18 42 20
rect 44 18 46 20
rect 40 12 46 18
rect 61 19 63 21
rect 65 19 67 21
rect 51 12 55 16
rect 61 12 67 19
rect 73 20 74 22
rect 76 20 77 22
rect 73 18 77 20
<< labels >>
rlabel alu0 12 36 12 36 6 an
rlabel alu0 33 23 33 23 6 an
rlabel alu0 27 36 27 36 6 bn
rlabel alu0 25 47 25 47 6 an
rlabel ndifct0 53 25 53 25 6 an
rlabel alu0 39 60 39 60 6 bn
rlabel alu0 75 40 75 40 6 bn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 52 36 52 36 6 a2
rlabel alu1 44 44 44 44 6 a2
rlabel alu1 52 52 52 52 6 a1
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 28 60 28 6 b
rlabel polyct1 68 36 68 36 6 b
rlabel alu1 60 48 60 48 6 a1
<< end >>
