magic
tech scmos
timestamp 1199469049
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -5 48 95 105
<< pwell >>
rect -5 -5 95 48
<< poly >>
rect 15 94 17 98
rect 27 94 29 98
rect 39 94 41 98
rect 51 94 53 98
rect 63 94 65 98
rect 75 94 77 98
rect 15 52 17 55
rect 27 52 29 55
rect 39 52 41 55
rect 51 52 53 55
rect 63 52 65 55
rect 15 50 23 52
rect 27 50 41 52
rect 15 49 19 50
rect 17 48 19 49
rect 21 48 23 50
rect 17 46 23 48
rect 35 48 37 50
rect 39 48 41 50
rect 35 46 41 48
rect 47 50 65 52
rect 47 48 49 50
rect 51 48 53 50
rect 47 46 53 48
rect 75 48 77 55
rect 75 46 83 48
rect 37 39 39 46
rect 49 39 51 46
rect 75 44 79 46
rect 81 44 83 46
rect 57 42 83 44
rect 57 39 59 42
rect 37 12 39 17
rect 49 2 51 6
rect 57 2 59 6
<< ndif >>
rect 28 21 37 39
rect 28 19 31 21
rect 33 19 37 21
rect 28 17 37 19
rect 39 29 49 39
rect 39 27 43 29
rect 45 27 49 29
rect 39 21 49 27
rect 39 19 43 21
rect 45 19 49 21
rect 39 17 49 19
rect 44 6 49 17
rect 51 6 57 39
rect 59 20 68 39
rect 59 18 63 20
rect 65 18 68 20
rect 59 10 68 18
rect 59 8 63 10
rect 65 8 68 10
rect 59 6 68 8
<< pdif >>
rect 6 91 15 94
rect 6 89 9 91
rect 11 89 15 91
rect 6 81 15 89
rect 6 79 9 81
rect 11 79 15 81
rect 6 55 15 79
rect 17 81 27 94
rect 17 79 21 81
rect 23 79 27 81
rect 17 55 27 79
rect 29 71 39 94
rect 29 69 33 71
rect 35 69 39 71
rect 29 55 39 69
rect 41 80 51 94
rect 41 78 45 80
rect 47 78 51 80
rect 41 72 51 78
rect 41 70 45 72
rect 47 70 51 72
rect 41 55 51 70
rect 53 91 63 94
rect 53 89 57 91
rect 59 89 63 91
rect 53 81 63 89
rect 53 79 57 81
rect 59 79 63 81
rect 53 55 63 79
rect 65 80 75 94
rect 65 78 69 80
rect 71 78 75 80
rect 65 72 75 78
rect 65 70 69 72
rect 71 70 75 72
rect 65 55 75 70
rect 77 91 86 94
rect 77 89 81 91
rect 83 89 86 91
rect 77 81 86 89
rect 77 79 81 81
rect 83 79 86 81
rect 77 71 86 79
rect 77 69 81 71
rect 83 69 86 71
rect 77 55 86 69
<< alu1 >>
rect -2 91 92 100
rect -2 89 9 91
rect 11 89 57 91
rect 59 89 81 91
rect 83 89 92 91
rect -2 88 92 89
rect 8 81 12 88
rect 8 79 9 81
rect 11 79 12 81
rect 8 77 12 79
rect 19 81 48 82
rect 19 79 21 81
rect 23 80 48 81
rect 23 79 45 80
rect 19 78 45 79
rect 47 78 48 80
rect 8 71 37 73
rect 8 69 33 71
rect 35 69 37 71
rect 8 68 37 69
rect 44 72 48 78
rect 56 81 60 88
rect 56 79 57 81
rect 59 79 60 81
rect 56 77 60 79
rect 68 80 72 82
rect 68 78 69 80
rect 71 78 72 80
rect 68 72 72 78
rect 44 70 45 72
rect 47 70 69 72
rect 71 70 72 72
rect 44 68 72 70
rect 80 81 84 88
rect 80 79 81 81
rect 83 79 84 81
rect 80 71 84 79
rect 80 69 81 71
rect 83 69 84 71
rect 8 32 12 68
rect 80 67 84 69
rect 17 58 83 62
rect 17 50 23 58
rect 17 48 19 50
rect 21 48 23 50
rect 17 47 23 48
rect 28 50 42 53
rect 28 48 37 50
rect 39 48 42 50
rect 28 47 42 48
rect 47 50 62 53
rect 47 48 49 50
rect 51 48 62 50
rect 47 47 62 48
rect 38 37 42 47
rect 8 29 46 32
rect 8 27 43 29
rect 45 27 46 29
rect 58 27 62 47
rect 77 46 83 58
rect 77 44 79 46
rect 81 44 83 46
rect 77 38 83 44
rect 30 21 34 23
rect 30 19 31 21
rect 33 19 34 21
rect 30 12 34 19
rect 42 21 46 27
rect 42 19 43 21
rect 45 19 46 21
rect 42 17 46 19
rect 62 20 66 22
rect 62 18 63 20
rect 65 18 66 20
rect 62 12 66 18
rect -2 10 92 12
rect -2 8 63 10
rect 65 8 92 10
rect -2 7 92 8
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 92 7
rect -2 0 92 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< nmos >>
rect 37 17 39 39
rect 49 6 51 39
rect 57 6 59 39
<< pmos >>
rect 15 55 17 94
rect 27 55 29 94
rect 39 55 41 94
rect 51 55 53 94
rect 63 55 65 94
rect 75 55 77 94
<< polyct1 >>
rect 19 48 21 50
rect 37 48 39 50
rect 49 48 51 50
rect 79 44 81 46
<< ndifct1 >>
rect 31 19 33 21
rect 43 27 45 29
rect 43 19 45 21
rect 63 18 65 20
rect 63 8 65 10
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 9 89 11 91
rect 9 79 11 81
rect 21 79 23 81
rect 33 69 35 71
rect 45 78 47 80
rect 45 70 47 72
rect 57 89 59 91
rect 57 79 59 81
rect 69 78 71 80
rect 69 70 71 72
rect 81 89 83 91
rect 81 79 83 81
rect 81 69 83 71
<< labels >>
rlabel pdifct1 22 80 22 80 6 n2
rlabel pdifct1 46 71 46 71 6 n2
rlabel pdifct1 46 79 46 79 6 n2
rlabel pdifct1 70 71 70 71 6 n2
rlabel pdifct1 70 79 70 79 6 n2
rlabel alu1 10 50 10 50 6 z
rlabel alu1 20 30 20 30 6 z
rlabel alu1 40 45 40 45 6 b
rlabel alu1 40 30 40 30 6 z
rlabel alu1 30 30 30 30 6 z
rlabel alu1 30 50 30 50 6 b
rlabel alu1 20 55 20 55 6 a1
rlabel alu1 20 70 20 70 6 z
rlabel alu1 40 60 40 60 6 a1
rlabel alu1 30 70 30 70 6 z
rlabel alu1 30 60 30 60 6 a1
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 60 40 60 40 6 a2
rlabel alu1 50 50 50 50 6 a2
rlabel alu1 60 60 60 60 6 a1
rlabel alu1 50 60 50 60 6 a1
rlabel alu1 45 94 45 94 6 vdd
rlabel alu1 80 50 80 50 6 a1
rlabel alu1 70 60 70 60 6 a1
<< end >>
