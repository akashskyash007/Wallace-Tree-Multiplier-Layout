magic
tech scmos
timestamp 1199202200
<< ab >>
rect 0 0 144 80
<< nwell >>
rect -5 36 149 88
<< pwell >>
rect -5 -8 149 36
<< poly >>
rect 9 70 11 74
rect 55 72 111 74
rect 55 64 57 72
rect 65 64 67 68
rect 75 64 77 68
rect 82 64 84 72
rect 92 64 94 68
rect 99 64 101 68
rect 19 56 21 61
rect 38 58 40 63
rect 45 58 47 63
rect 9 38 11 42
rect 19 39 21 42
rect 9 36 15 38
rect 19 37 34 39
rect 9 34 11 36
rect 13 34 15 36
rect 9 32 15 34
rect 27 35 30 37
rect 32 35 34 37
rect 27 33 34 35
rect 9 28 11 32
rect 27 30 29 33
rect 38 23 40 52
rect 45 48 47 52
rect 45 46 51 48
rect 45 44 47 46
rect 49 44 51 46
rect 45 42 51 44
rect 55 38 57 52
rect 45 36 57 38
rect 45 23 47 36
rect 65 33 67 52
rect 75 48 77 58
rect 71 46 77 48
rect 71 44 73 46
rect 75 44 77 46
rect 71 42 77 44
rect 51 30 57 32
rect 51 28 53 30
rect 55 28 57 30
rect 51 26 57 28
rect 55 23 57 26
rect 65 31 71 33
rect 65 29 67 31
rect 69 29 71 31
rect 65 27 71 29
rect 65 23 67 27
rect 75 23 77 42
rect 82 38 84 58
rect 109 62 111 72
rect 129 63 131 68
rect 92 48 94 51
rect 88 46 94 48
rect 88 44 90 46
rect 92 44 94 46
rect 88 42 94 44
rect 99 39 101 51
rect 109 48 111 51
rect 129 49 131 53
rect 109 46 117 48
rect 115 39 117 46
rect 122 47 131 49
rect 122 45 124 47
rect 126 45 131 47
rect 122 43 131 45
rect 82 36 94 38
rect 82 30 88 32
rect 82 28 84 30
rect 86 28 88 30
rect 82 26 88 28
rect 82 23 84 26
rect 92 23 94 36
rect 99 37 105 39
rect 99 35 101 37
rect 103 35 105 37
rect 99 33 105 35
rect 115 37 121 39
rect 115 35 117 37
rect 119 35 121 37
rect 115 33 121 35
rect 99 23 101 33
rect 119 30 121 33
rect 129 30 131 43
rect 27 18 29 23
rect 119 19 121 24
rect 129 18 131 23
rect 9 11 11 14
rect 38 11 40 17
rect 45 12 47 17
rect 9 9 40 11
rect 55 8 57 17
rect 65 12 67 17
rect 75 12 77 17
rect 82 8 84 17
rect 92 12 94 17
rect 99 12 101 17
rect 55 6 84 8
<< ndif >>
rect 20 28 27 30
rect 2 26 9 28
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 4 14 9 22
rect 11 20 16 28
rect 20 26 22 28
rect 24 26 27 28
rect 20 24 27 26
rect 22 23 27 24
rect 29 23 36 30
rect 112 28 119 30
rect 112 26 114 28
rect 116 26 119 28
rect 112 24 119 26
rect 121 28 129 30
rect 121 26 124 28
rect 126 26 129 28
rect 121 24 129 26
rect 11 18 18 20
rect 31 21 38 23
rect 31 19 33 21
rect 35 19 38 21
rect 11 16 14 18
rect 16 16 18 18
rect 31 17 38 19
rect 40 17 45 23
rect 47 21 55 23
rect 47 19 50 21
rect 52 19 55 21
rect 47 17 55 19
rect 57 21 65 23
rect 57 19 60 21
rect 62 19 65 21
rect 57 17 65 19
rect 67 21 75 23
rect 67 19 70 21
rect 72 19 75 21
rect 67 17 75 19
rect 77 17 82 23
rect 84 21 92 23
rect 84 19 87 21
rect 89 19 92 21
rect 84 17 92 19
rect 94 17 99 23
rect 101 21 108 23
rect 101 19 104 21
rect 106 19 108 21
rect 123 23 129 24
rect 131 28 138 30
rect 131 26 134 28
rect 136 26 138 28
rect 131 23 138 26
rect 101 17 108 19
rect 11 14 18 16
<< pdif >>
rect 4 56 9 70
rect 2 53 9 56
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 18 70
rect 11 66 14 68
rect 16 66 18 68
rect 11 64 18 66
rect 11 56 17 64
rect 50 58 55 64
rect 30 56 38 58
rect 11 54 19 56
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 48 26 56
rect 30 54 32 56
rect 34 54 38 56
rect 30 52 38 54
rect 40 52 45 58
rect 47 56 55 58
rect 47 54 50 56
rect 52 54 55 56
rect 47 52 55 54
rect 57 56 65 64
rect 57 54 60 56
rect 62 54 65 56
rect 57 52 65 54
rect 67 62 75 64
rect 67 60 70 62
rect 72 60 75 62
rect 67 58 75 60
rect 77 58 82 64
rect 84 62 92 64
rect 84 60 87 62
rect 89 60 92 62
rect 84 58 92 60
rect 67 52 73 58
rect 21 46 28 48
rect 21 44 24 46
rect 26 44 28 46
rect 21 42 28 44
rect 87 51 92 58
rect 94 51 99 64
rect 101 62 106 64
rect 101 60 109 62
rect 101 58 104 60
rect 106 58 109 60
rect 101 51 109 58
rect 111 57 116 62
rect 122 61 129 63
rect 122 59 124 61
rect 126 59 129 61
rect 111 55 118 57
rect 111 53 114 55
rect 116 53 118 55
rect 122 53 129 59
rect 131 59 136 63
rect 131 57 138 59
rect 131 55 134 57
rect 136 55 138 57
rect 131 53 138 55
rect 111 51 118 53
<< alu1 >>
rect -2 81 146 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 146 81
rect -2 68 146 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 15 46
rect 2 42 15 44
rect 2 28 6 42
rect 2 26 7 28
rect 2 24 4 26
rect 6 24 7 26
rect 2 22 7 24
rect 121 47 127 54
rect 121 46 124 47
rect 97 38 103 46
rect 113 45 124 46
rect 126 45 127 47
rect 113 42 127 45
rect 97 37 111 38
rect 97 35 101 37
rect 103 35 111 37
rect 97 34 111 35
rect -2 1 146 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 146 1
rect -2 -2 146 -1
<< ptie >>
rect 0 1 144 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 144 1
rect 0 -3 144 -1
<< ntie >>
rect 0 81 144 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 144 81
rect 0 77 144 79
<< nmos >>
rect 9 14 11 28
rect 27 23 29 30
rect 119 24 121 30
rect 38 17 40 23
rect 45 17 47 23
rect 55 17 57 23
rect 65 17 67 23
rect 75 17 77 23
rect 82 17 84 23
rect 92 17 94 23
rect 99 17 101 23
rect 129 23 131 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 56
rect 38 52 40 58
rect 45 52 47 58
rect 55 52 57 64
rect 65 52 67 64
rect 75 58 77 64
rect 82 58 84 64
rect 92 51 94 64
rect 99 51 101 64
rect 109 51 111 62
rect 129 53 131 63
<< polyct0 >>
rect 11 34 13 36
rect 30 35 32 37
rect 47 44 49 46
rect 73 44 75 46
rect 53 28 55 30
rect 67 29 69 31
rect 90 44 92 46
rect 84 28 86 30
rect 117 35 119 37
<< polyct1 >>
rect 124 45 126 47
rect 101 35 103 37
<< ndifct0 >>
rect 22 26 24 28
rect 114 26 116 28
rect 124 26 126 28
rect 33 19 35 21
rect 14 16 16 18
rect 50 19 52 21
rect 60 19 62 21
rect 70 19 72 21
rect 87 19 89 21
rect 104 19 106 21
rect 134 26 136 28
<< ndifct1 >>
rect 4 24 6 26
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
<< pdifct0 >>
rect 14 66 16 68
rect 14 52 16 54
rect 32 54 34 56
rect 50 54 52 56
rect 60 54 62 56
rect 70 60 72 62
rect 87 60 89 62
rect 24 44 26 46
rect 104 58 106 60
rect 124 59 126 61
rect 114 53 116 55
rect 134 55 136 57
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 13 66 14 68
rect 16 66 17 68
rect 13 54 17 66
rect 13 52 14 54
rect 16 52 17 54
rect 31 56 35 68
rect 69 62 73 68
rect 69 60 70 62
rect 72 60 73 62
rect 69 58 73 60
rect 81 62 91 63
rect 81 60 87 62
rect 89 60 91 62
rect 81 59 91 60
rect 102 60 108 68
rect 31 54 32 56
rect 34 54 35 56
rect 31 52 35 54
rect 38 56 54 57
rect 38 54 50 56
rect 52 54 54 56
rect 38 53 54 54
rect 59 56 63 58
rect 59 54 60 56
rect 62 54 63 56
rect 13 50 17 52
rect 21 46 28 47
rect 21 44 24 46
rect 26 44 28 46
rect 21 43 28 44
rect 21 37 25 43
rect 38 38 42 53
rect 59 47 63 54
rect 45 46 54 47
rect 45 44 47 46
rect 49 44 54 46
rect 45 43 54 44
rect 9 36 25 37
rect 9 34 11 36
rect 13 34 25 36
rect 28 37 44 38
rect 28 35 30 37
rect 32 35 44 37
rect 28 34 44 35
rect 9 33 25 34
rect 21 28 25 33
rect 21 26 22 28
rect 24 26 25 28
rect 21 24 25 26
rect 32 21 36 23
rect 13 18 17 20
rect 13 16 14 18
rect 16 16 17 18
rect 13 12 17 16
rect 32 19 33 21
rect 35 19 36 21
rect 32 12 36 19
rect 40 22 44 34
rect 50 32 54 43
rect 59 46 77 47
rect 59 44 73 46
rect 75 44 77 46
rect 59 43 77 44
rect 50 30 56 32
rect 50 28 53 30
rect 55 28 56 30
rect 50 26 56 28
rect 40 21 54 22
rect 40 19 50 21
rect 52 19 54 21
rect 40 18 54 19
rect 59 21 63 43
rect 81 40 85 59
rect 102 58 104 60
rect 106 58 108 60
rect 122 61 128 68
rect 122 59 124 61
rect 126 59 128 61
rect 122 58 128 59
rect 102 57 108 58
rect 133 57 137 59
rect 113 55 117 57
rect 113 54 114 55
rect 76 36 85 40
rect 89 53 114 54
rect 116 53 117 55
rect 133 55 134 57
rect 136 55 137 57
rect 89 50 117 53
rect 89 46 93 50
rect 89 44 90 46
rect 92 44 93 46
rect 76 33 80 36
rect 66 31 80 33
rect 89 32 93 44
rect 133 38 137 55
rect 115 37 137 38
rect 115 35 117 37
rect 119 35 137 37
rect 115 34 137 35
rect 66 29 67 31
rect 69 29 80 31
rect 66 27 80 29
rect 59 19 60 21
rect 62 19 63 21
rect 59 17 63 19
rect 69 21 73 23
rect 69 19 70 21
rect 72 19 73 21
rect 69 12 73 19
rect 76 22 80 27
rect 83 30 93 32
rect 83 28 84 30
rect 86 28 118 30
rect 83 26 114 28
rect 116 26 118 28
rect 112 25 118 26
rect 123 28 127 30
rect 123 26 124 28
rect 126 26 127 28
rect 76 21 91 22
rect 76 19 87 21
rect 89 19 91 21
rect 76 18 91 19
rect 102 21 108 22
rect 102 19 104 21
rect 106 19 108 21
rect 102 12 108 19
rect 123 12 127 26
rect 133 28 137 34
rect 133 26 134 28
rect 136 26 137 28
rect 133 24 137 26
<< labels >>
rlabel alu0 23 35 23 35 6 zn
rlabel alu0 17 35 17 35 6 zn
rlabel alu0 24 45 24 45 6 zn
rlabel alu0 47 20 47 20 6 n4
rlabel alu0 53 29 53 29 6 ci
rlabel alu0 36 36 36 36 6 n4
rlabel alu0 49 45 49 45 6 ci
rlabel alu0 46 55 46 55 6 n4
rlabel alu0 73 30 73 30 6 n1
rlabel alu0 68 45 68 45 6 n2
rlabel alu0 61 37 61 37 6 n2
rlabel alu0 83 20 83 20 6 n1
rlabel alu0 91 40 91 40 6 ci
rlabel alu0 86 61 86 61 6 n1
rlabel alu0 100 28 100 28 6 ci
rlabel alu0 126 36 126 36 6 cn
rlabel alu0 103 52 103 52 6 ci
rlabel alu0 135 41 135 41 6 cn
rlabel alu1 12 44 12 44 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 72 6 72 6 6 vss
rlabel alu1 100 40 100 40 6 d
rlabel alu1 72 74 72 74 6 vdd
rlabel alu1 108 36 108 36 6 d
rlabel alu1 116 44 116 44 6 cp
rlabel alu1 124 48 124 48 6 cp
<< end >>
