magic
tech scmos
timestamp 1199202906
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 12 39 14 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 36 21 42
rect 19 34 25 36
rect 10 24 12 33
rect 19 32 21 34
rect 23 32 25 34
rect 19 30 25 32
rect 21 27 23 30
rect 10 11 12 16
rect 21 15 23 19
<< ndif >>
rect 16 24 21 27
rect 2 16 10 24
rect 12 20 21 24
rect 12 18 15 20
rect 17 19 21 20
rect 23 23 30 27
rect 23 21 26 23
rect 28 21 30 23
rect 23 19 30 21
rect 17 18 19 19
rect 12 16 19 18
rect 2 11 8 16
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
<< pdif >>
rect 7 63 12 70
rect 5 61 12 63
rect 5 59 7 61
rect 9 59 12 61
rect 5 54 12 59
rect 5 52 7 54
rect 9 52 12 54
rect 5 50 12 52
rect 7 42 12 50
rect 14 42 19 70
rect 21 68 30 70
rect 21 66 26 68
rect 28 66 30 68
rect 21 61 30 66
rect 21 59 26 61
rect 28 59 30 61
rect 21 42 30 59
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 5 61 11 62
rect 5 59 7 61
rect 9 59 11 61
rect 5 55 11 59
rect 2 54 11 55
rect 2 52 7 54
rect 9 52 11 54
rect 2 51 11 52
rect 2 23 6 51
rect 18 43 22 47
rect 10 39 22 43
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 26 35 30 39
rect 10 33 14 35
rect 18 34 30 35
rect 18 32 21 34
rect 23 32 30 34
rect 18 31 30 32
rect 18 25 22 31
rect 2 21 14 23
rect 2 20 19 21
rect 2 18 15 20
rect 17 18 19 20
rect 2 17 19 18
rect -2 11 34 12
rect -2 9 4 11
rect 6 9 34 11
rect -2 1 34 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 10 16 12 24
rect 21 19 23 27
<< pmos >>
rect 12 42 14 70
rect 19 42 21 70
<< polyct1 >>
rect 11 35 13 37
rect 21 32 23 34
<< ndifct0 >>
rect 26 21 28 23
<< ndifct1 >>
rect 15 18 17 20
rect 4 9 6 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 26 66 28 68
rect 26 59 28 61
<< pdifct1 >>
rect 7 59 9 61
rect 7 52 9 54
<< alu0 >>
rect 25 66 26 68
rect 28 66 29 68
rect 25 61 29 66
rect 25 59 26 61
rect 28 59 29 61
rect 25 57 29 59
rect 25 23 29 25
rect 25 21 26 23
rect 28 21 29 23
rect 25 12 29 21
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 44 20 44 6 b
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 36 28 36 6 a
<< end >>
