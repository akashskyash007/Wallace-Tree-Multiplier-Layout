magic
tech scmos
timestamp 1199469451
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -2 48 82 104
<< pwell >>
rect -2 -4 82 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 31 94 33 98
rect 43 94 45 98
rect 55 94 57 98
rect 67 94 69 98
rect 11 53 13 56
rect 23 53 25 56
rect 11 51 25 53
rect 11 49 19 51
rect 21 50 25 51
rect 31 53 33 56
rect 43 53 45 56
rect 31 51 39 53
rect 31 50 35 51
rect 21 49 23 50
rect 11 47 23 49
rect 11 33 13 47
rect 21 33 23 47
rect 29 49 35 50
rect 37 49 39 51
rect 29 47 39 49
rect 43 51 51 53
rect 43 49 47 51
rect 49 49 51 51
rect 43 47 51 49
rect 29 33 31 47
rect 43 40 45 47
rect 55 43 57 56
rect 41 37 45 40
rect 49 41 57 43
rect 49 39 51 41
rect 53 40 57 41
rect 53 39 55 40
rect 49 37 55 39
rect 41 33 43 37
rect 53 26 55 37
rect 67 36 69 56
rect 59 34 69 36
rect 59 32 61 34
rect 63 33 69 34
rect 63 32 67 33
rect 59 30 67 32
rect 65 26 67 30
rect 11 11 13 16
rect 21 11 23 16
rect 29 11 31 16
rect 41 11 43 16
rect 53 4 55 9
rect 65 2 67 7
<< ndif >>
rect 3 31 11 33
rect 3 29 5 31
rect 7 29 11 31
rect 3 23 11 29
rect 3 21 5 23
rect 7 21 11 23
rect 3 19 11 21
rect 6 16 11 19
rect 13 16 21 33
rect 23 16 29 33
rect 31 31 41 33
rect 31 29 35 31
rect 37 29 41 31
rect 31 16 41 29
rect 43 26 48 33
rect 43 21 53 26
rect 43 19 47 21
rect 49 19 53 21
rect 43 16 53 19
rect 15 9 19 16
rect 48 9 53 16
rect 55 21 65 26
rect 55 19 59 21
rect 61 19 65 21
rect 55 11 65 19
rect 55 9 59 11
rect 61 9 65 11
rect 13 7 19 9
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
rect 57 7 65 9
rect 67 23 72 26
rect 67 21 75 23
rect 67 19 71 21
rect 73 19 75 21
rect 67 17 75 19
rect 67 7 72 17
<< pdif >>
rect 6 81 11 94
rect 3 79 11 81
rect 3 77 5 79
rect 7 77 11 79
rect 3 71 11 77
rect 3 69 5 71
rect 7 69 11 71
rect 3 67 11 69
rect 6 56 11 67
rect 13 91 23 94
rect 13 89 17 91
rect 19 89 23 91
rect 13 56 23 89
rect 25 56 31 94
rect 33 71 43 94
rect 33 69 37 71
rect 39 69 43 71
rect 33 56 43 69
rect 45 81 55 94
rect 45 79 49 81
rect 51 79 55 81
rect 45 56 55 79
rect 57 91 67 94
rect 57 89 61 91
rect 63 89 67 91
rect 57 81 67 89
rect 57 79 61 81
rect 63 79 67 81
rect 57 56 67 79
rect 69 74 74 94
rect 69 72 77 74
rect 69 70 73 72
rect 75 70 77 72
rect 69 64 77 70
rect 69 62 73 64
rect 75 62 77 64
rect 69 60 77 62
rect 69 56 74 60
<< alu1 >>
rect -2 91 82 100
rect -2 89 17 91
rect 19 89 61 91
rect 63 89 82 91
rect -2 88 82 89
rect 4 81 53 82
rect 4 79 49 81
rect 51 79 53 81
rect 4 77 5 79
rect 7 78 53 79
rect 60 81 64 88
rect 60 79 61 81
rect 63 79 64 81
rect 7 77 8 78
rect 60 77 64 79
rect 4 71 8 77
rect 68 72 77 73
rect 4 69 5 71
rect 7 69 8 71
rect 4 67 8 69
rect 26 71 41 72
rect 26 69 37 71
rect 39 69 41 71
rect 26 68 41 69
rect 46 68 63 72
rect 68 70 73 72
rect 75 70 77 72
rect 68 69 77 70
rect 8 53 12 63
rect 8 51 22 53
rect 8 49 19 51
rect 21 49 22 51
rect 8 47 22 49
rect 8 37 12 47
rect 4 31 8 33
rect 4 29 5 31
rect 7 29 8 31
rect 4 23 8 29
rect 26 32 30 68
rect 38 53 42 63
rect 34 51 42 53
rect 34 49 35 51
rect 37 49 42 51
rect 34 47 42 49
rect 46 51 52 68
rect 68 65 72 69
rect 68 64 77 65
rect 68 62 73 64
rect 75 62 77 64
rect 68 61 77 62
rect 68 52 72 61
rect 46 49 47 51
rect 49 49 52 51
rect 46 47 52 49
rect 57 48 72 52
rect 38 43 42 47
rect 38 41 55 43
rect 38 39 51 41
rect 53 39 55 41
rect 38 37 55 39
rect 60 34 64 36
rect 60 32 61 34
rect 63 32 64 34
rect 26 31 64 32
rect 26 29 35 31
rect 37 29 64 31
rect 26 28 64 29
rect 68 23 72 48
rect 4 21 5 23
rect 7 22 8 23
rect 7 21 51 22
rect 4 19 47 21
rect 49 19 51 21
rect 4 18 51 19
rect 58 21 62 23
rect 58 19 59 21
rect 61 19 62 21
rect 58 12 62 19
rect 68 21 74 23
rect 68 19 71 21
rect 73 19 74 21
rect 68 17 74 19
rect -2 11 82 12
rect -2 9 59 11
rect 61 9 82 11
rect -2 7 82 9
rect -2 5 15 7
rect 17 5 27 7
rect 29 5 37 7
rect 39 5 82 7
rect -2 0 82 5
<< ptie >>
rect 25 7 41 9
rect 25 5 27 7
rect 29 5 37 7
rect 39 5 41 7
rect 25 3 41 5
<< nmos >>
rect 11 16 13 33
rect 21 16 23 33
rect 29 16 31 33
rect 41 16 43 33
rect 53 9 55 26
rect 65 7 67 26
<< pmos >>
rect 11 56 13 94
rect 23 56 25 94
rect 31 56 33 94
rect 43 56 45 94
rect 55 56 57 94
rect 67 56 69 94
<< polyct1 >>
rect 19 49 21 51
rect 35 49 37 51
rect 47 49 49 51
rect 51 39 53 41
rect 61 32 63 34
<< ndifct1 >>
rect 5 29 7 31
rect 5 21 7 23
rect 35 29 37 31
rect 47 19 49 21
rect 59 19 61 21
rect 59 9 61 11
rect 15 5 17 7
rect 71 19 73 21
<< ptiect1 >>
rect 27 5 29 7
rect 37 5 39 7
<< pdifct1 >>
rect 5 77 7 79
rect 5 69 7 71
rect 17 89 19 91
rect 37 69 39 71
rect 49 79 51 81
rect 61 89 63 91
rect 61 79 63 81
rect 73 70 75 72
rect 73 62 75 64
<< labels >>
rlabel alu1 6 25 6 25 6 n4
rlabel alu1 10 50 10 50 6 a
rlabel alu1 6 74 6 74 6 n2
rlabel polyct1 20 50 20 50 6 a
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 40 50 40 50 6 b
rlabel alu1 33 70 33 70 6 zn
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 27 20 27 20 6 n4
rlabel alu1 45 30 45 30 6 zn
rlabel alu1 62 32 62 32 6 zn
rlabel alu1 50 40 50 40 6 b
rlabel alu1 60 50 60 50 6 z
rlabel alu1 50 60 50 60 6 c
rlabel alu1 60 70 60 70 6 c
rlabel alu1 28 80 28 80 6 n2
rlabel alu1 70 45 70 45 6 z
<< end >>
