magic
tech scmos
timestamp 1199202459
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 13 70 15 74
rect 20 70 22 74
rect 30 70 32 74
rect 37 70 39 74
rect 49 70 51 74
rect 56 70 58 74
rect 66 70 68 74
rect 73 70 75 74
rect 85 60 87 65
rect 13 42 15 45
rect 2 40 15 42
rect 20 42 22 45
rect 30 42 32 45
rect 20 40 33 42
rect 2 38 4 40
rect 6 38 13 40
rect 2 36 13 38
rect 27 38 29 40
rect 31 38 33 40
rect 27 36 33 38
rect 11 27 13 36
rect 17 34 23 36
rect 17 32 19 34
rect 21 32 23 34
rect 37 32 39 45
rect 49 42 51 45
rect 47 40 51 42
rect 56 42 58 45
rect 66 42 68 45
rect 56 40 69 42
rect 47 36 49 40
rect 63 38 65 40
rect 67 38 69 40
rect 63 36 69 38
rect 73 39 75 45
rect 73 37 79 39
rect 17 30 30 32
rect 18 27 20 30
rect 28 27 30 30
rect 35 30 39 32
rect 43 34 49 36
rect 43 32 45 34
rect 47 32 49 34
rect 43 30 49 32
rect 53 34 59 36
rect 53 32 55 34
rect 57 32 59 34
rect 73 35 75 37
rect 77 35 79 37
rect 85 36 87 42
rect 73 33 79 35
rect 83 33 87 36
rect 73 32 75 33
rect 53 30 66 32
rect 35 27 37 30
rect 47 27 49 30
rect 54 27 56 30
rect 64 27 66 30
rect 71 30 75 32
rect 83 30 85 33
rect 71 27 73 30
rect 11 8 13 16
rect 18 12 20 16
rect 28 12 30 16
rect 35 8 37 16
rect 11 6 37 8
rect 47 11 49 16
rect 54 11 56 16
rect 64 8 66 16
rect 71 12 73 16
rect 83 8 85 21
rect 64 6 85 8
<< ndif >>
rect 78 27 83 30
rect 2 20 11 27
rect 2 18 4 20
rect 6 18 11 20
rect 2 16 11 18
rect 13 16 18 27
rect 20 21 28 27
rect 20 19 23 21
rect 25 19 28 21
rect 20 16 28 19
rect 30 16 35 27
rect 37 16 47 27
rect 49 16 54 27
rect 56 20 64 27
rect 56 18 59 20
rect 61 18 64 20
rect 56 16 64 18
rect 66 16 71 27
rect 73 25 83 27
rect 73 23 78 25
rect 80 23 83 25
rect 73 21 83 23
rect 85 28 92 30
rect 85 26 88 28
rect 90 26 92 28
rect 85 24 92 26
rect 85 21 90 24
rect 73 16 81 21
rect 39 11 45 16
rect 39 9 41 11
rect 43 9 45 11
rect 39 7 45 9
<< pdif >>
rect 5 68 13 70
rect 5 66 8 68
rect 10 66 13 68
rect 5 45 13 66
rect 15 45 20 70
rect 22 61 30 70
rect 22 59 25 61
rect 27 59 30 61
rect 22 45 30 59
rect 32 45 37 70
rect 39 68 49 70
rect 39 66 43 68
rect 45 66 49 68
rect 39 45 49 66
rect 51 45 56 70
rect 58 61 66 70
rect 58 59 61 61
rect 63 59 66 61
rect 58 45 66 59
rect 68 45 73 70
rect 75 61 83 70
rect 75 59 79 61
rect 81 60 83 61
rect 81 59 85 60
rect 75 54 85 59
rect 75 52 79 54
rect 81 52 85 54
rect 75 45 85 52
rect 77 42 85 45
rect 87 55 92 60
rect 87 53 94 55
rect 87 51 90 53
rect 92 51 94 53
rect 87 46 94 51
rect 87 44 90 46
rect 92 44 94 46
rect 87 42 94 44
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 2 58 15 62
rect 21 61 65 62
rect 21 59 25 61
rect 27 59 61 61
rect 63 59 65 61
rect 21 58 65 59
rect 2 40 6 58
rect 2 38 4 40
rect 2 33 6 38
rect 10 22 14 47
rect 33 42 56 46
rect 33 34 39 42
rect 52 35 56 42
rect 73 37 79 38
rect 73 35 75 37
rect 77 35 79 37
rect 52 34 59 35
rect 52 32 55 34
rect 57 32 59 34
rect 73 33 79 35
rect 52 31 59 32
rect 41 26 47 30
rect 65 29 79 33
rect 65 26 71 29
rect 10 21 31 22
rect 10 19 23 21
rect 25 19 31 21
rect 10 18 31 19
rect -2 11 98 12
rect -2 9 41 11
rect 43 9 98 11
rect -2 1 98 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 11 16 13 27
rect 18 16 20 27
rect 28 16 30 27
rect 35 16 37 27
rect 47 16 49 27
rect 54 16 56 27
rect 64 16 66 27
rect 71 16 73 27
rect 83 21 85 30
<< pmos >>
rect 13 45 15 70
rect 20 45 22 70
rect 30 45 32 70
rect 37 45 39 70
rect 49 45 51 70
rect 56 45 58 70
rect 66 45 68 70
rect 73 45 75 70
rect 85 42 87 60
<< polyct0 >>
rect 29 38 31 40
rect 19 32 21 34
rect 65 38 67 40
rect 45 32 47 34
<< polyct1 >>
rect 4 38 6 40
rect 55 32 57 34
rect 75 35 77 37
<< ndifct0 >>
rect 4 18 6 20
rect 59 18 61 20
rect 78 23 80 25
rect 88 26 90 28
<< ndifct1 >>
rect 23 19 25 21
rect 41 9 43 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 8 66 10 68
rect 43 66 45 68
rect 79 59 81 61
rect 79 52 81 54
rect 90 51 92 53
rect 90 44 92 46
<< pdifct1 >>
rect 25 59 27 61
rect 61 59 63 61
<< alu0 >>
rect 6 66 8 68
rect 10 66 12 68
rect 6 65 12 66
rect 41 66 43 68
rect 45 66 47 68
rect 41 65 47 66
rect 19 58 21 62
rect 78 61 82 68
rect 78 59 79 61
rect 81 59 82 61
rect 19 55 23 58
rect 11 51 23 55
rect 78 54 82 59
rect 11 47 15 51
rect 26 50 68 54
rect 78 52 79 54
rect 81 52 82 54
rect 78 50 82 52
rect 89 53 93 55
rect 89 51 90 53
rect 92 51 93 53
rect 26 48 30 50
rect 6 36 7 42
rect 14 43 15 47
rect 20 44 30 48
rect 64 46 68 50
rect 89 46 93 51
rect 20 35 24 44
rect 27 40 33 41
rect 27 38 29 40
rect 31 38 33 40
rect 27 37 33 38
rect 17 34 24 35
rect 44 34 48 36
rect 17 32 19 34
rect 21 32 24 34
rect 17 31 24 32
rect 44 32 45 34
rect 47 32 48 34
rect 44 30 48 32
rect 64 44 90 46
rect 92 44 94 46
rect 64 42 94 44
rect 64 40 68 42
rect 64 38 65 40
rect 67 38 68 40
rect 64 36 68 38
rect 47 28 48 30
rect 90 29 94 42
rect 47 26 65 28
rect 86 28 94 29
rect 86 26 88 28
rect 90 26 94 28
rect 44 24 69 26
rect 76 25 82 26
rect 86 25 94 26
rect 76 23 78 25
rect 80 23 82 25
rect 3 20 7 22
rect 3 18 4 20
rect 6 18 7 20
rect 31 20 64 21
rect 31 18 59 20
rect 61 18 64 20
rect 3 12 7 18
rect 27 17 64 18
rect 76 12 82 23
<< labels >>
rlabel alu0 22 39 22 39 6 sn
rlabel alu0 91 48 91 48 6 sn
rlabel alu0 92 35 92 35 6 sn
rlabel alu0 79 44 79 44 6 sn
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 36 12 36 6 z
rlabel alu1 4 44 4 44 6 a0
rlabel alu1 12 60 12 60 6 a0
rlabel alu1 28 20 28 20 6 z
rlabel alu1 44 28 44 28 6 a1
rlabel alu1 36 40 36 40 6 s
rlabel alu1 44 44 44 44 6 s
rlabel alu1 28 60 28 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 68 28 68 28 6 a1
rlabel alu1 52 44 52 44 6 s
rlabel alu1 60 60 60 60 6 z
rlabel alu1 52 60 52 60 6 z
rlabel alu1 48 74 48 74 6 vdd
rlabel polyct1 76 36 76 36 6 a1
<< end >>
