magic
tech scmos
timestamp 1199203088
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 12 66 14 70
rect 22 66 24 70
rect 29 66 31 70
rect 12 45 14 51
rect 9 43 15 45
rect 9 41 11 43
rect 13 41 15 43
rect 9 39 15 41
rect 9 19 11 39
rect 39 64 41 68
rect 39 43 41 46
rect 39 41 55 43
rect 49 39 51 41
rect 53 39 55 41
rect 22 35 24 38
rect 17 33 24 35
rect 17 31 19 33
rect 21 31 24 33
rect 17 29 24 31
rect 29 35 31 38
rect 49 37 55 39
rect 29 33 35 35
rect 29 31 31 33
rect 33 31 35 33
rect 29 29 35 31
rect 19 19 21 29
rect 29 19 31 29
rect 49 26 51 37
rect 49 12 51 17
rect 9 2 11 6
rect 19 2 21 6
rect 29 2 31 6
<< ndif >>
rect 42 24 49 26
rect 42 22 44 24
rect 46 22 49 24
rect 42 20 49 22
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 6 9 13
rect 11 17 19 19
rect 11 15 14 17
rect 16 15 19 17
rect 11 6 19 15
rect 21 10 29 19
rect 21 8 24 10
rect 26 8 29 10
rect 21 6 29 8
rect 31 17 38 19
rect 44 17 49 20
rect 51 21 58 26
rect 51 19 54 21
rect 56 19 58 21
rect 51 17 58 19
rect 31 15 34 17
rect 36 15 38 17
rect 31 13 38 15
rect 31 6 36 13
<< pdif >>
rect 4 64 12 66
rect 4 62 7 64
rect 9 62 12 64
rect 4 51 12 62
rect 14 57 22 66
rect 14 55 17 57
rect 19 55 22 57
rect 14 51 22 55
rect 17 38 22 51
rect 24 38 29 66
rect 31 64 37 66
rect 31 62 39 64
rect 31 60 34 62
rect 36 60 39 62
rect 31 55 39 60
rect 31 53 34 55
rect 36 53 39 55
rect 31 46 39 53
rect 41 59 46 64
rect 41 57 48 59
rect 41 55 44 57
rect 46 55 48 57
rect 41 50 48 55
rect 41 48 44 50
rect 46 48 48 50
rect 41 46 48 48
rect 31 38 37 46
<< alu1 >>
rect -2 67 66 72
rect -2 65 56 67
rect 58 65 66 67
rect -2 64 66 65
rect 2 57 23 58
rect 2 55 17 57
rect 19 55 23 57
rect 2 54 23 55
rect 2 18 6 54
rect 10 43 14 45
rect 10 41 11 43
rect 13 41 14 43
rect 58 43 62 51
rect 10 26 14 41
rect 25 33 39 34
rect 25 31 31 33
rect 33 31 39 33
rect 25 30 39 31
rect 10 22 23 26
rect 33 22 39 30
rect 50 41 62 43
rect 50 39 51 41
rect 53 39 62 41
rect 50 37 62 39
rect 2 17 8 18
rect 2 15 4 17
rect 6 15 8 17
rect 2 13 8 15
rect -2 7 66 8
rect -2 5 48 7
rect 50 5 56 7
rect 58 5 66 7
rect -2 0 66 5
<< ptie >>
rect 46 7 60 9
rect 46 5 48 7
rect 50 5 56 7
rect 58 5 60 7
rect 46 3 60 5
<< ntie >>
rect 54 67 60 69
rect 54 65 56 67
rect 58 65 60 67
rect 54 46 60 65
<< nmos >>
rect 9 6 11 19
rect 19 6 21 19
rect 29 6 31 19
rect 49 17 51 26
<< pmos >>
rect 12 51 14 66
rect 22 38 24 66
rect 29 38 31 66
rect 39 46 41 64
<< polyct0 >>
rect 19 31 21 33
<< polyct1 >>
rect 11 41 13 43
rect 51 39 53 41
rect 31 31 33 33
<< ndifct0 >>
rect 44 22 46 24
rect 14 15 16 17
rect 24 8 26 10
rect 54 19 56 21
rect 34 15 36 17
<< ndifct1 >>
rect 4 15 6 17
<< ntiect1 >>
rect 56 65 58 67
<< ptiect1 >>
rect 48 5 50 7
rect 56 5 58 7
<< pdifct0 >>
rect 7 62 9 64
rect 34 60 36 62
rect 34 53 36 55
rect 44 55 46 57
rect 44 48 46 50
<< pdifct1 >>
rect 17 55 19 57
<< alu0 >>
rect 5 62 7 64
rect 9 62 11 64
rect 5 61 11 62
rect 33 62 37 64
rect 33 60 34 62
rect 36 60 37 62
rect 33 55 37 60
rect 33 53 34 55
rect 36 53 37 55
rect 33 51 37 53
rect 43 57 47 59
rect 43 55 44 57
rect 46 55 47 57
rect 43 50 47 55
rect 43 48 44 50
rect 46 48 47 50
rect 43 42 47 48
rect 18 38 47 42
rect 18 33 22 38
rect 18 31 19 33
rect 21 31 22 33
rect 18 29 22 31
rect 43 24 47 38
rect 43 22 44 24
rect 46 22 47 24
rect 43 20 47 22
rect 53 21 57 23
rect 53 19 54 21
rect 56 19 57 21
rect 12 17 38 18
rect 12 15 14 17
rect 16 15 34 17
rect 36 15 38 17
rect 12 14 38 15
rect 22 10 28 11
rect 22 8 24 10
rect 26 8 28 10
rect 53 8 57 19
<< labels >>
rlabel alu0 25 16 25 16 6 n1
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 36 12 36 6 b
rlabel alu1 12 56 12 56 6 z
rlabel alu1 20 24 20 24 6 b
rlabel alu1 28 32 28 32 6 a1
rlabel alu1 20 56 20 56 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 32 68 32 68 6 vdd
rlabel polyct1 52 40 52 40 6 a2
rlabel alu1 60 44 60 44 6 a2
<< end >>
