magic
tech scmos
timestamp 1199201690
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 20 58 22 63
rect 30 58 32 63
rect 9 39 11 42
rect 20 39 22 50
rect 30 47 32 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 30 11 33
rect 22 25 24 33
rect 29 25 31 41
rect 9 11 11 16
rect 22 13 24 18
rect 29 13 31 18
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 20 9 26
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 25 19 30
rect 11 18 22 25
rect 24 18 29 25
rect 31 22 38 25
rect 31 20 34 22
rect 36 20 38 22
rect 31 18 38 20
rect 11 16 19 18
rect 13 11 19 16
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 18 70
rect 11 66 14 68
rect 16 66 18 68
rect 11 61 18 66
rect 32 69 38 71
rect 32 67 34 69
rect 36 67 38 69
rect 32 65 38 67
rect 11 59 14 61
rect 16 59 18 61
rect 11 58 18 59
rect 34 58 38 65
rect 11 50 20 58
rect 22 54 30 58
rect 22 52 25 54
rect 27 52 30 54
rect 22 50 30 52
rect 32 50 38 58
rect 11 42 18 50
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 69 42 79
rect -2 68 34 69
rect 36 68 42 69
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 2 28 6 42
rect 34 46 38 55
rect 25 45 38 46
rect 25 43 31 45
rect 33 43 38 45
rect 25 42 38 43
rect 17 37 31 38
rect 17 35 21 37
rect 23 35 31 37
rect 17 34 31 35
rect 2 26 4 28
rect 2 23 6 26
rect 25 26 31 34
rect 2 20 14 23
rect 2 18 4 20
rect 6 18 14 20
rect 2 17 14 18
rect -2 11 42 12
rect -2 9 15 11
rect 17 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 16 11 30
rect 22 18 24 25
rect 29 18 31 25
<< pmos >>
rect 9 42 11 70
rect 20 50 22 58
rect 30 50 32 58
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 21 35 23 37
<< ndifct0 >>
rect 34 20 36 22
<< ndifct1 >>
rect 4 26 6 28
rect 4 18 6 20
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 66 16 68
rect 34 67 36 68
rect 14 59 16 61
rect 25 52 27 54
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 34 68 36 69
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 32 67 34 68
rect 36 67 38 68
rect 32 66 38 67
rect 12 61 18 66
rect 12 59 14 61
rect 16 59 18 61
rect 12 58 18 59
rect 10 54 29 55
rect 10 52 25 54
rect 27 52 29 54
rect 10 51 29 52
rect 10 37 14 51
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 6 23 7 30
rect 10 26 22 30
rect 18 23 22 26
rect 18 22 38 23
rect 18 20 34 22
rect 36 20 38 22
rect 18 19 38 20
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 19 53 19 53 6 zn
rlabel alu0 28 21 28 21 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 52 36 52 6 b
<< end >>
