magic
tech scmos
timestamp 1199203285
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 22 70 24 74
rect 29 70 31 74
rect 36 70 38 74
rect 9 39 11 42
rect 22 39 24 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 29 11 33
rect 19 23 21 33
rect 29 32 31 42
rect 36 39 38 42
rect 36 37 49 39
rect 41 35 45 37
rect 47 35 49 37
rect 41 33 49 35
rect 29 30 37 32
rect 29 28 33 30
rect 35 28 37 30
rect 29 26 37 28
rect 29 23 31 26
rect 41 23 43 33
rect 9 10 11 15
rect 19 10 21 15
rect 29 10 31 15
rect 41 10 43 15
<< ndif >>
rect 2 27 9 29
rect 2 25 4 27
rect 6 25 9 27
rect 2 23 9 25
rect 4 15 9 23
rect 11 23 16 29
rect 11 19 19 23
rect 11 17 14 19
rect 16 17 19 19
rect 11 15 19 17
rect 21 21 29 23
rect 21 19 24 21
rect 26 19 29 21
rect 21 15 29 19
rect 31 15 41 23
rect 43 21 50 23
rect 43 19 46 21
rect 48 19 50 21
rect 43 17 50 19
rect 43 15 48 17
rect 33 11 39 15
rect 33 9 35 11
rect 37 9 39 11
rect 33 7 39 9
<< pdif >>
rect 13 71 20 73
rect 13 70 15 71
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 55 9 60
rect 2 53 4 55
rect 6 53 9 55
rect 2 51 9 53
rect 4 42 9 51
rect 11 69 15 70
rect 17 70 20 71
rect 17 69 22 70
rect 11 42 22 69
rect 24 42 29 70
rect 31 42 36 70
rect 38 63 43 70
rect 38 61 45 63
rect 38 59 41 61
rect 43 59 45 61
rect 38 57 45 59
rect 38 42 43 57
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 15 71
rect 17 69 58 71
rect -2 68 58 69
rect 2 62 14 63
rect 2 60 4 62
rect 6 60 14 62
rect 2 57 14 60
rect 2 55 6 57
rect 2 53 4 55
rect 2 27 6 53
rect 34 49 46 55
rect 26 38 30 47
rect 17 37 30 38
rect 17 35 21 37
rect 23 35 30 37
rect 17 34 30 35
rect 34 30 38 39
rect 42 38 46 49
rect 42 37 49 38
rect 42 35 45 37
rect 47 35 49 37
rect 42 34 49 35
rect 2 25 4 27
rect 2 17 6 25
rect 31 28 33 30
rect 35 28 47 30
rect 31 26 47 28
rect -2 11 58 12
rect -2 9 35 11
rect 37 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 15 11 29
rect 19 15 21 23
rect 29 15 31 23
rect 41 15 43 23
<< pmos >>
rect 9 42 11 70
rect 22 42 24 70
rect 29 42 31 70
rect 36 42 38 70
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 21 35 23 37
rect 45 35 47 37
rect 33 28 35 30
<< ndifct0 >>
rect 14 17 16 19
rect 24 19 26 21
rect 46 19 48 21
<< ndifct1 >>
rect 4 25 6 27
rect 35 9 37 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 41 59 43 61
<< pdifct1 >>
rect 4 60 6 62
rect 4 53 6 55
rect 15 69 17 71
<< alu0 >>
rect 18 61 45 62
rect 18 59 41 61
rect 43 59 45 61
rect 18 58 45 59
rect 6 51 7 57
rect 18 47 22 58
rect 10 43 22 47
rect 10 37 14 43
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 31 30 34 31
rect 6 23 7 29
rect 10 25 26 29
rect 22 22 26 25
rect 22 21 50 22
rect 13 19 17 21
rect 13 17 14 19
rect 16 17 17 19
rect 22 19 24 21
rect 26 19 46 21
rect 48 19 50 21
rect 22 18 50 19
rect 13 12 17 17
<< labels >>
rlabel polyct0 12 36 12 36 6 zn
rlabel alu0 36 20 36 20 6 zn
rlabel alu0 31 60 31 60 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 36 20 36 6 a
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 32 36 32 6 b
rlabel alu1 28 44 28 44 6 a
rlabel alu1 36 52 36 52 6 c
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 b
rlabel alu1 44 48 44 48 6 c
<< end >>
