magic
tech scmos
timestamp 1199202633
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 10 59 16 61
rect 10 57 12 59
rect 14 57 16 59
rect 10 55 16 57
rect 10 52 12 55
rect 20 52 22 57
rect 10 39 12 42
rect 20 39 22 42
rect 9 36 12 39
rect 16 37 23 39
rect 9 30 11 36
rect 16 35 19 37
rect 21 35 23 37
rect 16 33 23 35
rect 16 30 18 33
rect 9 8 11 13
rect 16 8 18 13
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 13 9 17
rect 11 13 16 30
rect 18 17 26 30
rect 18 15 21 17
rect 23 15 26 17
rect 18 13 26 15
<< pdif >>
rect 2 69 8 71
rect 2 67 4 69
rect 6 67 8 69
rect 2 52 8 67
rect 24 53 30 55
rect 24 52 26 53
rect 2 42 10 52
rect 12 46 20 52
rect 12 44 15 46
rect 17 44 20 46
rect 12 42 20 44
rect 22 51 26 52
rect 28 51 30 53
rect 22 42 30 51
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 69 34 79
rect -2 68 4 69
rect 6 68 34 69
rect 9 59 23 62
rect 9 57 12 59
rect 14 58 23 59
rect 14 57 15 58
rect 9 50 15 57
rect 2 44 15 46
rect 17 44 19 46
rect 2 42 19 44
rect 2 30 6 42
rect 17 37 23 38
rect 17 35 19 37
rect 21 35 23 37
rect 17 31 23 35
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 17 25 30 31
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 13 11 30
rect 16 13 18 30
<< pmos >>
rect 10 42 12 52
rect 20 42 22 52
<< polyct1 >>
rect 12 57 14 59
rect 19 35 21 37
<< ndifct0 >>
rect 21 15 23 17
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 67 6 68
rect 26 51 28 53
<< pdifct1 >>
rect 4 68 6 69
rect 15 44 17 46
<< alu0 >>
rect 2 67 4 68
rect 6 67 8 68
rect 2 66 8 67
rect 26 54 30 68
rect 24 53 30 54
rect 24 51 26 53
rect 28 51 30 53
rect 24 50 30 51
rect 13 46 19 47
rect 20 17 24 19
rect 20 15 21 17
rect 23 15 24 17
rect 20 12 24 15
<< labels >>
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 12 56 12 56 6 b
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 32 20 32 6 a
rlabel alu1 20 60 20 60 6 b
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 28 28 28 6 a
<< end >>
