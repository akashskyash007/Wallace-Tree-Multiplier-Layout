magic
tech scmos
timestamp 1199201796
<< ab >>
rect 0 0 88 80
<< nwell >>
rect -5 36 93 88
<< pwell >>
rect -5 -8 93 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 53 70 55 74
rect 63 70 65 74
rect 73 70 75 74
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 16 37 28 39
rect 20 35 24 37
rect 26 35 28 37
rect 20 33 28 35
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 9 27 15 29
rect 10 24 12 27
rect 20 24 22 33
rect 33 31 35 42
rect 43 39 45 42
rect 53 39 55 42
rect 63 39 65 42
rect 43 37 49 39
rect 43 35 45 37
rect 47 35 49 37
rect 43 33 49 35
rect 53 37 65 39
rect 73 39 75 42
rect 73 37 79 39
rect 53 35 55 37
rect 57 35 59 37
rect 53 33 59 35
rect 73 35 75 37
rect 77 35 79 37
rect 73 33 79 35
rect 33 29 39 31
rect 47 30 49 33
rect 54 30 56 33
rect 33 27 35 29
rect 37 27 39 29
rect 33 25 39 27
rect 10 9 12 14
rect 20 9 22 14
rect 47 8 49 13
rect 54 8 56 13
<< ndif >>
rect 2 14 10 24
rect 12 21 20 24
rect 12 19 15 21
rect 17 19 20 21
rect 12 14 20 19
rect 22 14 31 24
rect 42 23 47 30
rect 40 21 47 23
rect 40 19 42 21
rect 44 19 47 21
rect 40 17 47 19
rect 2 11 8 14
rect 2 9 4 11
rect 6 9 8 11
rect 24 11 31 14
rect 42 13 47 17
rect 49 13 54 30
rect 56 24 63 30
rect 56 22 59 24
rect 61 22 63 24
rect 56 17 63 22
rect 56 15 59 17
rect 61 15 63 17
rect 56 13 63 15
rect 24 9 26 11
rect 28 9 31 11
rect 2 7 8 9
rect 24 7 31 9
<< pdif >>
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 42 9 58
rect 11 42 16 70
rect 18 54 26 70
rect 18 52 21 54
rect 23 52 26 54
rect 18 47 26 52
rect 18 45 21 47
rect 23 45 26 47
rect 18 42 26 45
rect 28 42 33 70
rect 35 61 43 70
rect 35 59 38 61
rect 40 59 43 61
rect 35 54 43 59
rect 35 52 38 54
rect 40 52 43 54
rect 35 42 43 52
rect 45 68 53 70
rect 45 66 48 68
rect 50 66 53 68
rect 45 61 53 66
rect 45 59 48 61
rect 50 59 53 61
rect 45 42 53 59
rect 55 60 63 70
rect 55 58 58 60
rect 60 58 63 60
rect 55 53 63 58
rect 55 51 58 53
rect 60 51 63 53
rect 55 42 63 51
rect 65 68 73 70
rect 65 66 68 68
rect 70 66 73 68
rect 65 61 73 66
rect 65 59 68 61
rect 70 59 73 61
rect 65 42 73 59
rect 75 63 80 70
rect 75 61 82 63
rect 75 59 78 61
rect 80 59 82 61
rect 75 54 82 59
rect 75 52 78 54
rect 80 52 82 54
rect 75 50 82 52
rect 75 42 80 50
<< alu1 >>
rect -2 81 90 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 90 81
rect -2 68 90 79
rect 2 54 25 55
rect 2 52 21 54
rect 23 52 25 54
rect 2 51 25 52
rect 2 22 6 51
rect 18 50 25 51
rect 19 47 25 50
rect 10 31 14 47
rect 19 45 21 47
rect 23 45 25 47
rect 19 44 25 45
rect 33 38 39 46
rect 22 37 39 38
rect 22 35 24 37
rect 26 35 39 37
rect 22 34 39 35
rect 43 42 78 46
rect 43 37 49 42
rect 43 35 45 37
rect 47 35 49 37
rect 43 34 49 35
rect 53 37 70 38
rect 53 35 55 37
rect 57 35 70 37
rect 53 34 70 35
rect 10 29 11 31
rect 13 30 14 31
rect 13 29 39 30
rect 10 27 35 29
rect 37 27 39 29
rect 10 26 39 27
rect 2 21 47 22
rect 2 19 15 21
rect 17 19 42 21
rect 44 19 47 21
rect 2 18 47 19
rect 66 17 70 34
rect 74 37 78 42
rect 74 35 75 37
rect 77 35 78 37
rect 74 25 78 35
rect -2 11 90 12
rect -2 9 4 11
rect 6 9 26 11
rect 28 9 90 11
rect -2 1 90 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 90 1
rect -2 -2 90 -1
<< ptie >>
rect 0 1 88 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 88 1
rect 0 -3 88 -1
<< ntie >>
rect 0 81 88 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 88 81
rect 0 77 88 79
<< nmos >>
rect 10 14 12 24
rect 20 14 22 24
rect 47 13 49 30
rect 54 13 56 30
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 53 42 55 70
rect 63 42 65 70
rect 73 42 75 70
<< polyct1 >>
rect 24 35 26 37
rect 11 29 13 31
rect 45 35 47 37
rect 55 35 57 37
rect 75 35 77 37
rect 35 27 37 29
<< ndifct0 >>
rect 59 22 61 24
rect 59 15 61 17
<< ndifct1 >>
rect 15 19 17 21
rect 42 19 44 21
rect 4 9 6 11
rect 26 9 28 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
<< pdifct0 >>
rect 4 60 6 62
rect 38 59 40 61
rect 38 52 40 54
rect 48 66 50 68
rect 48 59 50 61
rect 58 58 60 60
rect 58 51 60 53
rect 68 66 70 68
rect 68 59 70 61
rect 78 59 80 61
rect 78 52 80 54
<< pdifct1 >>
rect 21 52 23 54
rect 21 45 23 47
<< alu0 >>
rect 46 66 48 68
rect 50 66 52 68
rect 2 62 41 63
rect 2 60 4 62
rect 6 61 41 62
rect 6 60 38 61
rect 2 59 38 60
rect 40 59 41 61
rect 6 50 18 51
rect 37 54 41 59
rect 46 61 52 66
rect 66 66 68 68
rect 70 66 72 68
rect 46 59 48 61
rect 50 59 52 61
rect 46 58 52 59
rect 57 60 61 62
rect 57 58 58 60
rect 60 58 61 60
rect 66 61 72 66
rect 66 59 68 61
rect 70 59 72 61
rect 66 58 72 59
rect 77 61 81 63
rect 77 59 78 61
rect 80 59 81 61
rect 57 54 61 58
rect 77 54 81 59
rect 37 52 38 54
rect 40 53 78 54
rect 40 52 58 53
rect 37 51 58 52
rect 60 52 78 53
rect 80 52 81 54
rect 60 51 81 52
rect 37 50 81 51
rect 58 24 62 26
rect 58 22 59 24
rect 61 22 62 24
rect 58 17 62 22
rect 58 15 59 17
rect 61 15 62 17
rect 58 12 62 15
<< labels >>
rlabel alu0 39 56 39 56 6 n1
rlabel alu0 21 61 21 61 6 n1
rlabel alu0 59 56 59 56 6 n1
rlabel pdifct0 59 52 59 52 6 n1
rlabel alu0 79 56 79 56 6 n1
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel polyct1 36 28 36 28 6 b
rlabel alu1 28 36 28 36 6 c
rlabel alu1 28 28 28 28 6 b
rlabel alu1 36 40 36 40 6 c
rlabel alu1 20 52 20 52 6 z
rlabel alu1 44 6 44 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 60 36 60 36 6 a1
rlabel alu1 52 44 52 44 6 a2
rlabel alu1 60 44 60 44 6 a2
rlabel alu1 44 74 44 74 6 vdd
rlabel alu1 68 24 68 24 6 a1
rlabel alu1 76 32 76 32 6 a2
rlabel alu1 68 44 68 44 6 a2
<< end >>
