magic
tech scmos
timestamp 1199469569
<< ab >>
rect 0 0 30 100
<< nwell >>
rect -2 48 32 104
<< pwell >>
rect -2 -4 32 48
<< poly >>
rect 15 73 17 78
rect 15 50 17 61
rect 15 48 23 50
rect 15 46 19 48
rect 21 46 23 48
rect 15 44 23 46
rect 15 23 17 44
rect 15 12 17 17
<< ndif >>
rect 7 21 15 23
rect 7 19 9 21
rect 11 19 15 21
rect 7 17 15 19
rect 17 21 26 23
rect 17 19 21 21
rect 23 19 26 21
rect 17 17 26 19
<< pdif >>
rect 10 67 15 73
rect 7 65 15 67
rect 7 63 9 65
rect 11 63 15 65
rect 7 61 15 63
rect 17 71 26 73
rect 17 69 21 71
rect 23 69 26 71
rect 17 61 26 69
<< alu1 >>
rect -2 95 32 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 32 95
rect -2 88 32 93
rect 8 65 12 73
rect 20 71 24 88
rect 20 69 21 71
rect 23 69 24 71
rect 20 67 24 69
rect 8 63 9 65
rect 11 63 12 65
rect 8 32 12 63
rect 18 48 22 63
rect 18 46 19 48
rect 21 46 22 48
rect 18 37 22 46
rect 8 27 23 32
rect 8 21 12 27
rect 8 19 9 21
rect 11 19 12 21
rect 8 17 12 19
rect 20 21 24 23
rect 20 19 21 21
rect 23 19 24 21
rect 20 12 24 19
rect -2 7 32 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 32 7
rect -2 0 32 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 15 17 17 23
<< pmos >>
rect 15 61 17 73
<< polyct1 >>
rect 19 46 21 48
<< ndifct1 >>
rect 9 19 11 21
rect 21 19 23 21
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 9 63 11 65
rect 21 69 23 71
<< labels >>
rlabel alu1 10 45 10 45 6 z
rlabel alu1 15 6 15 6 6 vss
rlabel alu1 20 30 20 30 6 z
rlabel alu1 20 50 20 50 6 a
rlabel alu1 15 94 15 94 6 vdd
<< end >>
