magic
tech scmos
timestamp 1199203308
<< ab >>
rect 0 0 88 72
<< nwell >>
rect -5 32 93 77
<< pwell >>
rect -5 -5 93 32
<< poly >>
rect 9 66 11 70
rect 21 66 23 70
rect 28 66 30 70
rect 35 66 37 70
rect 42 66 44 70
rect 52 66 54 70
rect 59 66 61 70
rect 66 66 68 70
rect 73 66 75 70
rect 21 39 23 42
rect 9 29 11 38
rect 18 37 24 39
rect 18 35 20 37
rect 22 35 24 37
rect 18 33 24 35
rect 9 27 15 29
rect 9 25 11 27
rect 13 25 15 27
rect 9 23 15 25
rect 9 20 11 23
rect 21 18 23 33
rect 28 27 30 42
rect 35 33 37 42
rect 42 39 44 42
rect 52 39 54 42
rect 42 37 55 39
rect 49 33 55 37
rect 35 31 41 33
rect 39 27 41 31
rect 49 31 51 33
rect 53 31 55 33
rect 49 29 55 31
rect 27 25 33 27
rect 27 23 29 25
rect 31 23 33 25
rect 27 21 33 23
rect 39 25 45 27
rect 39 23 41 25
rect 43 23 45 25
rect 39 21 45 23
rect 31 18 33 21
rect 43 18 45 21
rect 53 18 55 29
rect 59 23 61 42
rect 66 33 68 42
rect 73 39 75 42
rect 73 37 82 39
rect 76 35 78 37
rect 80 35 82 37
rect 76 33 82 35
rect 65 31 71 33
rect 65 29 67 31
rect 69 29 71 31
rect 65 27 71 29
rect 59 21 67 23
rect 65 19 67 21
rect 65 17 71 19
rect 65 15 67 17
rect 69 15 71 17
rect 65 13 71 15
rect 9 2 11 6
rect 21 6 23 11
rect 31 6 33 11
rect 43 6 45 11
rect 53 6 55 11
<< ndif >>
rect 2 17 9 20
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 6 9 13
rect 11 18 19 20
rect 11 11 21 18
rect 23 16 31 18
rect 23 14 26 16
rect 28 14 31 16
rect 23 11 31 14
rect 33 11 43 18
rect 45 16 53 18
rect 45 14 48 16
rect 50 14 53 16
rect 45 11 53 14
rect 55 11 63 18
rect 11 7 19 11
rect 11 6 15 7
rect 13 5 15 6
rect 17 5 19 7
rect 35 7 41 11
rect 13 3 19 5
rect 35 5 37 7
rect 39 5 41 7
rect 57 7 63 11
rect 35 3 41 5
rect 57 5 59 7
rect 61 5 63 7
rect 57 3 63 5
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 21 66
rect 11 62 15 64
rect 17 62 21 64
rect 11 42 21 62
rect 23 42 28 66
rect 30 42 35 66
rect 37 42 42 66
rect 44 57 52 66
rect 44 55 47 57
rect 49 55 52 57
rect 44 42 52 55
rect 54 42 59 66
rect 61 42 66 66
rect 68 42 73 66
rect 75 64 82 66
rect 75 62 78 64
rect 80 62 82 64
rect 75 57 82 62
rect 75 55 78 57
rect 80 55 82 57
rect 75 42 82 55
rect 11 38 16 42
<< alu1 >>
rect -2 64 90 72
rect 2 49 6 59
rect 2 47 4 49
rect 2 42 6 47
rect 2 40 4 42
rect 2 19 6 40
rect 58 50 62 59
rect 18 46 79 50
rect 18 37 23 46
rect 18 35 20 37
rect 22 35 23 37
rect 18 33 23 35
rect 29 38 70 42
rect 29 27 33 38
rect 41 33 55 34
rect 41 31 51 33
rect 53 31 55 33
rect 41 30 55 31
rect 66 31 70 38
rect 66 29 67 31
rect 69 29 70 31
rect 74 37 79 46
rect 74 35 78 37
rect 74 29 79 35
rect 66 27 70 29
rect 2 17 14 19
rect 2 15 4 17
rect 6 15 14 17
rect 2 13 14 15
rect 26 25 33 27
rect 26 23 29 25
rect 31 23 33 25
rect 26 21 33 23
rect 39 25 61 26
rect 39 23 41 25
rect 43 23 61 25
rect 39 22 61 23
rect 57 18 61 22
rect 57 17 71 18
rect 57 15 67 17
rect 69 15 71 17
rect 57 14 71 15
rect -2 7 90 8
rect -2 5 15 7
rect 17 5 37 7
rect 39 5 59 7
rect 61 5 69 7
rect 71 5 77 7
rect 79 5 90 7
rect -2 0 90 5
<< ptie >>
rect 67 7 81 9
rect 67 5 69 7
rect 71 5 77 7
rect 79 5 81 7
rect 67 3 81 5
<< nmos >>
rect 9 6 11 20
rect 21 11 23 18
rect 31 11 33 18
rect 43 11 45 18
rect 53 11 55 18
<< pmos >>
rect 9 38 11 66
rect 21 42 23 66
rect 28 42 30 66
rect 35 42 37 66
rect 42 42 44 66
rect 52 42 54 66
rect 59 42 61 66
rect 66 42 68 66
rect 73 42 75 66
<< polyct0 >>
rect 11 25 13 27
rect 79 35 80 37
<< polyct1 >>
rect 20 35 22 37
rect 51 31 53 33
rect 29 23 31 25
rect 41 23 43 25
rect 78 35 79 37
rect 67 29 69 31
rect 67 15 69 17
<< ndifct0 >>
rect 26 14 28 16
rect 48 14 50 16
<< ndifct1 >>
rect 4 15 6 17
rect 15 5 17 7
rect 37 5 39 7
rect 59 5 61 7
<< ptiect1 >>
rect 69 5 71 7
rect 77 5 79 7
<< pdifct0 >>
rect 15 62 17 64
rect 47 55 49 57
rect 78 62 80 64
rect 78 55 80 57
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
<< alu0 >>
rect 13 62 15 64
rect 17 62 19 64
rect 13 61 19 62
rect 76 62 78 64
rect 80 62 82 64
rect 10 57 51 58
rect 10 55 47 57
rect 49 55 51 57
rect 10 54 51 55
rect 6 38 7 51
rect 10 27 14 54
rect 76 57 82 62
rect 76 55 78 57
rect 80 55 82 57
rect 76 54 82 55
rect 79 37 82 39
rect 80 35 82 37
rect 79 33 82 35
rect 10 25 11 27
rect 13 25 22 27
rect 10 23 22 25
rect 18 17 22 23
rect 18 16 52 17
rect 18 14 26 16
rect 28 14 48 16
rect 50 14 52 16
rect 18 13 52 14
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 35 15 35 15 6 zn
rlabel alu0 30 56 30 56 6 zn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 28 24 28 24 6 b
rlabel alu1 20 40 20 40 6 a
rlabel alu1 28 48 28 48 6 a
rlabel alu1 44 4 44 4 6 vss
rlabel alu1 44 24 44 24 6 c
rlabel alu1 44 32 44 32 6 d
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 48 36 48 6 a
rlabel alu1 44 48 44 48 6 a
rlabel alu1 44 68 44 68 6 vdd
rlabel alu1 60 16 60 16 6 c
rlabel polyct1 68 16 68 16 6 c
rlabel alu1 52 24 52 24 6 c
rlabel alu1 68 32 68 32 6 b
rlabel polyct1 52 32 52 32 6 d
rlabel alu1 52 40 52 40 6 b
rlabel alu1 60 40 60 40 6 b
rlabel alu1 52 48 52 48 6 a
rlabel alu1 60 52 60 52 6 a
rlabel alu1 68 48 68 48 6 a
rlabel alu1 76 40 76 40 6 a
<< end >>
