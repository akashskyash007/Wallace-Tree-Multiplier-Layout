magic
tech scmos
timestamp 1199973039
<< ab >>
rect 0 0 32 88
<< nwell >>
rect -5 40 37 97
<< pwell >>
rect -5 -9 37 40
<< poly >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 21 74 23 77
rect 9 43 11 46
rect 21 43 23 46
rect 2 41 14 43
rect 2 39 7 41
rect 9 39 14 41
rect 2 37 14 39
rect 18 41 30 43
rect 18 39 23 41
rect 25 39 30 41
rect 18 37 30 39
rect 9 34 11 37
rect 21 34 23 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 21 5 30 11
<< ndif >>
rect 2 25 9 34
rect 2 23 4 25
rect 6 23 9 25
rect 2 18 9 23
rect 2 16 4 18
rect 6 16 9 18
rect 2 14 9 16
rect 11 32 21 34
rect 11 30 15 32
rect 17 30 21 32
rect 11 24 21 30
rect 11 22 15 24
rect 17 22 21 24
rect 11 14 21 22
rect 23 25 30 34
rect 23 23 26 25
rect 28 23 30 25
rect 23 18 30 23
rect 23 16 26 18
rect 28 16 30 18
rect 23 14 30 16
rect 13 2 19 14
<< pdif >>
rect 13 74 19 86
rect 2 72 9 74
rect 2 70 4 72
rect 6 70 9 72
rect 2 46 9 70
rect 11 50 21 74
rect 11 48 15 50
rect 17 48 21 50
rect 11 46 21 48
rect 23 72 30 74
rect 23 70 26 72
rect 28 70 30 72
rect 23 46 30 70
<< alu1 >>
rect -2 89 34 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 34 89
rect -2 86 34 87
rect 3 81 7 86
rect 3 79 4 81
rect 6 79 7 81
rect 3 72 7 79
rect 3 70 4 72
rect 6 70 7 72
rect 3 68 7 70
rect 25 81 29 86
rect 25 79 26 81
rect 28 79 29 81
rect 25 72 29 79
rect 25 70 26 72
rect 28 70 29 72
rect 25 68 29 70
rect 6 59 26 63
rect 6 41 10 59
rect 6 39 7 41
rect 9 39 10 41
rect 6 33 10 39
rect 14 50 18 55
rect 14 48 15 50
rect 17 48 18 50
rect 14 32 18 48
rect 22 41 26 59
rect 22 39 23 41
rect 25 39 26 41
rect 22 33 26 39
rect 14 30 15 32
rect 17 30 18 32
rect 3 25 7 27
rect 3 23 4 25
rect 6 23 7 25
rect 3 18 7 23
rect 3 16 4 18
rect 6 16 7 18
rect 14 24 18 30
rect 14 22 15 24
rect 17 22 18 24
rect 14 17 18 22
rect 25 25 29 27
rect 25 23 26 25
rect 28 23 29 25
rect 25 18 29 23
rect 3 9 7 16
rect 3 7 4 9
rect 6 7 7 9
rect 3 2 7 7
rect 25 16 26 18
rect 28 16 29 18
rect 25 9 29 16
rect 25 7 26 9
rect 28 7 29 9
rect 25 2 29 7
rect -2 1 34 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< alu2 >>
rect -2 89 34 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 34 89
rect -2 81 34 87
rect -2 79 4 81
rect 6 79 26 81
rect 28 79 34 81
rect -2 76 34 79
rect -2 9 34 12
rect -2 7 4 9
rect 6 7 26 9
rect 28 7 34 9
rect -2 1 34 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 32 3
rect 25 -1 27 1
rect 29 -1 32 1
rect 25 -3 32 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 32 91
rect 25 87 27 89
rect 29 87 32 89
rect 25 85 32 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
<< polyct1 >>
rect 7 39 9 41
rect 23 39 25 41
<< ndifct1 >>
rect 4 23 6 25
rect 4 16 6 18
rect 15 30 17 32
rect 15 22 17 24
rect 26 23 28 25
rect 26 16 28 18
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
<< pdifct1 >>
rect 4 70 6 72
rect 15 48 17 50
rect 26 70 28 72
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 4 79 6 81
rect 26 79 28 81
rect 4 7 6 9
rect 26 7 28 9
rect 7 -1 9 1
rect 23 -1 25 1
<< labels >>
rlabel alu1 8 48 8 48 6 a
rlabel alu1 16 36 16 36 6 z
rlabel alu1 24 48 24 48 6 a
rlabel alu2 16 6 16 6 6 vss
rlabel alu2 16 6 16 6 6 vss
rlabel alu2 16 82 16 82 6 vdd
<< end >>
