magic
tech scmos
timestamp 1199203476
<< ab >>
rect 0 0 104 72
<< nwell >>
rect -5 32 109 77
<< pwell >>
rect -5 -5 109 32
<< poly >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 53 66 55 70
rect 63 64 65 69
rect 73 64 75 69
rect 83 57 85 62
rect 93 57 95 61
rect 9 19 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 16 33 28 35
rect 16 31 24 33
rect 26 31 28 33
rect 16 29 28 31
rect 23 26 25 29
rect 33 26 35 38
rect 43 35 45 46
rect 53 43 55 46
rect 63 43 65 46
rect 73 43 75 46
rect 53 41 65 43
rect 43 33 57 35
rect 43 31 51 33
rect 53 31 57 33
rect 43 29 57 31
rect 63 31 65 41
rect 69 41 75 43
rect 69 39 71 41
rect 73 39 75 41
rect 69 37 75 39
rect 83 31 85 38
rect 93 35 95 38
rect 93 33 102 35
rect 93 31 98 33
rect 100 31 102 33
rect 63 29 102 31
rect 43 26 45 29
rect 55 26 57 29
rect 78 26 80 29
rect 5 17 11 19
rect 5 15 7 17
rect 9 15 11 17
rect 5 13 11 15
rect 55 15 57 20
rect 63 16 69 18
rect 43 8 45 13
rect 23 2 25 7
rect 33 4 35 7
rect 63 14 65 16
rect 67 14 69 16
rect 63 12 69 14
rect 63 4 65 12
rect 33 2 65 4
rect 78 2 80 7
<< ndif >>
rect 18 19 23 26
rect 16 17 23 19
rect 16 15 18 17
rect 20 15 23 17
rect 16 13 23 15
rect 18 7 23 13
rect 25 24 33 26
rect 25 22 28 24
rect 30 22 33 24
rect 25 7 33 22
rect 35 24 43 26
rect 35 22 38 24
rect 40 22 43 24
rect 35 13 43 22
rect 45 20 55 26
rect 57 24 64 26
rect 57 22 60 24
rect 62 22 64 24
rect 57 20 64 22
rect 71 24 78 26
rect 71 22 73 24
rect 75 22 78 24
rect 45 13 53 20
rect 35 7 40 13
rect 47 10 53 13
rect 47 8 49 10
rect 51 8 53 10
rect 47 6 53 8
rect 71 17 78 22
rect 71 15 73 17
rect 75 15 78 17
rect 71 13 78 15
rect 73 7 78 13
rect 80 18 88 26
rect 80 16 83 18
rect 85 16 88 18
rect 80 11 88 16
rect 80 9 83 11
rect 85 9 88 11
rect 80 7 88 9
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 38 16 66
rect 18 57 26 66
rect 18 55 21 57
rect 23 55 26 57
rect 18 42 26 55
rect 18 40 21 42
rect 23 40 26 42
rect 18 38 26 40
rect 28 38 33 66
rect 35 64 43 66
rect 35 62 38 64
rect 40 62 43 64
rect 35 46 43 62
rect 45 50 53 66
rect 45 48 48 50
rect 50 48 53 50
rect 45 46 53 48
rect 55 64 60 66
rect 55 57 63 64
rect 55 55 58 57
rect 60 55 63 57
rect 55 46 63 55
rect 65 57 73 64
rect 65 55 68 57
rect 70 55 73 57
rect 65 50 73 55
rect 65 48 68 50
rect 70 48 73 50
rect 65 46 73 48
rect 75 57 81 64
rect 75 55 83 57
rect 75 53 78 55
rect 80 53 83 55
rect 75 46 83 53
rect 35 38 41 46
rect 77 38 83 46
rect 85 49 93 57
rect 85 47 88 49
rect 90 47 93 49
rect 85 42 93 47
rect 85 40 88 42
rect 90 40 93 42
rect 85 38 93 40
rect 95 55 102 57
rect 95 53 98 55
rect 100 53 102 55
rect 95 48 102 53
rect 95 46 98 48
rect 100 46 102 48
rect 95 38 102 46
<< alu1 >>
rect -2 67 106 72
rect -2 65 89 67
rect 91 65 97 67
rect 99 65 106 67
rect -2 64 106 65
rect 18 57 63 58
rect 18 55 21 57
rect 23 55 58 57
rect 60 55 63 57
rect 18 54 63 55
rect 18 44 22 54
rect 18 43 24 44
rect 10 42 24 43
rect 10 40 21 42
rect 23 40 24 42
rect 10 38 24 40
rect 10 26 14 38
rect 49 41 75 42
rect 49 39 71 41
rect 73 39 75 41
rect 49 38 75 39
rect 49 33 55 38
rect 49 31 51 33
rect 53 31 55 33
rect 49 30 55 31
rect 97 33 102 35
rect 97 31 98 33
rect 100 31 102 33
rect 10 24 32 26
rect 10 22 28 24
rect 30 22 32 24
rect 26 21 32 22
rect 97 19 102 31
rect 90 13 102 19
rect -2 7 106 8
rect -2 5 5 7
rect 7 5 97 7
rect 99 5 106 7
rect -2 0 106 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 95 7 101 24
rect 95 5 97 7
rect 99 5 101 7
rect 95 3 101 5
<< ntie >>
rect 87 67 101 69
rect 87 65 89 67
rect 91 65 97 67
rect 99 65 101 67
rect 87 63 101 65
<< nmos >>
rect 23 7 25 26
rect 33 7 35 26
rect 43 13 45 26
rect 55 20 57 26
rect 78 7 80 26
<< pmos >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 46 45 66
rect 53 46 55 66
rect 63 46 65 64
rect 73 46 75 64
rect 83 38 85 57
rect 93 38 95 57
<< polyct0 >>
rect 24 31 26 33
rect 7 15 9 17
rect 65 14 67 16
<< polyct1 >>
rect 51 31 53 33
rect 71 39 73 41
rect 98 31 100 33
<< ndifct0 >>
rect 18 15 20 17
rect 38 22 40 24
rect 60 22 62 24
rect 73 22 75 24
rect 49 8 51 10
rect 73 15 75 17
rect 83 16 85 18
rect 83 9 85 11
<< ndifct1 >>
rect 28 22 30 24
<< ntiect1 >>
rect 89 65 91 67
rect 97 65 99 67
<< ptiect1 >>
rect 5 5 7 7
rect 97 5 99 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 38 62 40 64
rect 48 48 50 50
rect 68 55 70 57
rect 68 48 70 50
rect 78 53 80 55
rect 88 47 90 49
rect 88 40 90 42
rect 98 53 100 55
rect 98 46 100 48
<< pdifct1 >>
rect 21 55 23 57
rect 21 40 23 42
rect 58 55 60 57
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 36 62 38 64
rect 40 62 42 64
rect 36 61 42 62
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 67 57 71 59
rect 67 55 68 57
rect 70 55 71 57
rect 46 50 52 51
rect 67 50 71 55
rect 77 55 81 64
rect 77 53 78 55
rect 80 53 81 55
rect 77 51 81 53
rect 97 55 101 64
rect 97 53 98 55
rect 100 53 101 55
rect 36 48 48 50
rect 50 48 68 50
rect 70 48 71 50
rect 36 46 71 48
rect 87 49 91 51
rect 87 47 88 49
rect 90 47 91 49
rect 36 34 40 46
rect 87 42 91 47
rect 97 48 101 53
rect 97 46 98 48
rect 100 46 101 48
rect 97 44 101 46
rect 22 33 40 34
rect 22 31 24 33
rect 26 31 40 33
rect 22 30 40 31
rect 87 40 88 42
rect 90 40 91 42
rect 87 34 91 40
rect 72 30 91 34
rect 36 26 40 30
rect 36 24 64 26
rect 36 22 38 24
rect 40 22 60 24
rect 62 22 64 24
rect 36 21 42 22
rect 58 21 64 22
rect 72 24 76 30
rect 72 22 73 24
rect 75 22 76 24
rect 72 18 76 22
rect 5 17 76 18
rect 5 15 7 17
rect 9 15 18 17
rect 20 16 73 17
rect 20 15 65 16
rect 5 14 65 15
rect 67 15 73 16
rect 75 15 76 17
rect 67 14 76 15
rect 63 13 76 14
rect 82 18 86 20
rect 82 16 83 18
rect 85 16 86 18
rect 82 11 86 16
rect 47 10 53 11
rect 47 8 49 10
rect 51 8 53 10
rect 82 9 83 11
rect 85 9 86 11
rect 82 8 86 9
<< labels >>
rlabel alu0 31 32 31 32 6 an
rlabel alu0 50 24 50 24 6 an
rlabel alu0 53 48 53 48 6 an
rlabel alu0 69 52 69 52 6 an
rlabel alu0 40 16 40 16 6 bn
rlabel ndifct0 74 23 74 23 6 bn
rlabel alu0 89 40 89 40 6 bn
rlabel alu1 20 24 20 24 6 z
rlabel alu1 12 36 12 36 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 52 4 52 4 6 vss
rlabel alu1 68 40 68 40 6 a
rlabel alu1 60 40 60 40 6 a
rlabel alu1 52 36 52 36 6 a
rlabel alu1 60 56 60 56 6 z
rlabel alu1 52 56 52 56 6 z
rlabel alu1 52 68 52 68 6 vdd
rlabel alu1 92 16 92 16 6 b
rlabel alu1 100 24 100 24 6 b
<< end >>
