magic
tech scmos
timestamp 1199202805
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 37 70 39 74
rect 49 70 51 74
rect 15 63 17 67
rect 25 63 27 67
rect 15 46 17 49
rect 25 46 27 49
rect 15 44 27 46
rect 17 42 19 44
rect 21 42 23 44
rect 17 40 23 42
rect 7 37 13 39
rect 7 35 9 37
rect 11 35 13 37
rect 7 33 14 35
rect 12 30 14 33
rect 19 30 21 40
rect 37 39 39 42
rect 33 37 39 39
rect 33 35 35 37
rect 37 35 39 37
rect 49 39 51 42
rect 49 37 55 39
rect 49 35 51 37
rect 53 35 55 37
rect 26 33 39 35
rect 26 30 28 33
rect 36 30 38 33
rect 43 30 45 35
rect 49 33 55 35
rect 50 30 52 33
rect 12 11 14 16
rect 19 8 21 16
rect 26 12 28 16
rect 36 12 38 16
rect 43 8 45 16
rect 50 11 52 16
rect 19 6 45 8
<< ndif >>
rect 2 27 12 30
rect 2 25 4 27
rect 6 25 12 27
rect 2 20 12 25
rect 2 18 4 20
rect 6 18 12 20
rect 2 16 12 18
rect 14 16 19 30
rect 21 16 26 30
rect 28 28 36 30
rect 28 26 31 28
rect 33 26 36 28
rect 28 16 36 26
rect 38 16 43 30
rect 45 16 50 30
rect 52 27 60 30
rect 52 25 55 27
rect 57 25 60 27
rect 52 20 60 25
rect 52 18 55 20
rect 57 18 60 20
rect 52 16 60 18
<< pdif >>
rect 29 68 37 70
rect 29 66 31 68
rect 33 66 37 68
rect 29 63 37 66
rect 6 61 15 63
rect 6 59 9 61
rect 11 59 15 61
rect 6 49 15 59
rect 17 61 25 63
rect 17 59 20 61
rect 22 59 25 61
rect 17 53 25 59
rect 17 51 20 53
rect 22 51 25 53
rect 17 49 25 51
rect 27 61 37 63
rect 27 59 31 61
rect 33 59 37 61
rect 27 49 37 59
rect 29 42 37 49
rect 39 61 49 70
rect 39 59 43 61
rect 45 59 49 61
rect 39 53 49 59
rect 39 51 43 53
rect 45 51 49 53
rect 39 42 49 51
rect 51 68 59 70
rect 51 66 54 68
rect 56 66 59 68
rect 51 61 59 66
rect 51 59 54 61
rect 56 59 59 61
rect 51 42 59 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 18 61 23 63
rect 18 59 20 61
rect 22 59 23 61
rect 9 46 14 55
rect 18 54 23 59
rect 41 61 47 62
rect 41 59 43 61
rect 45 59 47 61
rect 41 54 47 59
rect 18 53 47 54
rect 18 51 20 53
rect 22 51 43 53
rect 45 51 47 53
rect 18 50 47 51
rect 9 44 22 46
rect 9 42 19 44
rect 21 42 22 44
rect 7 37 14 38
rect 7 35 9 37
rect 11 35 14 37
rect 7 34 14 35
rect 10 22 14 34
rect 18 33 22 42
rect 26 26 30 50
rect 34 42 47 46
rect 34 37 38 42
rect 34 35 35 37
rect 37 35 38 37
rect 34 33 38 35
rect 42 37 55 38
rect 42 35 51 37
rect 53 35 55 37
rect 42 34 55 35
rect 42 22 46 34
rect 10 18 46 22
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 12 16 14 30
rect 19 16 21 30
rect 26 16 28 30
rect 36 16 38 30
rect 43 16 45 30
rect 50 16 52 30
<< pmos >>
rect 15 49 17 63
rect 25 49 27 63
rect 37 42 39 70
rect 49 42 51 70
<< polyct1 >>
rect 19 42 21 44
rect 9 35 11 37
rect 35 35 37 37
rect 51 35 53 37
<< ndifct0 >>
rect 4 25 6 27
rect 4 18 6 20
rect 31 26 33 28
rect 55 25 57 27
rect 55 18 57 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 31 66 33 68
rect 9 59 11 61
rect 31 59 33 61
rect 54 66 56 68
rect 54 59 56 61
<< pdifct1 >>
rect 20 59 22 61
rect 20 51 22 53
rect 43 59 45 61
rect 43 51 45 53
<< alu0 >>
rect 7 61 13 68
rect 29 66 31 68
rect 33 66 35 68
rect 7 59 9 61
rect 11 59 13 61
rect 7 58 13 59
rect 29 61 35 66
rect 52 66 54 68
rect 56 66 58 68
rect 29 59 31 61
rect 33 59 35 61
rect 29 58 35 59
rect 52 61 58 66
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
rect 3 27 7 29
rect 3 25 4 27
rect 6 25 7 27
rect 3 20 7 25
rect 3 18 4 20
rect 6 18 7 20
rect 30 28 35 29
rect 30 26 31 28
rect 33 26 35 28
rect 26 25 35 26
rect 54 27 58 29
rect 54 25 55 27
rect 57 25 58 27
rect 54 20 58 25
rect 54 18 55 20
rect 57 18 58 20
rect 3 12 7 18
rect 54 12 58 18
<< labels >>
rlabel alu1 12 28 12 28 6 a
rlabel alu1 12 48 12 48 6 b
rlabel alu1 20 20 20 20 6 a
rlabel alu1 28 20 28 20 6 a
rlabel alu1 20 36 20 36 6 b
rlabel alu1 28 44 28 44 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 20 36 20 6 a
rlabel polyct1 36 36 36 36 6 c
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 44 44 44 6 c
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel polyct1 52 36 52 36 6 a
<< end >>
