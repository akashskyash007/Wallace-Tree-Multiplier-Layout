magic
tech scmos
timestamp 1199201915
<< ab >>
rect 0 0 144 72
<< nwell >>
rect -5 32 149 77
<< pwell >>
rect -5 -5 149 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 99 66 101 70
rect 109 66 111 70
rect 119 66 121 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 33 31 35
rect 9 31 11 33
rect 13 31 21 33
rect 9 29 21 31
rect 19 23 21 29
rect 29 23 31 33
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 39 33 61 35
rect 39 31 45 33
rect 47 31 57 33
rect 59 31 61 33
rect 39 29 61 31
rect 39 26 41 29
rect 49 26 51 29
rect 59 26 61 29
rect 69 35 71 38
rect 79 35 81 38
rect 89 35 91 38
rect 69 33 91 35
rect 69 31 77 33
rect 79 31 85 33
rect 87 31 91 33
rect 69 29 91 31
rect 69 26 71 29
rect 79 26 81 29
rect 89 26 91 29
rect 99 35 101 38
rect 109 35 111 38
rect 119 35 121 38
rect 99 33 121 35
rect 99 26 101 33
rect 108 31 110 33
rect 112 31 117 33
rect 119 31 121 33
rect 108 29 121 31
rect 109 26 111 29
rect 119 26 121 29
rect 19 7 21 12
rect 29 7 31 12
rect 39 3 41 8
rect 49 3 51 8
rect 59 3 61 8
rect 69 3 71 8
rect 79 3 81 8
rect 89 3 91 8
rect 99 3 101 8
rect 109 3 111 8
rect 119 3 121 8
<< ndif >>
rect 34 23 39 26
rect 12 21 19 23
rect 12 19 14 21
rect 16 19 19 21
rect 12 17 19 19
rect 14 12 19 17
rect 21 16 29 23
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 31 21 39 23
rect 31 19 34 21
rect 36 19 39 21
rect 31 12 39 19
rect 34 8 39 12
rect 41 16 49 26
rect 41 14 44 16
rect 46 14 49 16
rect 41 8 49 14
rect 51 24 59 26
rect 51 22 54 24
rect 56 22 59 24
rect 51 8 59 22
rect 61 23 69 26
rect 61 21 64 23
rect 66 21 69 23
rect 61 16 69 21
rect 61 14 64 16
rect 66 14 69 16
rect 61 8 69 14
rect 71 24 79 26
rect 71 22 74 24
rect 76 22 79 24
rect 71 8 79 22
rect 81 16 89 26
rect 81 14 84 16
rect 86 14 89 16
rect 81 8 89 14
rect 91 24 99 26
rect 91 22 94 24
rect 96 22 99 24
rect 91 17 99 22
rect 91 15 94 17
rect 96 15 99 17
rect 91 8 99 15
rect 101 12 109 26
rect 101 10 104 12
rect 106 10 109 12
rect 101 8 109 10
rect 111 24 119 26
rect 111 22 114 24
rect 116 22 119 24
rect 111 17 119 22
rect 111 15 114 17
rect 116 15 119 17
rect 111 8 119 15
rect 121 20 128 26
rect 121 18 124 20
rect 126 18 128 20
rect 121 12 128 18
rect 121 10 124 12
rect 126 10 128 12
rect 121 8 128 10
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 49 29 66
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 50 39 55
rect 31 48 34 50
rect 36 48 39 50
rect 31 38 39 48
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 38 49 55
rect 51 49 59 66
rect 51 47 54 49
rect 56 47 59 49
rect 51 42 59 47
rect 51 40 54 42
rect 56 40 59 42
rect 51 38 59 40
rect 61 64 69 66
rect 61 62 64 64
rect 66 62 69 64
rect 61 57 69 62
rect 61 55 64 57
rect 66 55 69 57
rect 61 38 69 55
rect 71 49 79 66
rect 71 47 74 49
rect 76 47 79 49
rect 71 42 79 47
rect 71 40 74 42
rect 76 40 79 42
rect 71 38 79 40
rect 81 64 89 66
rect 81 62 84 64
rect 86 62 89 64
rect 81 57 89 62
rect 81 55 84 57
rect 86 55 89 57
rect 81 38 89 55
rect 91 49 99 66
rect 91 47 94 49
rect 96 47 99 49
rect 91 42 99 47
rect 91 40 94 42
rect 96 40 99 42
rect 91 38 99 40
rect 101 64 109 66
rect 101 62 104 64
rect 106 62 109 64
rect 101 57 109 62
rect 101 55 104 57
rect 106 55 109 57
rect 101 38 109 55
rect 111 57 119 66
rect 111 55 114 57
rect 116 55 119 57
rect 111 50 119 55
rect 111 48 114 50
rect 116 48 119 50
rect 111 38 119 48
rect 121 64 128 66
rect 121 62 124 64
rect 126 62 128 64
rect 121 57 128 62
rect 121 55 124 57
rect 126 55 128 57
rect 121 38 128 55
<< alu1 >>
rect -2 67 146 72
rect -2 65 134 67
rect 136 65 146 67
rect -2 64 146 65
rect 2 49 7 59
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 2 40 4 42
rect 6 40 24 42
rect 26 40 30 42
rect 2 38 30 40
rect 2 33 15 34
rect 2 31 11 33
rect 13 31 15 33
rect 2 30 15 31
rect 2 13 6 30
rect 26 26 30 38
rect 41 34 47 42
rect 81 34 87 42
rect 122 34 127 51
rect 41 33 63 34
rect 41 31 45 33
rect 47 31 57 33
rect 59 31 63 33
rect 41 30 63 31
rect 73 33 95 34
rect 73 31 77 33
rect 79 31 85 33
rect 87 31 95 33
rect 73 30 95 31
rect 105 33 127 34
rect 105 31 110 33
rect 112 31 117 33
rect 119 31 127 33
rect 105 30 127 31
rect 13 24 58 26
rect 13 22 54 24
rect 56 22 58 24
rect 13 21 17 22
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect 33 21 58 22
rect 33 19 34 21
rect 36 19 38 21
rect 33 13 38 19
rect -2 7 146 8
rect -2 5 5 7
rect 7 5 134 7
rect 136 5 146 7
rect -2 0 146 5
<< ptie >>
rect 3 7 9 13
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 132 7 138 24
rect 132 5 134 7
rect 136 5 138 7
rect 132 3 138 5
<< ntie >>
rect 132 67 138 69
rect 132 65 134 67
rect 136 65 138 67
rect 132 40 138 65
<< nmos >>
rect 19 12 21 23
rect 29 12 31 23
rect 39 8 41 26
rect 49 8 51 26
rect 59 8 61 26
rect 69 8 71 26
rect 79 8 81 26
rect 89 8 91 26
rect 99 8 101 26
rect 109 8 111 26
rect 119 8 121 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 69 38 71 66
rect 79 38 81 66
rect 89 38 91 66
rect 99 38 101 66
rect 109 38 111 66
rect 119 38 121 66
<< polyct1 >>
rect 11 31 13 33
rect 45 31 47 33
rect 57 31 59 33
rect 77 31 79 33
rect 85 31 87 33
rect 110 31 112 33
rect 117 31 119 33
<< ndifct0 >>
rect 24 14 26 16
rect 44 14 46 16
rect 64 21 66 23
rect 64 14 66 16
rect 74 22 76 24
rect 84 14 86 16
rect 94 22 96 24
rect 94 15 96 17
rect 104 10 106 12
rect 114 22 116 24
rect 114 15 116 17
rect 124 18 126 20
rect 124 10 126 12
<< ndifct1 >>
rect 14 19 16 21
rect 34 19 36 21
rect 54 22 56 24
<< ntiect1 >>
rect 134 65 136 67
<< ptiect1 >>
rect 5 5 7 7
rect 134 5 136 7
<< pdifct0 >>
rect 14 55 16 57
rect 14 48 16 50
rect 24 47 26 49
rect 34 55 36 57
rect 34 48 36 50
rect 44 62 46 64
rect 44 55 46 57
rect 54 47 56 49
rect 54 40 56 42
rect 64 62 66 64
rect 64 55 66 57
rect 74 47 76 49
rect 74 40 76 42
rect 84 62 86 64
rect 84 55 86 57
rect 94 47 96 49
rect 94 40 96 42
rect 104 62 106 64
rect 104 55 106 57
rect 114 55 116 57
rect 114 48 116 50
rect 124 62 126 64
rect 124 55 126 57
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 24 40 26 42
<< alu0 >>
rect 42 62 44 64
rect 46 62 48 64
rect 12 57 38 58
rect 12 55 14 57
rect 16 55 34 57
rect 36 55 38 57
rect 12 54 38 55
rect 42 57 48 62
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 62 62 64 64
rect 66 62 68 64
rect 62 57 68 62
rect 62 55 64 57
rect 66 55 68 57
rect 62 54 68 55
rect 82 62 84 64
rect 86 62 88 64
rect 82 57 88 62
rect 82 55 84 57
rect 86 55 88 57
rect 82 54 88 55
rect 102 62 104 64
rect 106 62 108 64
rect 102 57 108 62
rect 122 62 124 64
rect 126 62 128 64
rect 102 55 104 57
rect 106 55 108 57
rect 102 54 108 55
rect 113 57 117 59
rect 113 55 114 57
rect 116 55 117 57
rect 12 50 18 54
rect 32 50 38 54
rect 113 50 117 55
rect 122 57 128 62
rect 122 55 124 57
rect 126 55 128 57
rect 122 54 128 55
rect 12 48 14 50
rect 16 48 18 50
rect 12 47 18 48
rect 22 49 28 50
rect 22 47 24 49
rect 26 47 28 49
rect 22 42 28 47
rect 32 48 34 50
rect 36 49 114 50
rect 36 48 54 49
rect 32 47 54 48
rect 56 47 74 49
rect 76 47 94 49
rect 96 48 114 49
rect 116 48 117 50
rect 96 47 117 48
rect 32 46 117 47
rect 53 42 57 46
rect 53 40 54 42
rect 56 40 57 42
rect 53 38 57 40
rect 73 42 77 46
rect 93 42 97 46
rect 73 40 74 42
rect 76 40 77 42
rect 73 38 77 40
rect 93 40 94 42
rect 96 40 97 42
rect 93 38 97 40
rect 63 23 67 25
rect 63 21 64 23
rect 66 21 67 23
rect 72 24 118 25
rect 72 22 74 24
rect 76 22 94 24
rect 96 22 114 24
rect 116 22 118 24
rect 72 21 118 22
rect 23 16 27 18
rect 23 14 24 16
rect 26 14 27 16
rect 23 8 27 14
rect 63 17 67 21
rect 93 17 97 21
rect 42 16 88 17
rect 42 14 44 16
rect 46 14 64 16
rect 66 14 84 16
rect 86 14 88 16
rect 42 13 88 14
rect 93 15 94 17
rect 96 15 97 17
rect 93 13 97 15
rect 113 17 118 21
rect 113 15 114 17
rect 116 15 118 17
rect 103 12 107 14
rect 113 13 118 15
rect 123 20 127 22
rect 123 18 124 20
rect 126 18 127 20
rect 103 10 104 12
rect 106 10 107 12
rect 103 8 107 10
rect 123 12 127 18
rect 123 10 124 12
rect 126 10 127 12
rect 123 8 127 10
<< labels >>
rlabel alu0 15 52 15 52 6 n3
rlabel alu0 65 19 65 19 6 n2
rlabel alu0 55 44 55 44 6 n3
rlabel alu0 25 56 25 56 6 n3
rlabel alu0 35 52 35 52 6 n3
rlabel ndifct0 65 15 65 15 6 n2
rlabel alu0 95 19 95 19 6 n1
rlabel alu0 95 44 95 44 6 n3
rlabel alu0 75 44 75 44 6 n3
rlabel alu0 115 19 115 19 6 n1
rlabel ndifct0 95 23 95 23 6 n1
rlabel alu0 115 52 115 52 6 n3
rlabel alu1 4 20 4 20 6 b
rlabel alu1 28 28 28 28 6 z
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 20 24 20 24 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 4 52 4 52 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 60 32 60 32 6 a3
rlabel alu1 52 32 52 32 6 a3
rlabel alu1 52 24 52 24 6 z
rlabel alu1 44 24 44 24 6 z
rlabel alu1 44 36 44 36 6 a3
rlabel alu1 72 4 72 4 6 vss
rlabel alu1 76 32 76 32 6 a2
rlabel alu1 92 32 92 32 6 a2
rlabel alu1 84 36 84 36 6 a2
rlabel alu1 72 68 72 68 6 vdd
rlabel alu1 108 32 108 32 6 a1
rlabel alu1 116 32 116 32 6 a1
rlabel alu1 124 40 124 40 6 a1
<< end >>
