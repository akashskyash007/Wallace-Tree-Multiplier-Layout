magic
tech scmos
timestamp 1199202400
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 31 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 9 30 11 33
rect 19 30 21 33
rect 9 9 11 14
rect 19 9 21 14
<< ndif >>
rect 2 18 9 30
rect 2 16 4 18
rect 6 16 9 18
rect 2 14 9 16
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 14 19 19
rect 21 21 28 30
rect 21 19 24 21
rect 26 19 28 21
rect 21 17 28 19
rect 21 14 27 17
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 42 19 59
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 68 38 70
rect 31 66 34 68
rect 36 66 38 68
rect 31 61 38 66
rect 31 59 34 61
rect 36 59 38 61
rect 31 42 38 59
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 24 46
rect 26 44 31 46
rect 2 42 31 44
rect 2 30 6 42
rect 15 37 31 38
rect 15 35 17 37
rect 19 35 31 37
rect 15 34 31 35
rect 2 28 17 30
rect 2 26 14 28
rect 16 26 17 28
rect 25 26 31 34
rect 2 25 17 26
rect 13 21 17 25
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 14 11 30
rect 19 14 21 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
<< polyct1 >>
rect 17 35 19 37
<< ndifct0 >>
rect 4 16 6 18
rect 24 19 26 21
<< ndifct1 >>
rect 14 26 16 28
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 66 16 68
rect 14 59 16 61
rect 24 51 26 53
rect 34 66 36 68
rect 34 59 36 61
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 44 26 46
<< alu0 >>
rect 13 66 14 68
rect 16 66 17 68
rect 13 61 17 66
rect 13 59 14 61
rect 16 59 17 61
rect 13 57 17 59
rect 32 66 34 68
rect 36 66 38 68
rect 32 61 38 66
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 23 53 27 55
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 3 18 7 20
rect 3 16 4 18
rect 6 16 7 18
rect 22 21 28 22
rect 22 19 24 21
rect 26 19 28 21
rect 3 12 7 16
rect 22 12 28 19
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 44 28 44 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 20 74 20 74 6 vdd
<< end >>
