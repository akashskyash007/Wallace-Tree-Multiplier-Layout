magic
tech scmos
timestamp 1199202844
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 9 39 11 49
rect 19 46 21 49
rect 29 46 31 49
rect 19 44 25 46
rect 19 42 21 44
rect 23 42 25 44
rect 19 40 25 42
rect 29 44 35 46
rect 29 42 31 44
rect 33 42 35 44
rect 29 40 35 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 36 15 37
rect 13 35 17 36
rect 9 33 17 35
rect 15 30 17 33
rect 22 30 24 40
rect 29 30 31 40
rect 39 39 41 49
rect 39 37 47 39
rect 39 35 43 37
rect 45 35 47 37
rect 36 33 47 35
rect 36 30 38 33
rect 15 6 17 10
rect 22 6 24 10
rect 29 6 31 10
rect 36 6 38 10
<< ndif >>
rect 10 22 15 30
rect 8 20 15 22
rect 8 18 10 20
rect 12 18 15 20
rect 8 16 15 18
rect 10 10 15 16
rect 17 10 22 30
rect 24 10 29 30
rect 31 10 36 30
rect 38 11 47 30
rect 38 10 42 11
rect 40 9 42 10
rect 44 9 47 11
rect 40 7 47 9
<< pdif >>
rect 43 71 49 73
rect 43 69 45 71
rect 47 69 49 71
rect 43 66 49 69
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 49 9 62
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 49 19 52
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 49 29 62
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 49 39 52
rect 41 49 49 66
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 45 71
rect 47 69 58 71
rect -2 68 58 69
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 55 38 59
rect 2 54 38 55
rect 2 52 14 54
rect 16 52 34 54
rect 36 52 38 54
rect 2 51 38 52
rect 2 49 14 51
rect 2 21 6 49
rect 42 47 46 63
rect 18 44 24 47
rect 18 42 21 44
rect 23 42 24 44
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 18 37 24 42
rect 34 43 46 47
rect 18 33 30 37
rect 34 33 38 43
rect 42 37 46 39
rect 42 35 43 37
rect 45 35 46 37
rect 10 25 22 29
rect 2 20 14 21
rect 2 18 10 20
rect 12 18 14 20
rect 2 17 14 18
rect 18 17 22 25
rect 26 17 30 33
rect 42 23 46 35
rect 34 17 46 23
rect -2 11 58 12
rect -2 9 42 11
rect 44 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 15 10 17 30
rect 22 10 24 30
rect 29 10 31 30
rect 36 10 38 30
<< pmos >>
rect 9 49 11 66
rect 19 49 21 66
rect 29 49 31 66
rect 39 49 41 66
<< polyct0 >>
rect 31 42 33 44
<< polyct1 >>
rect 21 42 23 44
rect 11 35 13 37
rect 43 35 45 37
<< ndifct1 >>
rect 10 18 12 20
rect 42 9 44 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 62 6 64
rect 14 59 16 61
rect 24 62 26 64
<< pdifct1 >>
rect 45 69 47 71
rect 14 52 16 54
rect 34 59 36 61
rect 34 52 36 54
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 23 64 27 68
rect 3 60 7 62
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 23 62 24 64
rect 26 62 27 64
rect 23 60 27 62
rect 13 55 17 59
rect 29 44 34 45
rect 29 42 31 44
rect 33 42 34 44
rect 29 41 34 42
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 d
rlabel alu1 12 32 12 32 6 d
rlabel alu1 20 40 20 40 6 c
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 20 36 20 6 a
rlabel alu1 28 24 28 24 6 c
rlabel alu1 36 40 36 40 6 b
rlabel alu1 36 60 36 60 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 56 44 56 6 b
<< end >>
