magic
tech scmos
timestamp 1199203220
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 59 11 64
rect 19 59 21 64
rect 29 59 31 64
rect 36 59 38 64
rect 46 55 48 60
rect 53 55 55 60
rect 9 35 11 39
rect 19 35 21 39
rect 9 33 21 35
rect 9 31 17 33
rect 19 31 21 33
rect 9 29 21 31
rect 29 30 31 39
rect 36 36 38 39
rect 46 36 48 39
rect 36 34 48 36
rect 53 36 55 39
rect 53 34 62 36
rect 38 32 48 34
rect 38 30 42 32
rect 44 30 48 32
rect 56 32 58 34
rect 60 32 62 34
rect 56 30 62 32
rect 9 26 11 29
rect 28 28 34 30
rect 28 26 30 28
rect 32 26 34 28
rect 28 24 34 26
rect 38 28 48 30
rect 28 21 30 24
rect 38 21 40 28
rect 28 6 30 11
rect 38 6 40 11
rect 9 2 11 6
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 6 9 13
rect 11 21 26 26
rect 11 18 28 21
rect 11 16 14 18
rect 16 16 28 18
rect 11 11 28 16
rect 30 19 38 21
rect 30 17 33 19
rect 35 17 38 19
rect 30 11 38 17
rect 40 15 48 21
rect 40 13 43 15
rect 45 13 48 15
rect 40 11 48 13
rect 11 10 26 11
rect 11 8 14 10
rect 16 8 22 10
rect 24 8 26 10
rect 11 6 26 8
<< pdif >>
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 39 9 48
rect 11 50 19 59
rect 11 48 14 50
rect 16 48 19 50
rect 11 43 19 48
rect 11 41 14 43
rect 16 41 19 43
rect 11 39 19 41
rect 21 57 29 59
rect 21 55 24 57
rect 26 55 29 57
rect 21 39 29 55
rect 31 39 36 59
rect 38 55 43 59
rect 38 49 46 55
rect 38 47 41 49
rect 43 47 46 49
rect 38 39 46 47
rect 48 39 53 55
rect 55 53 62 55
rect 55 51 58 53
rect 60 51 62 53
rect 55 39 62 51
<< alu1 >>
rect -2 67 66 72
rect -2 65 49 67
rect 51 65 57 67
rect 59 65 66 67
rect -2 64 66 65
rect 13 50 17 52
rect 13 48 14 50
rect 16 48 17 50
rect 13 43 17 48
rect 2 41 14 43
rect 16 41 17 43
rect 2 38 17 41
rect 2 26 6 38
rect 58 42 62 43
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 17 7 22
rect 29 38 62 42
rect 29 28 33 38
rect 29 26 30 28
rect 32 26 33 28
rect 29 24 33 26
rect 41 32 47 34
rect 41 30 42 32
rect 44 30 47 32
rect 58 34 62 38
rect 60 32 62 34
rect 41 27 47 30
rect 58 29 62 32
rect 41 21 54 27
rect 2 15 4 17
rect 6 15 7 17
rect 2 13 7 15
rect -2 7 66 8
rect -2 5 57 7
rect 59 5 66 7
rect -2 0 66 5
<< ptie >>
rect 55 7 61 26
rect 55 5 57 7
rect 59 5 61 7
rect 55 3 61 5
<< ntie >>
rect 47 67 61 69
rect 47 65 49 67
rect 51 65 57 67
rect 59 65 61 67
rect 47 63 61 65
<< nmos >>
rect 9 6 11 26
rect 28 11 30 21
rect 38 11 40 21
<< pmos >>
rect 9 39 11 59
rect 19 39 21 59
rect 29 39 31 59
rect 36 39 38 59
rect 46 39 48 55
rect 53 39 55 55
<< polyct0 >>
rect 17 31 19 33
<< polyct1 >>
rect 42 30 44 32
rect 58 32 60 34
rect 30 26 32 28
<< ndifct0 >>
rect 14 16 16 18
rect 33 17 35 19
rect 43 13 45 15
rect 14 8 16 10
rect 22 8 24 10
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
<< ntiect1 >>
rect 49 65 51 67
rect 57 65 59 67
<< ptiect1 >>
rect 57 5 59 7
<< pdifct0 >>
rect 4 55 6 57
rect 4 48 6 50
rect 24 55 26 57
rect 41 47 43 49
rect 58 51 60 53
<< pdifct1 >>
rect 14 48 16 50
rect 14 41 16 43
<< alu0 >>
rect 2 57 8 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 50 8 55
rect 22 57 28 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 57 53 61 64
rect 2 48 4 50
rect 6 48 8 50
rect 2 47 8 48
rect 57 51 58 53
rect 60 51 61 53
rect 21 49 45 50
rect 57 49 61 51
rect 21 47 41 49
rect 43 47 45 49
rect 21 46 45 47
rect 21 34 25 46
rect 15 33 25 34
rect 15 31 17 33
rect 19 31 25 33
rect 15 30 25 31
rect 21 20 25 30
rect 56 31 58 38
rect 13 18 17 20
rect 13 16 14 18
rect 16 16 17 18
rect 21 19 37 20
rect 21 17 33 19
rect 35 17 37 19
rect 21 16 37 17
rect 13 10 17 16
rect 42 15 46 17
rect 42 13 43 15
rect 45 13 46 15
rect 13 8 14 10
rect 16 8 17 10
rect 21 10 25 12
rect 21 8 22 10
rect 24 8 25 10
rect 42 8 46 13
<< labels >>
rlabel alu0 29 18 29 18 6 zn
rlabel alu0 20 32 20 32 6 zn
rlabel alu0 33 48 33 48 6 zn
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 44 28 44 28 6 b
rlabel alu1 44 40 44 40 6 a
rlabel alu1 36 40 36 40 6 a
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 24 52 24 6 b
rlabel alu1 60 36 60 36 6 a
rlabel alu1 52 40 52 40 6 a
<< end >>
