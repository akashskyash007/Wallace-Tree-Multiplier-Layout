magic
tech scmos
timestamp 1199472698
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -2 48 52 104
<< pwell >>
rect -2 -4 52 48
<< alu1 >>
rect -2 95 52 100
rect -2 93 5 95
rect 7 93 14 95
rect 16 93 24 95
rect 26 93 34 95
rect 36 93 43 95
rect 45 93 52 95
rect -2 88 52 93
rect -2 7 52 12
rect -2 5 5 7
rect 7 5 14 7
rect 16 5 24 7
rect 26 5 34 7
rect 36 5 43 7
rect 45 5 52 7
rect -2 0 52 5
<< ptie >>
rect 3 7 47 39
rect 3 5 5 7
rect 7 5 14 7
rect 16 5 24 7
rect 26 5 34 7
rect 36 5 43 7
rect 45 5 47 7
rect 3 3 47 5
<< ntie >>
rect 3 95 47 97
rect 3 93 5 95
rect 7 93 14 95
rect 16 93 24 95
rect 26 93 34 95
rect 36 93 43 95
rect 45 93 47 95
rect 3 55 47 93
<< ntiect1 >>
rect 5 93 7 95
rect 14 93 16 95
rect 24 93 26 95
rect 34 93 36 95
rect 43 93 45 95
<< ptiect1 >>
rect 5 5 7 7
rect 14 5 16 7
rect 24 5 26 7
rect 34 5 36 7
rect 43 5 45 7
<< labels >>
rlabel ptiect1 25 6 25 6 6 vss
rlabel ntiect1 25 94 25 94 6 vdd
<< end >>
