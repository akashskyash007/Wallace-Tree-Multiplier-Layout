magic
tech scmos
timestamp 1199469786
<< ab >>
rect 0 0 40 100
<< nwell >>
rect -2 48 42 104
<< pwell >>
rect -2 -4 42 48
<< poly >>
rect 13 83 15 88
rect 25 83 27 88
rect 13 46 15 71
rect 25 63 27 71
rect 25 61 31 63
rect 25 59 27 61
rect 29 59 31 61
rect 25 57 31 59
rect 13 44 23 46
rect 17 42 19 44
rect 21 42 23 44
rect 17 40 23 42
rect 19 37 21 40
rect 27 37 29 57
rect 19 22 21 27
rect 27 22 29 27
<< ndif >>
rect 14 33 19 37
rect 11 31 19 33
rect 11 29 13 31
rect 15 29 19 31
rect 11 27 19 29
rect 21 27 27 37
rect 29 31 37 37
rect 29 29 33 31
rect 35 29 37 31
rect 29 27 37 29
<< pdif >>
rect 3 81 13 83
rect 3 79 7 81
rect 9 79 13 81
rect 3 71 13 79
rect 15 75 25 83
rect 15 73 19 75
rect 21 73 25 75
rect 15 71 25 73
rect 27 81 37 83
rect 27 79 31 81
rect 33 79 37 81
rect 27 71 37 79
<< alu1 >>
rect -2 95 42 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 42 95
rect -2 88 42 93
rect 6 81 10 88
rect 6 79 7 81
rect 9 79 10 81
rect 6 77 10 79
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 77 34 79
rect 17 75 23 76
rect 17 73 19 75
rect 21 73 23 75
rect 8 68 23 73
rect 8 32 12 68
rect 18 61 32 63
rect 18 59 27 61
rect 29 59 32 61
rect 18 57 32 59
rect 18 44 22 53
rect 28 47 32 57
rect 18 42 19 44
rect 21 43 22 44
rect 21 42 32 43
rect 18 37 32 42
rect 8 31 17 32
rect 8 29 13 31
rect 15 29 17 31
rect 8 27 17 29
rect 32 31 36 33
rect 32 29 33 31
rect 35 29 36 31
rect 32 12 36 29
rect -2 7 42 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 42 7
rect -2 0 42 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 19 27 21 37
rect 27 27 29 37
<< pmos >>
rect 13 71 15 83
rect 25 71 27 83
<< polyct1 >>
rect 27 59 29 61
rect 19 42 21 44
<< ndifct1 >>
rect 13 29 15 31
rect 33 29 35 31
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 7 79 9 81
rect 19 73 21 75
rect 31 79 33 81
<< labels >>
rlabel alu1 10 50 10 50 6 z
rlabel ptiect1 20 6 20 6 6 vss
rlabel alu1 20 45 20 45 6 b
rlabel alu1 20 60 20 60 6 a
rlabel alu1 20 70 20 70 6 z
rlabel ntiect1 20 94 20 94 6 vdd
rlabel alu1 30 40 30 40 6 b
rlabel alu1 30 55 30 55 6 a
<< end >>
