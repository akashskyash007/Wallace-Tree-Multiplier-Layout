magic
tech scmos
timestamp 1199542746
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -5 48 55 105
<< pwell >>
rect -5 -5 55 48
<< poly >>
rect 19 94 21 98
rect 27 94 29 98
rect 35 94 37 98
rect 19 53 21 56
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 11 47 23 49
rect 11 25 13 47
rect 27 43 29 56
rect 35 53 37 56
rect 35 51 39 53
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 23 37 33 39
rect 23 25 25 37
rect 37 33 39 51
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 35 27 43 29
rect 35 24 37 27
rect 11 11 13 15
rect 23 11 25 15
rect 35 10 37 14
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 25 24 30 25
rect 25 21 35 24
rect 25 19 29 21
rect 31 19 35 21
rect 25 15 35 19
rect 15 11 21 15
rect 27 14 35 15
rect 37 14 45 24
rect 15 9 17 11
rect 19 9 21 11
rect 39 11 45 14
rect 15 7 21 9
rect 39 9 41 11
rect 43 9 45 11
rect 39 7 45 9
<< pdif >>
rect 14 85 19 94
rect 7 81 19 85
rect 7 79 9 81
rect 11 79 19 81
rect 7 71 19 79
rect 7 69 9 71
rect 11 69 19 71
rect 7 61 19 69
rect 7 59 9 61
rect 11 59 19 61
rect 7 56 19 59
rect 21 56 27 94
rect 29 56 35 94
rect 37 91 45 94
rect 37 89 41 91
rect 43 89 45 91
rect 37 56 45 89
rect 7 55 13 56
<< alu1 >>
rect -2 91 52 100
rect -2 89 41 91
rect 43 89 52 91
rect -2 88 52 89
rect 8 81 12 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 71 12 79
rect 8 69 9 71
rect 11 69 12 71
rect 8 61 12 69
rect 8 59 9 61
rect 11 59 12 61
rect 8 22 12 59
rect 18 51 22 83
rect 18 49 19 51
rect 21 49 22 51
rect 18 27 22 49
rect 28 41 32 83
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 31 42 83
rect 38 29 39 31
rect 41 29 42 31
rect 3 21 33 22
rect 3 19 5 21
rect 7 19 29 21
rect 31 19 33 21
rect 3 18 33 19
rect 38 17 42 29
rect -2 11 52 12
rect -2 9 17 11
rect 19 9 41 11
rect 43 9 52 11
rect -2 0 52 9
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 14 37 24
<< pmos >>
rect 19 56 21 94
rect 27 56 29 94
rect 35 56 37 94
<< polyct1 >>
rect 19 49 21 51
rect 29 39 31 41
rect 39 29 41 31
<< ndifct1 >>
rect 5 19 7 21
rect 29 19 31 21
rect 17 9 19 11
rect 41 9 43 11
<< pdifct1 >>
rect 9 79 11 81
rect 9 69 11 71
rect 9 59 11 61
rect 41 89 43 91
<< labels >>
rlabel alu1 20 20 20 20 6 nq
rlabel alu1 10 50 10 50 6 nq
rlabel alu1 20 55 20 55 6 i1
rlabel alu1 25 6 25 6 6 vss
rlabel ndifct1 30 20 30 20 6 nq
rlabel alu1 30 55 30 55 6 i0
rlabel alu1 25 94 25 94 6 vdd
rlabel alu1 40 50 40 50 6 i2
<< end >>
