magic
tech scmos
timestamp 1199202196
<< ab >>
rect 0 0 144 72
<< nwell >>
rect -5 32 149 77
<< pwell >>
rect -5 -5 149 32
<< poly >>
rect 9 66 11 70
rect 55 68 111 70
rect 55 60 57 68
rect 65 60 67 64
rect 75 60 77 64
rect 82 60 84 68
rect 92 60 94 64
rect 99 60 101 64
rect 19 52 21 57
rect 38 54 40 59
rect 45 54 47 59
rect 9 34 11 38
rect 19 35 21 38
rect 9 32 15 34
rect 19 33 34 35
rect 9 30 11 32
rect 13 30 15 32
rect 9 28 15 30
rect 27 31 30 33
rect 32 31 34 33
rect 27 29 34 31
rect 9 24 11 28
rect 27 26 29 29
rect 38 19 40 48
rect 45 44 47 48
rect 45 42 51 44
rect 45 40 47 42
rect 49 40 51 42
rect 45 38 51 40
rect 55 34 57 48
rect 45 32 57 34
rect 45 19 47 32
rect 65 29 67 48
rect 75 44 77 54
rect 71 42 77 44
rect 71 40 73 42
rect 75 40 77 42
rect 71 38 77 40
rect 51 26 57 28
rect 51 24 53 26
rect 55 24 57 26
rect 51 22 57 24
rect 55 19 57 22
rect 65 27 71 29
rect 65 25 67 27
rect 69 25 71 27
rect 65 23 71 25
rect 65 19 67 23
rect 75 19 77 38
rect 82 34 84 54
rect 109 58 111 68
rect 129 59 131 64
rect 92 44 94 47
rect 88 42 94 44
rect 88 40 90 42
rect 92 40 94 42
rect 88 38 94 40
rect 99 35 101 47
rect 109 44 111 47
rect 129 45 131 49
rect 109 42 117 44
rect 115 35 117 42
rect 122 43 131 45
rect 122 41 124 43
rect 126 41 131 43
rect 122 39 131 41
rect 82 32 94 34
rect 82 26 88 28
rect 82 24 84 26
rect 86 24 88 26
rect 82 22 88 24
rect 82 19 84 22
rect 92 19 94 32
rect 99 33 105 35
rect 99 31 101 33
rect 103 31 105 33
rect 99 29 105 31
rect 115 33 121 35
rect 115 31 117 33
rect 119 31 121 33
rect 115 29 121 31
rect 99 19 101 29
rect 119 26 121 29
rect 129 26 131 39
rect 27 14 29 19
rect 119 15 121 20
rect 129 14 131 19
rect 9 7 11 10
rect 38 7 40 13
rect 45 8 47 13
rect 9 5 40 7
rect 55 4 57 13
rect 65 8 67 13
rect 75 8 77 13
rect 82 4 84 13
rect 92 8 94 13
rect 99 8 101 13
rect 55 2 84 4
<< ndif >>
rect 20 24 27 26
rect 2 22 9 24
rect 2 20 4 22
rect 6 20 9 22
rect 2 18 9 20
rect 4 10 9 18
rect 11 16 16 24
rect 20 22 22 24
rect 24 22 27 24
rect 20 20 27 22
rect 22 19 27 20
rect 29 19 36 26
rect 112 24 119 26
rect 112 22 114 24
rect 116 22 119 24
rect 112 20 119 22
rect 121 24 129 26
rect 121 22 124 24
rect 126 22 129 24
rect 121 20 129 22
rect 11 14 18 16
rect 31 17 38 19
rect 31 15 33 17
rect 35 15 38 17
rect 11 12 14 14
rect 16 12 18 14
rect 31 13 38 15
rect 40 13 45 19
rect 47 17 55 19
rect 47 15 50 17
rect 52 15 55 17
rect 47 13 55 15
rect 57 17 65 19
rect 57 15 60 17
rect 62 15 65 17
rect 57 13 65 15
rect 67 17 75 19
rect 67 15 70 17
rect 72 15 75 17
rect 67 13 75 15
rect 77 13 82 19
rect 84 17 92 19
rect 84 15 87 17
rect 89 15 92 17
rect 84 13 92 15
rect 94 13 99 19
rect 101 17 108 19
rect 101 15 104 17
rect 106 15 108 17
rect 123 19 129 20
rect 131 24 138 26
rect 131 22 134 24
rect 136 22 138 24
rect 131 19 138 22
rect 101 13 108 15
rect 11 10 18 12
<< pdif >>
rect 4 52 9 66
rect 2 49 9 52
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 18 66
rect 11 62 14 64
rect 16 62 18 64
rect 11 60 18 62
rect 11 52 17 60
rect 50 54 55 60
rect 30 52 38 54
rect 11 50 19 52
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 44 26 52
rect 30 50 32 52
rect 34 50 38 52
rect 30 48 38 50
rect 40 48 45 54
rect 47 52 55 54
rect 47 50 50 52
rect 52 50 55 52
rect 47 48 55 50
rect 57 52 65 60
rect 57 50 60 52
rect 62 50 65 52
rect 57 48 65 50
rect 67 58 75 60
rect 67 56 70 58
rect 72 56 75 58
rect 67 54 75 56
rect 77 54 82 60
rect 84 58 92 60
rect 84 56 87 58
rect 89 56 92 58
rect 84 54 92 56
rect 67 48 73 54
rect 21 42 28 44
rect 21 40 24 42
rect 26 40 28 42
rect 21 38 28 40
rect 87 47 92 54
rect 94 47 99 60
rect 101 58 106 60
rect 101 56 109 58
rect 101 54 104 56
rect 106 54 109 56
rect 101 47 109 54
rect 111 53 116 58
rect 122 57 129 59
rect 122 55 124 57
rect 126 55 129 57
rect 111 51 118 53
rect 111 49 114 51
rect 116 49 118 51
rect 122 49 129 55
rect 131 55 136 59
rect 131 53 138 55
rect 131 51 134 53
rect 136 51 138 53
rect 131 49 138 51
rect 111 47 118 49
<< alu1 >>
rect -2 67 146 72
rect -2 65 28 67
rect 30 65 38 67
rect 40 65 119 67
rect 121 65 146 67
rect -2 64 146 65
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 2 40 4 42
rect 6 40 15 42
rect 2 38 15 40
rect 2 24 6 38
rect 2 22 7 24
rect 2 20 4 22
rect 6 20 7 22
rect 2 18 7 20
rect 121 43 127 50
rect 121 42 124 43
rect 97 34 103 42
rect 113 41 124 42
rect 126 41 127 43
rect 113 38 127 41
rect 97 33 111 34
rect 97 31 101 33
rect 103 31 111 33
rect 97 30 111 31
rect -2 7 146 8
rect -2 5 120 7
rect 122 5 131 7
rect 133 5 146 7
rect -2 0 146 5
<< ptie >>
rect 112 7 141 9
rect 112 5 120 7
rect 122 5 131 7
rect 133 5 141 7
rect 112 3 141 5
<< ntie >>
rect 22 67 46 69
rect 22 65 28 67
rect 30 65 38 67
rect 40 65 46 67
rect 22 63 46 65
rect 117 67 123 69
rect 117 65 119 67
rect 121 65 123 67
rect 117 63 123 65
<< nmos >>
rect 9 10 11 24
rect 27 19 29 26
rect 119 20 121 26
rect 38 13 40 19
rect 45 13 47 19
rect 55 13 57 19
rect 65 13 67 19
rect 75 13 77 19
rect 82 13 84 19
rect 92 13 94 19
rect 99 13 101 19
rect 129 19 131 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 52
rect 38 48 40 54
rect 45 48 47 54
rect 55 48 57 60
rect 65 48 67 60
rect 75 54 77 60
rect 82 54 84 60
rect 92 47 94 60
rect 99 47 101 60
rect 109 47 111 58
rect 129 49 131 59
<< polyct0 >>
rect 11 30 13 32
rect 30 31 32 33
rect 47 40 49 42
rect 73 40 75 42
rect 53 24 55 26
rect 67 25 69 27
rect 90 40 92 42
rect 84 24 86 26
rect 117 31 119 33
<< polyct1 >>
rect 124 41 126 43
rect 101 31 103 33
<< ndifct0 >>
rect 22 22 24 24
rect 114 22 116 24
rect 124 22 126 24
rect 33 15 35 17
rect 14 12 16 14
rect 50 15 52 17
rect 60 15 62 17
rect 70 15 72 17
rect 87 15 89 17
rect 104 15 106 17
rect 134 22 136 24
<< ndifct1 >>
rect 4 20 6 22
<< ntiect1 >>
rect 28 65 30 67
rect 38 65 40 67
rect 119 65 121 67
<< ptiect1 >>
rect 120 5 122 7
rect 131 5 133 7
<< pdifct0 >>
rect 14 62 16 64
rect 14 48 16 50
rect 32 50 34 52
rect 50 50 52 52
rect 60 50 62 52
rect 70 56 72 58
rect 87 56 89 58
rect 24 40 26 42
rect 104 54 106 56
rect 124 55 126 57
rect 114 49 116 51
rect 134 51 136 53
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
<< alu0 >>
rect 13 62 14 64
rect 16 62 17 64
rect 13 50 17 62
rect 13 48 14 50
rect 16 48 17 50
rect 31 52 35 64
rect 69 58 73 64
rect 69 56 70 58
rect 72 56 73 58
rect 69 54 73 56
rect 81 58 91 59
rect 81 56 87 58
rect 89 56 91 58
rect 81 55 91 56
rect 102 56 108 64
rect 31 50 32 52
rect 34 50 35 52
rect 31 48 35 50
rect 38 52 54 53
rect 38 50 50 52
rect 52 50 54 52
rect 38 49 54 50
rect 59 52 63 54
rect 59 50 60 52
rect 62 50 63 52
rect 13 46 17 48
rect 21 42 28 43
rect 21 40 24 42
rect 26 40 28 42
rect 21 39 28 40
rect 21 33 25 39
rect 38 34 42 49
rect 59 43 63 50
rect 45 42 54 43
rect 45 40 47 42
rect 49 40 54 42
rect 45 39 54 40
rect 9 32 25 33
rect 9 30 11 32
rect 13 30 25 32
rect 28 33 44 34
rect 28 31 30 33
rect 32 31 44 33
rect 28 30 44 31
rect 9 29 25 30
rect 21 24 25 29
rect 21 22 22 24
rect 24 22 25 24
rect 21 20 25 22
rect 32 17 36 19
rect 13 14 17 16
rect 13 12 14 14
rect 16 12 17 14
rect 13 8 17 12
rect 32 15 33 17
rect 35 15 36 17
rect 32 8 36 15
rect 40 18 44 30
rect 50 28 54 39
rect 59 42 77 43
rect 59 40 73 42
rect 75 40 77 42
rect 59 39 77 40
rect 50 26 56 28
rect 50 24 53 26
rect 55 24 56 26
rect 50 22 56 24
rect 40 17 54 18
rect 40 15 50 17
rect 52 15 54 17
rect 40 14 54 15
rect 59 17 63 39
rect 81 36 85 55
rect 102 54 104 56
rect 106 54 108 56
rect 122 57 128 64
rect 122 55 124 57
rect 126 55 128 57
rect 122 54 128 55
rect 102 53 108 54
rect 133 53 137 55
rect 113 51 117 53
rect 113 50 114 51
rect 76 32 85 36
rect 89 49 114 50
rect 116 49 117 51
rect 133 51 134 53
rect 136 51 137 53
rect 89 46 117 49
rect 89 42 93 46
rect 89 40 90 42
rect 92 40 93 42
rect 76 29 80 32
rect 66 27 80 29
rect 89 28 93 40
rect 133 34 137 51
rect 115 33 137 34
rect 115 31 117 33
rect 119 31 137 33
rect 115 30 137 31
rect 66 25 67 27
rect 69 25 80 27
rect 66 23 80 25
rect 59 15 60 17
rect 62 15 63 17
rect 59 13 63 15
rect 69 17 73 19
rect 69 15 70 17
rect 72 15 73 17
rect 69 8 73 15
rect 76 18 80 23
rect 83 26 93 28
rect 83 24 84 26
rect 86 24 118 26
rect 83 22 114 24
rect 116 22 118 24
rect 112 21 118 22
rect 123 24 127 26
rect 123 22 124 24
rect 126 22 127 24
rect 76 17 91 18
rect 76 15 87 17
rect 89 15 91 17
rect 76 14 91 15
rect 102 17 108 18
rect 102 15 104 17
rect 106 15 108 17
rect 102 8 108 15
rect 123 8 127 22
rect 133 24 137 30
rect 133 22 134 24
rect 136 22 137 24
rect 133 20 137 22
<< labels >>
rlabel alu0 17 31 17 31 6 zn
rlabel alu0 23 31 23 31 6 zn
rlabel alu0 47 16 47 16 6 n4
rlabel alu0 36 32 36 32 6 n4
rlabel alu0 53 25 53 25 6 ci
rlabel alu0 46 51 46 51 6 n4
rlabel alu0 49 41 49 41 6 ci
rlabel alu0 61 33 61 33 6 n2
rlabel alu0 83 16 83 16 6 n1
rlabel alu0 73 26 73 26 6 n1
rlabel alu0 91 36 91 36 6 ci
rlabel alu0 68 41 68 41 6 n2
rlabel alu0 86 57 86 57 6 n1
rlabel alu0 100 24 100 24 6 ci
rlabel alu0 126 32 126 32 6 cn
rlabel alu0 115 49 115 49 6 ci
rlabel alu0 135 37 135 37 6 cn
rlabel alu1 12 40 12 40 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 72 4 72 4 6 vss
rlabel alu1 100 36 100 36 6 d
rlabel alu1 72 68 72 68 6 vdd
rlabel alu1 108 32 108 32 6 d
rlabel alu1 116 40 116 40 6 cp
rlabel alu1 124 44 124 44 6 cp
<< end >>
