magic
tech scmos
timestamp 1199470350
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 25 94 27 98
rect 37 94 39 98
rect 45 94 47 98
rect 57 94 59 98
rect 65 94 67 98
rect 25 52 27 55
rect 25 50 31 52
rect 25 48 27 50
rect 29 48 31 50
rect 12 46 31 48
rect 12 36 14 46
rect 37 43 39 55
rect 45 52 47 55
rect 45 50 53 52
rect 45 48 49 50
rect 51 48 53 50
rect 45 46 53 48
rect 35 41 41 43
rect 35 40 37 41
rect 33 39 37 40
rect 39 39 41 41
rect 33 37 41 39
rect 33 34 35 37
rect 45 34 47 46
rect 57 43 59 55
rect 65 52 67 55
rect 65 50 73 52
rect 65 49 69 50
rect 67 48 69 49
rect 71 48 73 50
rect 67 46 73 48
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 57 34 59 37
rect 67 34 69 46
rect 12 12 14 17
rect 33 12 35 17
rect 45 12 47 17
rect 57 12 59 17
rect 67 12 69 17
<< ndif >>
rect 3 31 12 36
rect 3 29 6 31
rect 8 29 12 31
rect 3 21 12 29
rect 3 19 6 21
rect 8 19 12 21
rect 3 17 12 19
rect 14 34 22 36
rect 14 32 18 34
rect 20 32 22 34
rect 14 30 22 32
rect 14 17 19 30
rect 28 23 33 34
rect 25 21 33 23
rect 25 19 27 21
rect 29 19 33 21
rect 25 17 33 19
rect 35 31 45 34
rect 35 29 39 31
rect 41 29 45 31
rect 35 17 45 29
rect 47 21 57 34
rect 47 19 51 21
rect 53 19 57 21
rect 47 17 57 19
rect 59 17 67 34
rect 69 31 74 34
rect 69 29 77 31
rect 69 27 73 29
rect 75 27 77 29
rect 69 21 77 27
rect 69 19 73 21
rect 75 19 77 21
rect 69 17 77 19
rect 61 10 65 17
rect 61 8 67 10
rect 61 6 63 8
rect 65 6 67 8
rect 61 4 67 6
<< pdif >>
rect 20 69 25 94
rect 17 67 25 69
rect 17 65 19 67
rect 21 65 25 67
rect 17 59 25 65
rect 17 57 19 59
rect 21 57 25 59
rect 17 55 25 57
rect 27 91 37 94
rect 27 89 31 91
rect 33 89 37 91
rect 27 81 37 89
rect 27 79 31 81
rect 33 79 37 81
rect 27 55 37 79
rect 39 55 45 94
rect 47 81 57 94
rect 47 79 51 81
rect 53 79 57 81
rect 47 73 57 79
rect 47 71 51 73
rect 53 71 57 73
rect 47 55 57 71
rect 59 55 65 94
rect 67 91 76 94
rect 67 89 71 91
rect 73 89 76 91
rect 67 81 76 89
rect 67 79 71 81
rect 73 79 76 81
rect 67 55 76 79
<< alu1 >>
rect -2 95 82 100
rect -2 93 9 95
rect 11 93 82 95
rect -2 91 82 93
rect -2 89 31 91
rect 33 89 71 91
rect 73 89 82 91
rect -2 88 82 89
rect 18 67 22 83
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 77 34 79
rect 50 81 54 83
rect 50 79 51 81
rect 53 79 54 81
rect 50 73 54 79
rect 70 81 74 88
rect 70 79 71 81
rect 73 79 74 81
rect 70 77 74 79
rect 50 72 51 73
rect 18 65 19 67
rect 21 65 22 67
rect 18 59 22 65
rect 18 57 19 59
rect 21 57 22 59
rect 18 42 22 57
rect 28 71 51 72
rect 53 71 54 73
rect 28 68 54 71
rect 28 52 32 68
rect 58 67 72 73
rect 26 50 32 52
rect 26 48 27 50
rect 29 48 32 50
rect 26 46 32 48
rect 7 38 22 42
rect 17 34 22 38
rect 5 31 9 33
rect 5 29 6 31
rect 8 29 9 31
rect 5 21 9 29
rect 17 32 18 34
rect 20 32 22 34
rect 17 27 22 32
rect 28 32 32 46
rect 38 58 53 63
rect 38 43 42 58
rect 36 41 42 43
rect 36 39 37 41
rect 39 39 42 41
rect 36 37 42 39
rect 48 50 52 53
rect 48 48 49 50
rect 51 48 52 50
rect 48 32 52 48
rect 57 42 62 63
rect 68 50 72 67
rect 68 48 69 50
rect 71 48 72 50
rect 68 46 72 48
rect 57 41 73 42
rect 57 39 59 41
rect 61 39 73 41
rect 57 38 73 39
rect 28 31 43 32
rect 28 29 39 31
rect 41 29 43 31
rect 28 28 43 29
rect 48 27 63 32
rect 71 29 77 30
rect 71 27 73 29
rect 75 27 77 29
rect 71 22 77 27
rect 5 19 6 21
rect 8 19 9 21
rect 5 12 9 19
rect 25 21 77 22
rect 25 19 27 21
rect 29 19 51 21
rect 53 19 73 21
rect 75 19 77 21
rect 25 18 77 19
rect -2 8 82 12
rect -2 7 63 8
rect -2 5 9 7
rect 11 5 19 7
rect 21 6 63 7
rect 65 6 82 8
rect 21 5 82 6
rect -2 0 82 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 13 97
rect 7 93 9 95
rect 11 93 13 95
rect 7 91 13 93
<< nmos >>
rect 12 17 14 36
rect 33 17 35 34
rect 45 17 47 34
rect 57 17 59 34
rect 67 17 69 34
<< pmos >>
rect 25 55 27 94
rect 37 55 39 94
rect 45 55 47 94
rect 57 55 59 94
rect 65 55 67 94
<< polyct1 >>
rect 27 48 29 50
rect 49 48 51 50
rect 37 39 39 41
rect 69 48 71 50
rect 59 39 61 41
<< ndifct1 >>
rect 6 29 8 31
rect 6 19 8 21
rect 18 32 20 34
rect 27 19 29 21
rect 39 29 41 31
rect 51 19 53 21
rect 73 27 75 29
rect 73 19 75 21
rect 63 6 65 8
<< ntiect1 >>
rect 9 93 11 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 19 65 21 67
rect 19 57 21 59
rect 31 89 33 91
rect 31 79 33 81
rect 51 79 53 81
rect 51 71 53 73
rect 71 89 73 91
rect 71 79 73 81
<< labels >>
rlabel ndifct1 28 20 28 20 6 n3
rlabel polyct1 28 49 28 49 6 zn
rlabel ndifct1 52 20 52 20 6 n3
rlabel ndifct1 40 30 40 30 6 zn
rlabel pdifct1 52 72 52 72 6 zn
rlabel pdifct1 52 80 52 80 6 zn
rlabel ndifct1 74 20 74 20 6 n3
rlabel ndifct1 74 28 74 28 6 n3
rlabel alu1 10 40 10 40 6 z
rlabel alu1 20 55 20 55 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 50 40 50 40 6 b2
rlabel alu1 40 50 40 50 6 b1
rlabel alu1 50 60 50 60 6 b1
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 60 30 60 30 6 b2
rlabel alu1 70 40 70 40 6 a2
rlabel alu1 60 50 60 50 6 a2
rlabel alu1 60 70 60 70 6 a1
rlabel alu1 70 60 70 60 6 a1
<< end >>
