magic
tech scmos
timestamp 1199202122
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 26 67 48 69
rect 9 58 11 63
rect 19 58 21 63
rect 26 58 28 67
rect 36 58 38 63
rect 46 58 48 67
rect 58 62 60 67
rect 9 37 11 42
rect 19 37 21 42
rect 9 35 21 37
rect 9 32 11 35
rect 5 30 11 32
rect 19 30 21 35
rect 26 30 28 42
rect 36 39 38 42
rect 32 37 38 39
rect 32 35 34 37
rect 36 35 38 37
rect 32 33 38 35
rect 36 30 38 33
rect 46 39 48 42
rect 58 39 60 42
rect 46 37 53 39
rect 46 35 49 37
rect 51 35 53 37
rect 46 33 53 35
rect 57 37 63 39
rect 57 35 59 37
rect 61 35 63 37
rect 57 33 63 35
rect 46 30 48 33
rect 58 30 60 33
rect 5 28 7 30
rect 9 28 11 30
rect 5 26 11 28
rect 9 23 11 26
rect 19 18 21 23
rect 26 18 28 23
rect 36 18 38 23
rect 46 18 48 23
rect 9 11 11 16
rect 58 15 60 20
<< ndif >>
rect 13 23 19 30
rect 21 23 26 30
rect 28 28 36 30
rect 28 26 31 28
rect 33 26 36 28
rect 28 23 36 26
rect 38 27 46 30
rect 38 25 41 27
rect 43 25 46 27
rect 38 23 46 25
rect 48 23 58 30
rect 2 20 9 23
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 17 23
rect 50 20 58 23
rect 60 28 67 30
rect 60 26 63 28
rect 65 26 67 28
rect 60 24 67 26
rect 60 20 65 24
rect 50 19 56 20
rect 50 17 52 19
rect 54 17 56 19
rect 13 11 19 16
rect 50 15 56 17
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 65 19 69
rect 13 58 17 65
rect 50 60 58 62
rect 50 58 52 60
rect 54 58 58 60
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 4 42 9 45
rect 11 42 19 58
rect 21 42 26 58
rect 28 54 36 58
rect 28 52 31 54
rect 33 52 36 54
rect 28 42 36 52
rect 38 56 46 58
rect 38 54 41 56
rect 43 54 46 56
rect 38 49 46 54
rect 38 47 41 49
rect 43 47 46 49
rect 38 42 46 47
rect 48 42 58 58
rect 60 60 67 62
rect 60 58 63 60
rect 65 58 67 60
rect 60 53 67 58
rect 60 51 63 53
rect 65 51 67 53
rect 60 49 67 51
rect 60 42 65 49
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 71 74 79
rect -2 69 15 71
rect 17 69 74 71
rect -2 68 74 69
rect 10 54 35 55
rect 10 52 31 54
rect 33 52 35 54
rect 10 51 35 52
rect 10 49 22 51
rect 2 31 6 39
rect 2 30 14 31
rect 2 28 7 30
rect 9 28 14 30
rect 2 25 14 28
rect 18 30 22 49
rect 26 38 30 47
rect 49 46 55 54
rect 49 42 63 46
rect 26 37 39 38
rect 26 35 34 37
rect 36 35 39 37
rect 26 34 39 35
rect 18 28 35 30
rect 57 37 63 42
rect 57 35 59 37
rect 61 35 63 37
rect 57 34 63 35
rect 18 26 31 28
rect 33 26 35 28
rect 18 25 35 26
rect -2 11 74 12
rect -2 9 15 11
rect 17 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 19 23 21 30
rect 26 23 28 30
rect 36 23 38 30
rect 46 23 48 30
rect 9 16 11 23
rect 58 20 60 30
<< pmos >>
rect 9 42 11 58
rect 19 42 21 58
rect 26 42 28 58
rect 36 42 38 58
rect 46 42 48 58
rect 58 42 60 62
<< polyct0 >>
rect 49 35 51 37
<< polyct1 >>
rect 34 35 36 37
rect 59 35 61 37
rect 7 28 9 30
<< ndifct0 >>
rect 41 25 43 27
rect 4 18 6 20
rect 63 26 65 28
rect 52 17 54 19
<< ndifct1 >>
rect 31 26 33 28
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 52 58 54 60
rect 4 54 6 56
rect 4 47 6 49
rect 41 54 43 56
rect 41 47 43 49
rect 63 58 65 60
rect 63 51 65 53
<< pdifct1 >>
rect 15 69 17 71
rect 31 52 33 54
<< alu0 >>
rect 3 59 44 63
rect 3 56 7 59
rect 3 54 4 56
rect 6 54 7 56
rect 40 56 44 59
rect 50 60 56 68
rect 50 58 52 60
rect 54 58 56 60
rect 50 57 56 58
rect 62 60 66 62
rect 62 58 63 60
rect 65 58 66 60
rect 3 49 7 54
rect 40 54 41 56
rect 43 54 44 56
rect 3 47 4 49
rect 6 47 7 49
rect 3 45 7 47
rect 40 49 44 54
rect 40 47 41 49
rect 43 47 44 49
rect 40 45 44 47
rect 62 53 66 58
rect 62 51 63 53
rect 65 51 70 53
rect 62 49 70 51
rect 48 37 52 39
rect 48 35 49 37
rect 51 35 52 37
rect 48 29 52 35
rect 66 29 70 49
rect 40 27 44 29
rect 40 25 41 27
rect 43 25 44 27
rect 48 28 70 29
rect 48 26 63 28
rect 65 26 70 28
rect 48 25 70 26
rect 40 21 44 25
rect 2 20 44 21
rect 2 18 4 20
rect 6 18 44 20
rect 2 17 44 18
rect 51 19 55 21
rect 51 17 52 19
rect 54 17 55 19
rect 51 12 55 17
<< labels >>
rlabel alu0 5 54 5 54 6 n1
rlabel alu0 42 23 42 23 6 n3
rlabel alu0 23 19 23 19 6 n3
rlabel alu0 50 32 50 32 6 bn
rlabel alu0 42 54 42 54 6 n1
rlabel alu0 59 27 59 27 6 bn
rlabel alu0 64 55 64 55 6 bn
rlabel alu1 12 28 12 28 6 a
rlabel alu1 4 32 4 32 6 a
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 28 28 28 6 z
rlabel alu1 28 44 28 44 6 c
rlabel alu1 20 40 20 40 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 36 36 36 6 c
rlabel alu1 52 48 52 48 6 b
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 40 60 40 6 b
<< end >>
