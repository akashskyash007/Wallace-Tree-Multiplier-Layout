magic
tech scmos
timestamp 1199201878
<< ab >>
rect 0 0 144 80
<< nwell >>
rect -5 36 149 88
<< pwell >>
rect -5 -8 149 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 99 70 101 74
rect 109 70 111 74
rect 119 70 121 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 99 39 101 42
rect 109 39 111 42
rect 9 37 15 39
rect 19 37 34 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 25 35 27 37
rect 29 35 34 37
rect 25 33 34 35
rect 32 30 34 33
rect 39 37 51 39
rect 39 35 43 37
rect 45 35 51 37
rect 39 33 51 35
rect 39 30 41 33
rect 49 30 51 33
rect 56 37 63 39
rect 56 35 59 37
rect 61 35 63 37
rect 56 33 63 35
rect 68 37 74 39
rect 68 35 70 37
rect 72 35 74 37
rect 68 33 74 35
rect 56 30 58 33
rect 72 30 74 33
rect 79 37 91 39
rect 79 35 83 37
rect 85 35 91 37
rect 79 33 91 35
rect 79 30 81 33
rect 89 30 91 33
rect 96 37 111 39
rect 96 35 99 37
rect 101 35 107 37
rect 109 35 111 37
rect 96 33 111 35
rect 119 39 121 42
rect 119 37 127 39
rect 119 35 123 37
rect 125 35 127 37
rect 119 33 127 35
rect 96 30 98 33
rect 32 6 34 11
rect 39 6 41 11
rect 49 6 51 11
rect 56 6 58 11
rect 72 6 74 11
rect 79 6 81 11
rect 89 6 91 11
rect 96 6 98 11
<< ndif >>
rect 23 11 32 30
rect 34 11 39 30
rect 41 21 49 30
rect 41 19 44 21
rect 46 19 49 21
rect 41 11 49 19
rect 51 11 56 30
rect 58 13 72 30
rect 58 11 64 13
rect 66 11 72 13
rect 74 11 79 30
rect 81 21 89 30
rect 81 19 84 21
rect 86 19 89 21
rect 81 11 89 19
rect 91 11 96 30
rect 98 22 106 30
rect 98 20 101 22
rect 103 20 106 22
rect 98 15 106 20
rect 98 13 101 15
rect 103 13 106 15
rect 98 11 106 13
rect 23 9 26 11
rect 28 9 30 11
rect 23 7 30 9
rect 60 9 70 11
<< pdif >>
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 55 9 60
rect 2 53 4 55
rect 6 53 9 55
rect 2 51 9 53
rect 4 42 9 51
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 62 29 70
rect 21 60 24 62
rect 26 60 29 62
rect 21 42 29 60
rect 31 53 39 70
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 62 49 70
rect 41 60 44 62
rect 46 60 49 62
rect 41 42 49 60
rect 51 53 59 70
rect 51 51 54 53
rect 56 51 59 53
rect 51 42 59 51
rect 61 61 69 70
rect 61 59 64 61
rect 66 59 69 61
rect 61 54 69 59
rect 61 52 64 54
rect 66 52 69 54
rect 61 42 69 52
rect 71 68 79 70
rect 71 66 74 68
rect 76 66 79 68
rect 71 61 79 66
rect 71 59 74 61
rect 76 59 79 61
rect 71 42 79 59
rect 81 60 89 70
rect 81 58 84 60
rect 86 58 89 60
rect 81 53 89 58
rect 81 51 84 53
rect 86 51 89 53
rect 81 42 89 51
rect 91 68 99 70
rect 91 66 94 68
rect 96 66 99 68
rect 91 61 99 66
rect 91 59 94 61
rect 96 59 99 61
rect 91 42 99 59
rect 101 60 109 70
rect 101 58 104 60
rect 106 58 109 60
rect 101 53 109 58
rect 101 51 104 53
rect 106 51 109 53
rect 101 42 109 51
rect 111 68 119 70
rect 111 66 114 68
rect 116 66 119 68
rect 111 61 119 66
rect 111 59 114 61
rect 116 59 119 61
rect 111 42 119 59
rect 121 55 126 70
rect 121 53 128 55
rect 121 51 124 53
rect 126 51 128 53
rect 121 46 128 51
rect 121 44 124 46
rect 126 44 128 46
rect 121 42 128 44
<< alu1 >>
rect -2 81 146 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 146 81
rect -2 68 146 79
rect 12 53 58 54
rect 12 51 14 53
rect 16 51 34 53
rect 36 51 54 53
rect 56 51 58 53
rect 12 50 58 51
rect 12 47 18 50
rect 2 46 18 47
rect 2 44 14 46
rect 16 44 18 46
rect 2 43 18 44
rect 2 22 6 43
rect 25 42 63 46
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 30 47 35
rect 57 37 63 42
rect 57 35 59 37
rect 61 35 63 37
rect 57 34 63 35
rect 69 42 103 46
rect 69 37 73 42
rect 97 38 103 42
rect 69 35 70 37
rect 72 35 73 37
rect 69 30 73 35
rect 10 26 47 30
rect 65 26 73 30
rect 81 37 87 38
rect 81 35 83 37
rect 85 35 87 37
rect 81 30 87 35
rect 97 37 111 38
rect 97 35 99 37
rect 101 35 107 37
rect 109 35 111 37
rect 97 34 111 35
rect 122 37 126 39
rect 122 35 123 37
rect 125 35 126 37
rect 122 30 126 35
rect 81 26 126 30
rect 2 21 88 22
rect 2 19 44 21
rect 46 19 84 21
rect 86 19 88 21
rect 2 18 88 19
rect 122 17 126 26
rect -2 11 64 12
rect 66 11 146 12
rect -2 9 26 11
rect 28 9 146 11
rect -2 1 146 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 146 1
rect -2 -2 146 -1
<< ptie >>
rect 0 1 144 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 144 1
rect 0 -3 144 -1
<< ntie >>
rect 0 81 144 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 144 81
rect 0 77 144 79
<< nmos >>
rect 32 11 34 30
rect 39 11 41 30
rect 49 11 51 30
rect 56 11 58 30
rect 72 11 74 30
rect 79 11 81 30
rect 89 11 91 30
rect 96 11 98 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 42 81 70
rect 89 42 91 70
rect 99 42 101 70
rect 109 42 111 70
rect 119 42 121 70
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 43 35 45 37
rect 59 35 61 37
rect 70 35 72 37
rect 83 35 85 37
rect 99 35 101 37
rect 107 35 109 37
rect 123 35 125 37
<< ndifct0 >>
rect 64 12 66 13
rect 101 20 103 22
rect 101 13 103 15
<< ndifct1 >>
rect 44 19 46 21
rect 64 11 66 12
rect 84 19 86 21
rect 26 9 28 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
<< pdifct0 >>
rect 4 60 6 62
rect 4 53 6 55
rect 24 60 26 62
rect 44 60 46 62
rect 64 59 66 61
rect 64 52 66 54
rect 74 66 76 68
rect 74 59 76 61
rect 84 58 86 60
rect 84 51 86 53
rect 94 66 96 68
rect 94 59 96 61
rect 104 58 106 60
rect 104 51 106 53
rect 114 66 116 68
rect 114 59 116 61
rect 124 51 126 53
rect 124 44 126 46
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
rect 34 51 36 53
rect 54 51 56 53
<< alu0 >>
rect 72 66 74 68
rect 76 66 78 68
rect 2 62 67 63
rect 2 60 4 62
rect 6 60 24 62
rect 26 60 44 62
rect 46 61 67 62
rect 46 60 64 61
rect 2 59 64 60
rect 66 59 67 61
rect 2 55 7 59
rect 2 53 4 55
rect 6 53 7 55
rect 63 54 67 59
rect 72 61 78 66
rect 92 66 94 68
rect 96 66 98 68
rect 72 59 74 61
rect 76 59 78 61
rect 72 58 78 59
rect 83 60 87 62
rect 83 58 84 60
rect 86 58 87 60
rect 92 61 98 66
rect 112 66 114 68
rect 116 66 118 68
rect 92 59 94 61
rect 96 59 98 61
rect 92 58 98 59
rect 103 60 107 62
rect 103 58 104 60
rect 106 58 107 60
rect 112 61 118 66
rect 112 59 114 61
rect 116 59 118 61
rect 112 58 118 59
rect 83 54 87 58
rect 103 54 107 58
rect 2 51 7 53
rect 63 52 64 54
rect 66 53 128 54
rect 66 52 84 53
rect 63 51 84 52
rect 86 51 104 53
rect 106 51 124 53
rect 126 51 128 53
rect 63 50 128 51
rect 122 46 128 50
rect 122 44 124 46
rect 126 44 128 46
rect 122 43 128 44
rect 99 22 105 23
rect 99 20 101 22
rect 103 20 105 22
rect 99 15 105 20
rect 62 13 68 14
rect 62 12 64 13
rect 66 12 68 13
rect 99 13 101 15
rect 103 13 105 15
rect 99 12 105 13
<< labels >>
rlabel alu0 4 57 4 57 6 n3
rlabel alu0 65 56 65 56 6 n3
rlabel alu0 34 61 34 61 6 n3
rlabel alu0 105 56 105 56 6 n3
rlabel alu0 85 56 85 56 6 n3
rlabel alu0 125 48 125 48 6 n3
rlabel alu0 95 52 95 52 6 n3
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 b2
rlabel polyct1 12 36 12 36 6 b2
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 b2
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 b2
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 44 32 44 32 6 b2
rlabel alu1 28 40 28 40 6 b1
rlabel alu1 36 44 36 44 6 b1
rlabel alu1 44 44 44 44 6 b1
rlabel alu1 52 44 52 44 6 b1
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 72 6 72 6 6 vss
rlabel alu1 60 20 60 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 68 28 68 28 6 a1
rlabel alu1 76 20 76 20 6 z
rlabel alu1 84 20 84 20 6 z
rlabel alu1 84 32 84 32 6 a2
rlabel alu1 60 40 60 40 6 b1
rlabel alu1 76 44 76 44 6 a1
rlabel alu1 84 44 84 44 6 a1
rlabel alu1 72 74 72 74 6 vdd
rlabel alu1 100 28 100 28 6 a2
rlabel alu1 108 28 108 28 6 a2
rlabel alu1 92 28 92 28 6 a2
rlabel alu1 100 40 100 40 6 a1
rlabel polyct1 108 36 108 36 6 a1
rlabel alu1 92 44 92 44 6 a1
rlabel alu1 116 28 116 28 6 a2
rlabel alu1 124 28 124 28 6 a2
<< end >>
