magic
tech scmos
timestamp 1199201905
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 9 33 11 43
rect 19 40 21 43
rect 29 40 31 43
rect 19 38 25 40
rect 19 36 21 38
rect 23 36 25 38
rect 19 34 25 36
rect 29 38 35 40
rect 29 36 31 38
rect 33 36 35 38
rect 29 34 35 36
rect 39 39 41 43
rect 39 37 47 39
rect 39 35 43 37
rect 45 35 47 37
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 23 30 25 34
rect 31 30 33 34
rect 39 33 47 35
rect 39 30 41 33
rect 9 27 15 29
rect 13 24 15 27
rect 13 12 15 17
rect 23 9 25 14
rect 31 9 33 14
rect 39 9 41 14
<< ndif >>
rect 18 24 23 30
rect 4 17 13 24
rect 15 21 23 24
rect 15 19 18 21
rect 20 19 23 21
rect 15 17 23 19
rect 4 11 11 17
rect 18 14 23 17
rect 25 14 31 30
rect 33 14 39 30
rect 41 18 48 30
rect 41 16 44 18
rect 46 16 48 18
rect 41 14 48 16
rect 4 9 7 11
rect 9 9 11 11
rect 4 7 11 9
<< pdif >>
rect 4 64 9 70
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 54 9 60
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 43 9 50
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 43 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 43 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 43 39 52
rect 41 68 48 70
rect 41 66 44 68
rect 46 66 48 68
rect 41 61 48 66
rect 41 59 44 61
rect 46 59 48 61
rect 41 43 48 59
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 62 8 63
rect 2 60 4 62
rect 6 60 8 62
rect 2 54 8 60
rect 2 52 4 54
rect 6 52 8 54
rect 2 51 8 52
rect 2 22 6 51
rect 10 41 24 47
rect 41 46 47 54
rect 17 38 24 41
rect 17 36 21 38
rect 23 36 24 38
rect 17 34 24 36
rect 29 42 47 46
rect 29 38 35 42
rect 29 36 31 38
rect 33 36 35 38
rect 29 35 35 36
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 31 47 35
rect 10 29 11 30
rect 13 29 30 30
rect 10 26 30 29
rect 2 21 22 22
rect 2 19 18 21
rect 20 19 22 21
rect 2 17 22 19
rect 26 17 30 26
rect 34 25 47 31
rect -2 11 58 12
rect -2 9 7 11
rect 9 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 13 17 15 24
rect 23 14 25 30
rect 31 14 33 30
rect 39 14 41 30
<< pmos >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
<< polyct0 >>
rect 11 30 13 31
<< polyct1 >>
rect 21 36 23 38
rect 31 36 33 38
rect 43 35 45 37
rect 11 29 13 30
<< ndifct0 >>
rect 44 16 46 18
<< ndifct1 >>
rect 18 19 20 21
rect 7 9 9 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 14 59 16 61
rect 14 52 16 54
rect 24 66 26 68
rect 24 59 26 61
rect 34 59 36 61
rect 34 52 36 54
rect 44 66 46 68
rect 44 59 46 61
<< pdifct1 >>
rect 4 60 6 62
rect 4 52 6 54
<< alu0 >>
rect 22 66 24 68
rect 26 66 28 68
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 61 28 66
rect 42 66 44 68
rect 46 66 48 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 33 61 37 63
rect 33 59 34 61
rect 36 59 37 61
rect 33 54 37 59
rect 42 61 48 66
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 13 52 14 54
rect 16 52 34 54
rect 36 52 37 54
rect 13 50 37 52
rect 10 31 14 33
rect 10 30 11 31
rect 13 30 14 31
rect 43 18 47 20
rect 43 16 44 18
rect 46 16 47 18
rect 43 12 47 16
<< labels >>
rlabel alu0 15 56 15 56 6 n3
rlabel alu0 35 56 35 56 6 n3
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 40 20 40 6 a3
rlabel alu1 12 44 12 44 6 a3
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 20 28 20 6 b
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 36 44 36 44 6 a2
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 44 48 44 48 6 a2
<< end >>
