magic
tech scmos
timestamp 1199202696
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 90 60 92 65
rect 100 60 102 65
rect 9 39 11 43
rect 19 39 21 43
rect 29 39 31 43
rect 39 39 41 43
rect 49 39 51 43
rect 59 39 61 43
rect 69 39 71 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 33 39
rect 19 35 27 37
rect 29 35 33 37
rect 19 33 33 35
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 37 51 39
rect 38 35 43 37
rect 45 35 51 37
rect 38 33 51 35
rect 55 37 71 39
rect 79 39 81 43
rect 90 39 92 43
rect 100 39 102 43
rect 79 37 92 39
rect 96 37 102 39
rect 55 35 59 37
rect 61 35 63 37
rect 55 33 63 35
rect 81 35 83 37
rect 85 35 87 37
rect 81 33 87 35
rect 96 35 98 37
rect 100 35 102 37
rect 96 33 102 35
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 12 11 14 16
rect 19 11 21 16
rect 31 6 33 11
rect 38 6 40 11
rect 48 6 50 11
rect 55 6 57 11
<< ndif >>
rect 5 28 12 30
rect 5 26 7 28
rect 9 26 12 28
rect 5 21 12 26
rect 5 19 7 21
rect 9 19 12 21
rect 5 16 12 19
rect 14 16 19 30
rect 21 16 31 30
rect 23 11 31 16
rect 33 11 38 30
rect 40 21 48 30
rect 40 19 43 21
rect 45 19 48 21
rect 40 11 48 19
rect 50 11 55 30
rect 57 11 66 30
rect 23 9 25 11
rect 27 9 29 11
rect 23 7 29 9
rect 59 9 61 11
rect 63 9 66 11
rect 59 7 66 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 43 9 59
rect 11 60 19 70
rect 11 58 14 60
rect 16 58 19 60
rect 11 53 19 58
rect 11 51 14 53
rect 16 51 19 53
rect 11 43 19 51
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 43 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 43 39 51
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 61 49 66
rect 41 59 44 61
rect 46 59 49 61
rect 41 43 49 59
rect 51 60 59 70
rect 51 58 54 60
rect 56 58 59 60
rect 51 53 59 58
rect 51 51 54 53
rect 56 51 59 53
rect 51 43 59 51
rect 61 68 69 70
rect 61 66 64 68
rect 66 66 69 68
rect 61 61 69 66
rect 61 59 64 61
rect 66 59 69 61
rect 61 43 69 59
rect 71 61 79 70
rect 71 59 74 61
rect 76 59 79 61
rect 71 53 79 59
rect 71 51 74 53
rect 76 51 79 53
rect 71 43 79 51
rect 81 68 88 70
rect 81 66 84 68
rect 86 66 88 68
rect 81 61 88 66
rect 81 59 84 61
rect 86 60 88 61
rect 86 59 90 60
rect 81 43 90 59
rect 92 53 100 60
rect 92 51 95 53
rect 97 51 100 53
rect 92 43 100 51
rect 102 58 110 60
rect 102 56 105 58
rect 107 56 110 58
rect 102 50 110 56
rect 102 48 105 50
rect 107 48 110 50
rect 102 43 110 48
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 68 114 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 73 61 78 63
rect 73 59 74 61
rect 76 59 78 61
rect 73 54 78 59
rect 2 53 99 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 51 54 53
rect 56 51 74 53
rect 76 51 95 53
rect 97 51 99 53
rect 2 50 99 51
rect 2 29 6 50
rect 25 42 97 46
rect 10 37 20 39
rect 10 35 11 37
rect 13 35 20 37
rect 10 33 20 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 16 30 20 33
rect 41 30 47 35
rect 57 37 63 42
rect 93 38 97 42
rect 57 35 59 37
rect 61 35 63 37
rect 57 34 63 35
rect 81 37 87 38
rect 81 35 83 37
rect 85 35 87 37
rect 81 30 87 35
rect 93 37 103 38
rect 93 35 98 37
rect 100 35 103 37
rect 93 34 103 35
rect 2 28 11 29
rect 2 26 7 28
rect 9 26 11 28
rect 16 26 87 30
rect 2 25 11 26
rect 7 22 11 25
rect 7 21 47 22
rect 9 19 43 21
rect 45 19 47 21
rect 7 18 47 19
rect -2 11 114 12
rect -2 9 25 11
rect 27 9 61 11
rect 63 9 114 11
rect -2 1 114 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 12 16 14 30
rect 19 16 21 30
rect 31 11 33 30
rect 38 11 40 30
rect 48 11 50 30
rect 55 11 57 30
<< pmos >>
rect 9 43 11 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
rect 49 43 51 70
rect 59 43 61 70
rect 69 43 71 70
rect 79 43 81 70
rect 90 43 92 60
rect 100 43 102 60
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 43 35 45 37
rect 59 35 61 37
rect 83 35 85 37
rect 98 35 100 37
<< ndifct1 >>
rect 7 26 9 28
rect 7 19 9 21
rect 43 19 45 21
rect 25 9 27 11
rect 61 9 63 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 58 16 60
rect 24 66 26 68
rect 24 59 26 61
rect 44 66 46 68
rect 44 59 46 61
rect 54 58 56 60
rect 64 66 66 68
rect 64 59 66 61
rect 84 66 86 68
rect 84 59 86 61
rect 105 56 107 58
rect 105 48 107 50
<< pdifct1 >>
rect 14 51 16 53
rect 34 59 36 61
rect 34 51 36 53
rect 54 51 56 53
rect 74 59 76 61
rect 74 51 76 53
rect 95 51 97 53
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 60 17 62
rect 13 58 14 60
rect 16 58 17 60
rect 22 61 28 66
rect 42 66 44 68
rect 46 66 48 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 13 54 17 58
rect 42 61 48 66
rect 62 66 64 68
rect 66 66 68 68
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 53 60 57 62
rect 53 58 54 60
rect 56 58 57 60
rect 62 61 68 66
rect 82 66 84 68
rect 86 66 88 68
rect 62 59 64 61
rect 66 59 68 61
rect 62 58 68 59
rect 53 54 57 58
rect 82 61 88 66
rect 82 59 84 61
rect 86 59 88 61
rect 82 58 88 59
rect 104 58 108 68
rect 104 56 105 58
rect 107 56 108 58
rect 104 50 108 56
rect 104 48 105 50
rect 107 48 108 50
rect 104 46 108 48
rect 5 18 7 25
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 b
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 b
rlabel polyct1 28 36 28 36 6 a
rlabel alu1 28 40 28 40 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 56 6 56 6 6 vss
rlabel ndifct1 44 20 44 20 6 z
rlabel alu1 52 28 52 28 6 b
rlabel alu1 60 28 60 28 6 b
rlabel alu1 44 32 44 32 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 52 44 52 44 6 a
rlabel alu1 60 40 60 40 6 a
rlabel alu1 52 52 52 52 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 56 74 56 74 6 vdd
rlabel alu1 68 28 68 28 6 b
rlabel alu1 76 28 76 28 6 b
rlabel alu1 84 32 84 32 6 b
rlabel alu1 68 44 68 44 6 a
rlabel alu1 76 44 76 44 6 a
rlabel alu1 84 44 84 44 6 a
rlabel alu1 84 52 84 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 76 56 76 56 6 z
rlabel alu1 92 44 92 44 6 a
rlabel alu1 100 36 100 36 6 a
rlabel alu1 92 52 92 52 6 z
<< end >>
