magic
tech scmos
timestamp 1199203235
<< ab >>
rect 0 0 104 80
<< nwell >>
rect -5 36 109 88
<< pwell >>
rect -5 -8 109 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 66 31 71
rect 39 66 41 71
rect 49 66 51 71
rect 56 66 58 71
rect 66 66 68 71
rect 73 66 75 71
rect 83 60 85 65
rect 90 60 92 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 9 37 41 39
rect 45 37 51 39
rect 9 30 11 37
rect 19 30 21 37
rect 29 35 33 37
rect 35 35 37 37
rect 29 33 37 35
rect 45 35 47 37
rect 49 35 51 37
rect 45 33 51 35
rect 56 39 58 42
rect 66 39 68 42
rect 56 37 68 39
rect 56 35 64 37
rect 66 35 68 37
rect 56 33 68 35
rect 73 39 75 42
rect 83 39 85 42
rect 90 39 92 42
rect 73 37 85 39
rect 89 37 95 39
rect 29 30 31 33
rect 9 13 11 18
rect 46 28 48 33
rect 56 28 58 33
rect 73 31 75 37
rect 89 35 91 37
rect 93 35 95 37
rect 89 33 95 35
rect 72 29 78 31
rect 72 27 74 29
rect 76 27 78 29
rect 72 25 78 27
rect 19 6 21 10
rect 29 6 31 10
rect 46 6 48 10
rect 56 6 58 10
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 18 9 24
rect 11 22 19 30
rect 11 20 14 22
rect 16 20 19 22
rect 11 18 19 20
rect 13 10 19 18
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 21 29 26
rect 21 19 24 21
rect 26 19 29 21
rect 21 10 29 19
rect 31 28 44 30
rect 31 15 46 28
rect 31 13 34 15
rect 36 13 46 15
rect 31 10 46 13
rect 48 20 56 28
rect 48 18 51 20
rect 53 18 56 20
rect 48 10 56 18
rect 58 21 65 28
rect 58 19 61 21
rect 63 19 65 21
rect 58 14 65 19
rect 58 12 61 14
rect 63 12 65 14
rect 58 10 65 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 66 27 70
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 42 29 62
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 42 39 52
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 56 49 62
rect 41 54 44 56
rect 46 54 49 56
rect 41 42 49 54
rect 51 42 56 66
rect 58 55 66 66
rect 58 53 61 55
rect 63 53 66 55
rect 58 47 66 53
rect 58 45 61 47
rect 63 45 66 47
rect 58 42 66 45
rect 68 42 73 66
rect 75 60 81 66
rect 75 58 83 60
rect 75 56 78 58
rect 80 56 83 58
rect 75 42 83 56
rect 85 42 90 60
rect 92 55 97 60
rect 92 53 99 55
rect 92 51 95 53
rect 97 51 99 53
rect 92 46 99 51
rect 92 44 95 46
rect 97 44 99 46
rect 92 42 99 44
<< alu1 >>
rect -2 81 106 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 106 81
rect -2 68 106 79
rect 33 61 39 63
rect 33 59 34 61
rect 36 59 39 61
rect 33 54 39 59
rect 9 52 14 54
rect 16 52 34 54
rect 36 52 39 54
rect 9 50 39 52
rect 18 39 22 50
rect 2 38 22 39
rect 2 34 27 38
rect 45 37 55 38
rect 45 35 47 37
rect 49 35 55 37
rect 45 34 55 35
rect 62 37 95 38
rect 62 35 64 37
rect 66 35 91 37
rect 93 35 95 37
rect 62 34 95 35
rect 2 28 7 34
rect 2 26 4 28
rect 6 26 7 28
rect 2 24 7 26
rect 23 28 27 34
rect 23 26 24 28
rect 26 26 27 28
rect 23 21 27 26
rect 49 30 55 34
rect 49 29 78 30
rect 49 27 74 29
rect 76 27 78 29
rect 49 26 78 27
rect 89 26 95 34
rect 23 19 24 21
rect 26 19 27 21
rect 23 17 27 19
rect 74 17 78 26
rect -2 1 106 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 106 1
rect -2 -2 106 -1
<< ptie >>
rect 0 1 104 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 104 1
rect 0 -3 104 -1
<< ntie >>
rect 0 81 104 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 104 81
rect 0 77 104 79
<< nmos >>
rect 9 18 11 30
rect 19 10 21 30
rect 29 10 31 30
rect 46 10 48 28
rect 56 10 58 28
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 66
rect 39 42 41 66
rect 49 42 51 66
rect 56 42 58 66
rect 66 42 68 66
rect 73 42 75 66
rect 83 42 85 60
rect 90 42 92 60
<< polyct0 >>
rect 33 35 35 37
<< polyct1 >>
rect 47 35 49 37
rect 64 35 66 37
rect 91 35 93 37
rect 74 27 76 29
<< ndifct0 >>
rect 14 20 16 22
rect 34 13 36 15
rect 51 18 53 20
rect 61 19 63 21
rect 61 12 63 14
<< ndifct1 >>
rect 4 26 6 28
rect 24 26 26 28
rect 24 19 26 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 59 16 61
rect 24 62 26 64
rect 44 62 46 64
rect 44 54 46 56
rect 61 53 63 55
rect 61 45 63 47
rect 78 56 80 58
rect 95 51 97 53
rect 95 44 97 46
<< pdifct1 >>
rect 14 52 16 54
rect 34 59 36 61
rect 34 52 36 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 23 64 27 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 23 62 24 64
rect 26 62 27 64
rect 43 64 47 68
rect 23 60 27 62
rect 13 54 17 59
rect 43 62 44 64
rect 46 62 47 64
rect 43 56 47 62
rect 77 58 81 68
rect 43 54 44 56
rect 46 54 47 56
rect 43 52 47 54
rect 60 55 64 57
rect 60 53 61 55
rect 63 53 64 55
rect 77 56 78 58
rect 80 56 81 58
rect 77 54 81 56
rect 60 47 64 53
rect 60 46 61 47
rect 37 45 61 46
rect 63 46 64 47
rect 94 53 98 55
rect 94 51 95 53
rect 97 51 98 53
rect 94 46 98 51
rect 63 45 95 46
rect 37 44 95 45
rect 97 44 98 46
rect 37 42 98 44
rect 37 38 41 42
rect 31 37 41 38
rect 31 35 33 37
rect 35 35 41 37
rect 31 34 41 35
rect 13 22 17 24
rect 13 20 14 22
rect 16 20 17 22
rect 13 12 17 20
rect 37 26 41 34
rect 37 22 45 26
rect 41 21 45 22
rect 59 21 65 22
rect 41 20 55 21
rect 41 18 51 20
rect 53 18 55 20
rect 41 17 55 18
rect 59 19 61 21
rect 63 19 65 21
rect 33 15 37 17
rect 33 13 34 15
rect 36 13 37 15
rect 33 12 37 13
rect 59 14 65 19
rect 59 12 61 14
rect 63 12 65 14
<< labels >>
rlabel alu0 36 36 36 36 6 zn
rlabel alu0 48 19 48 19 6 zn
rlabel alu0 62 49 62 49 6 zn
rlabel alu0 96 48 96 48 6 zn
rlabel alu1 12 36 12 36 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 52 6 52 6 6 vss
rlabel alu1 76 20 76 20 6 a
rlabel alu1 52 32 52 32 6 a
rlabel alu1 68 36 68 36 6 b
rlabel alu1 76 36 76 36 6 b
rlabel alu1 68 28 68 28 6 a
rlabel alu1 60 28 60 28 6 a
rlabel alu1 52 74 52 74 6 vdd
rlabel alu1 84 36 84 36 6 b
rlabel alu1 92 32 92 32 6 b
<< end >>
