magic
tech scmos
timestamp 1199542317
<< ab >>
rect 0 0 140 100
<< nwell >>
rect -5 48 145 105
<< pwell >>
rect -5 -5 145 48
<< poly >>
rect 25 94 27 98
rect 37 94 39 98
rect 49 94 51 98
rect 57 94 59 98
rect 69 94 71 98
rect 81 94 83 98
rect 89 94 91 98
rect 113 94 115 98
rect 125 94 127 98
rect 13 70 15 74
rect 13 53 15 56
rect 5 51 15 53
rect 5 49 7 51
rect 9 49 15 51
rect 5 47 15 49
rect 13 37 15 47
rect 25 53 27 75
rect 37 73 39 76
rect 31 71 39 73
rect 31 69 33 71
rect 35 69 39 71
rect 31 67 39 69
rect 25 51 33 53
rect 25 49 29 51
rect 31 49 33 51
rect 25 47 33 49
rect 13 25 15 29
rect 25 23 27 47
rect 37 41 39 67
rect 49 63 51 75
rect 45 61 51 63
rect 45 59 47 61
rect 49 59 51 61
rect 45 57 51 59
rect 47 51 53 53
rect 57 51 59 75
rect 69 73 71 76
rect 81 73 83 76
rect 47 49 49 51
rect 51 49 59 51
rect 47 47 53 49
rect 37 39 51 41
rect 31 31 39 33
rect 31 29 33 31
rect 35 29 39 31
rect 31 27 39 29
rect 37 23 39 27
rect 49 23 51 39
rect 57 23 59 49
rect 67 71 71 73
rect 77 71 83 73
rect 67 33 69 71
rect 77 53 79 71
rect 89 63 91 76
rect 101 69 103 73
rect 83 61 91 63
rect 83 59 85 61
rect 87 59 91 61
rect 83 57 91 59
rect 73 51 79 53
rect 101 51 103 55
rect 73 49 75 51
rect 77 49 103 51
rect 73 47 79 49
rect 77 39 79 47
rect 63 31 69 33
rect 63 29 65 31
rect 67 29 69 31
rect 63 27 69 29
rect 73 37 79 39
rect 83 41 91 43
rect 83 39 85 41
rect 87 39 91 41
rect 83 37 91 39
rect 73 23 75 37
rect 79 31 85 33
rect 79 29 81 31
rect 83 29 85 31
rect 79 27 85 29
rect 69 21 75 23
rect 69 18 71 21
rect 81 19 83 27
rect 89 19 91 37
rect 101 35 103 49
rect 113 43 115 55
rect 109 41 115 43
rect 125 41 127 55
rect 109 39 111 41
rect 113 39 127 41
rect 109 37 115 39
rect 113 34 115 37
rect 125 35 127 39
rect 101 25 103 29
rect 25 7 27 11
rect 37 7 39 11
rect 49 7 51 11
rect 57 7 59 11
rect 113 11 115 15
rect 125 11 127 15
rect 69 2 71 6
rect 81 3 83 7
rect 89 3 91 7
<< ndif >>
rect 5 29 13 37
rect 15 33 23 37
rect 15 31 19 33
rect 21 31 23 33
rect 15 29 23 31
rect 5 21 11 29
rect 41 31 47 33
rect 41 29 43 31
rect 45 29 47 31
rect 41 23 47 29
rect 5 19 7 21
rect 9 19 11 21
rect 5 17 11 19
rect 17 21 25 23
rect 17 19 19 21
rect 21 19 25 21
rect 17 11 25 19
rect 27 11 37 23
rect 39 11 49 23
rect 51 11 57 23
rect 59 21 67 23
rect 59 19 63 21
rect 65 19 67 21
rect 59 18 67 19
rect 93 33 101 35
rect 93 31 95 33
rect 97 31 101 33
rect 93 29 101 31
rect 103 34 108 35
rect 120 34 125 35
rect 103 29 113 34
rect 93 21 99 23
rect 93 19 95 21
rect 97 19 99 21
rect 76 18 81 19
rect 59 11 69 18
rect 61 6 69 11
rect 71 11 81 18
rect 71 9 75 11
rect 77 9 81 11
rect 71 7 81 9
rect 83 7 89 19
rect 91 7 99 19
rect 105 15 113 29
rect 115 31 125 34
rect 115 29 119 31
rect 121 29 125 31
rect 115 21 125 29
rect 115 19 119 21
rect 121 19 125 21
rect 115 15 125 19
rect 127 31 135 35
rect 127 29 131 31
rect 133 29 135 31
rect 127 21 135 29
rect 127 19 131 21
rect 133 19 135 21
rect 127 15 135 19
rect 105 11 111 15
rect 105 9 107 11
rect 109 9 111 11
rect 105 7 111 9
rect 71 6 78 7
<< pdif >>
rect 105 94 111 95
rect 129 94 135 95
rect 5 81 11 83
rect 5 79 7 81
rect 9 79 11 81
rect 5 70 11 79
rect 17 81 25 94
rect 17 79 19 81
rect 21 79 25 81
rect 17 75 25 79
rect 27 76 37 94
rect 39 76 49 94
rect 27 75 32 76
rect 5 56 13 70
rect 15 61 23 70
rect 15 59 19 61
rect 21 59 23 61
rect 15 56 23 59
rect 41 75 49 76
rect 51 75 57 94
rect 59 81 69 94
rect 59 79 63 81
rect 65 79 69 81
rect 59 76 69 79
rect 71 91 81 94
rect 71 89 75 91
rect 77 89 81 91
rect 71 76 81 89
rect 83 76 89 94
rect 91 81 99 94
rect 91 79 95 81
rect 97 79 99 81
rect 91 76 99 79
rect 105 93 113 94
rect 105 91 107 93
rect 109 91 113 93
rect 59 75 64 76
rect 41 71 47 75
rect 41 69 43 71
rect 45 69 47 71
rect 41 67 47 69
rect 105 69 113 91
rect 93 61 101 69
rect 93 59 95 61
rect 97 59 101 61
rect 93 55 101 59
rect 103 55 113 69
rect 115 81 125 94
rect 115 79 119 81
rect 121 79 125 81
rect 115 71 125 79
rect 115 69 119 71
rect 121 69 125 71
rect 115 61 125 69
rect 115 59 119 61
rect 121 59 125 61
rect 115 55 125 59
rect 127 93 135 94
rect 127 91 131 93
rect 133 91 135 93
rect 127 81 135 91
rect 127 79 131 81
rect 133 79 135 81
rect 127 71 135 79
rect 127 69 131 71
rect 133 69 135 71
rect 127 61 135 69
rect 127 59 131 61
rect 133 59 135 61
rect 127 55 135 59
<< alu1 >>
rect -2 93 142 100
rect -2 91 107 93
rect 109 91 131 93
rect 133 91 142 93
rect -2 89 75 91
rect 77 89 142 91
rect -2 88 142 89
rect 6 81 10 88
rect 6 79 7 81
rect 9 79 10 81
rect 6 77 10 79
rect 17 81 67 82
rect 17 79 19 81
rect 21 79 63 81
rect 65 79 67 81
rect 17 78 67 79
rect 94 81 98 83
rect 94 79 95 81
rect 97 79 98 81
rect 8 72 12 73
rect 94 72 98 79
rect 118 81 122 83
rect 118 79 119 81
rect 121 79 122 81
rect 8 71 37 72
rect 8 69 33 71
rect 35 69 37 71
rect 8 68 37 69
rect 41 71 112 72
rect 41 69 43 71
rect 45 69 112 71
rect 41 68 112 69
rect 8 52 12 68
rect 5 51 12 52
rect 5 49 7 51
rect 9 49 12 51
rect 5 48 12 49
rect 8 27 12 48
rect 18 62 22 63
rect 18 61 51 62
rect 18 59 19 61
rect 21 59 47 61
rect 49 59 51 61
rect 18 58 51 59
rect 18 33 22 58
rect 28 51 32 53
rect 28 49 29 51
rect 31 49 32 51
rect 28 41 32 49
rect 39 51 53 52
rect 39 49 49 51
rect 51 49 53 51
rect 39 48 53 49
rect 58 42 62 68
rect 18 31 19 33
rect 21 32 22 33
rect 52 38 62 42
rect 68 52 72 63
rect 84 62 88 63
rect 77 61 88 62
rect 77 59 85 61
rect 87 59 88 61
rect 77 58 88 59
rect 93 61 102 62
rect 93 59 95 61
rect 97 59 102 61
rect 93 58 102 59
rect 84 52 88 58
rect 68 51 79 52
rect 68 49 75 51
rect 77 49 79 51
rect 68 48 79 49
rect 84 48 93 52
rect 52 32 56 38
rect 68 37 72 48
rect 84 42 88 48
rect 77 41 88 42
rect 77 39 85 41
rect 87 39 88 41
rect 77 38 88 39
rect 84 37 88 38
rect 98 36 102 58
rect 94 33 102 36
rect 94 32 95 33
rect 21 31 37 32
rect 18 29 33 31
rect 35 29 37 31
rect 18 28 37 29
rect 41 31 56 32
rect 41 29 43 31
rect 45 29 56 31
rect 41 28 56 29
rect 63 31 95 32
rect 97 32 102 33
rect 108 42 112 68
rect 118 71 122 79
rect 118 69 119 71
rect 121 69 122 71
rect 118 61 122 69
rect 118 59 119 61
rect 121 59 122 61
rect 118 52 122 59
rect 130 81 134 88
rect 130 79 131 81
rect 133 79 134 81
rect 130 71 134 79
rect 130 69 131 71
rect 133 69 134 71
rect 130 61 134 69
rect 130 59 131 61
rect 133 59 134 61
rect 130 57 134 59
rect 118 47 124 52
rect 120 42 124 47
rect 108 41 115 42
rect 108 39 111 41
rect 113 39 115 41
rect 108 38 115 39
rect 120 38 133 42
rect 97 31 98 32
rect 63 29 65 31
rect 67 29 81 31
rect 83 29 98 31
rect 63 28 98 29
rect 6 21 10 23
rect 108 22 112 38
rect 120 33 124 38
rect 6 19 7 21
rect 9 19 10 21
rect 6 12 10 19
rect 17 21 67 22
rect 17 19 19 21
rect 21 19 63 21
rect 65 19 67 21
rect 17 18 67 19
rect 93 21 112 22
rect 93 19 95 21
rect 97 19 112 21
rect 93 18 112 19
rect 118 31 124 33
rect 118 29 119 31
rect 121 29 124 31
rect 118 28 124 29
rect 130 31 134 33
rect 130 29 131 31
rect 133 29 134 31
rect 118 21 122 28
rect 118 19 119 21
rect 121 19 122 21
rect 118 17 122 19
rect 130 21 134 29
rect 130 19 131 21
rect 133 19 134 21
rect 130 12 134 19
rect -2 11 142 12
rect -2 9 75 11
rect 77 9 107 11
rect 109 9 142 11
rect -2 7 142 9
rect -2 5 119 7
rect 121 5 142 7
rect -2 0 142 5
<< ptie >>
rect 117 7 128 9
rect 117 5 119 7
rect 121 5 128 7
rect 117 3 128 5
<< nmos >>
rect 13 29 15 37
rect 25 11 27 23
rect 37 11 39 23
rect 49 11 51 23
rect 57 11 59 23
rect 101 29 103 35
rect 69 6 71 18
rect 81 7 83 19
rect 89 7 91 19
rect 113 15 115 34
rect 125 15 127 35
<< pmos >>
rect 25 75 27 94
rect 37 76 39 94
rect 13 56 15 70
rect 49 75 51 94
rect 57 75 59 94
rect 69 76 71 94
rect 81 76 83 94
rect 89 76 91 94
rect 101 55 103 69
rect 113 55 115 94
rect 125 55 127 94
<< polyct1 >>
rect 7 49 9 51
rect 33 69 35 71
rect 29 49 31 51
rect 47 59 49 61
rect 49 49 51 51
rect 33 29 35 31
rect 85 59 87 61
rect 75 49 77 51
rect 65 29 67 31
rect 85 39 87 41
rect 81 29 83 31
rect 111 39 113 41
<< ndifct1 >>
rect 19 31 21 33
rect 43 29 45 31
rect 7 19 9 21
rect 19 19 21 21
rect 63 19 65 21
rect 95 31 97 33
rect 95 19 97 21
rect 75 9 77 11
rect 119 29 121 31
rect 119 19 121 21
rect 131 29 133 31
rect 131 19 133 21
rect 107 9 109 11
<< ptiect1 >>
rect 119 5 121 7
<< pdifct1 >>
rect 7 79 9 81
rect 19 79 21 81
rect 19 59 21 61
rect 63 79 65 81
rect 75 89 77 91
rect 95 79 97 81
rect 107 91 109 93
rect 43 69 45 71
rect 95 59 97 61
rect 119 79 121 81
rect 119 69 121 71
rect 119 59 121 61
rect 131 91 133 93
rect 131 79 133 81
rect 131 69 133 71
rect 131 59 133 61
<< labels >>
rlabel alu1 10 50 10 50 6 cmd1
rlabel alu1 20 70 20 70 6 cmd1
rlabel polyct1 30 50 30 50 6 i2
rlabel polyct1 50 50 50 50 6 i1
rlabel alu1 30 70 30 70 6 cmd1
rlabel alu1 70 6 70 6 6 vss
rlabel alu1 80 40 80 40 6 i0
rlabel alu1 70 50 70 50 6 cmd0
rlabel alu1 80 60 80 60 6 i0
rlabel alu1 70 94 70 94 6 vdd
rlabel alu1 90 50 90 50 6 i0
rlabel alu1 120 25 120 25 6 q
rlabel alu1 130 40 130 40 6 q
rlabel alu1 120 65 120 65 6 q
<< end >>
