magic
tech scmos
timestamp 1199202557
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 10 66 12 71
rect 20 66 22 71
rect 32 60 34 65
rect 10 38 12 42
rect 20 38 22 42
rect 32 39 34 42
rect 9 36 15 38
rect 9 34 11 36
rect 13 34 15 36
rect 9 32 15 34
rect 19 36 25 38
rect 19 34 21 36
rect 23 34 25 36
rect 19 32 25 34
rect 32 37 39 39
rect 32 35 35 37
rect 37 35 39 37
rect 32 33 39 35
rect 12 29 14 32
rect 19 29 21 32
rect 33 29 35 33
rect 33 15 35 20
rect 12 6 14 10
rect 19 6 21 10
<< ndif >>
rect 7 22 12 29
rect 5 20 12 22
rect 5 18 7 20
rect 9 18 12 20
rect 5 16 12 18
rect 7 10 12 16
rect 14 10 19 29
rect 21 21 33 29
rect 21 19 27 21
rect 29 20 33 21
rect 35 27 42 29
rect 35 25 38 27
rect 40 25 42 27
rect 35 23 42 25
rect 35 20 40 23
rect 29 19 31 20
rect 21 14 31 19
rect 21 12 27 14
rect 29 12 31 14
rect 21 10 31 12
<< pdif >>
rect 2 63 10 66
rect 2 61 4 63
rect 6 61 10 63
rect 2 42 10 61
rect 12 62 20 66
rect 12 60 15 62
rect 17 60 20 62
rect 12 42 20 60
rect 22 63 30 66
rect 22 61 26 63
rect 28 61 30 63
rect 22 60 30 61
rect 22 42 32 60
rect 34 56 39 60
rect 34 54 41 56
rect 34 52 37 54
rect 39 52 41 54
rect 34 50 41 52
rect 34 42 39 50
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 10 62 19 63
rect 10 60 15 62
rect 17 60 19 62
rect 10 59 19 60
rect 10 55 14 59
rect 2 49 14 55
rect 2 21 6 49
rect 10 36 14 39
rect 10 34 11 36
rect 13 34 14 36
rect 10 29 14 34
rect 26 41 38 47
rect 34 37 38 41
rect 34 35 35 37
rect 37 35 38 37
rect 34 33 38 35
rect 10 25 22 29
rect 2 20 11 21
rect 2 18 7 20
rect 9 18 11 20
rect 2 17 11 18
rect 18 17 22 25
rect -2 1 50 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 12 10 14 29
rect 19 10 21 29
rect 33 20 35 29
<< pmos >>
rect 10 42 12 66
rect 20 42 22 66
rect 32 42 34 60
<< polyct0 >>
rect 21 34 23 36
<< polyct1 >>
rect 11 34 13 36
rect 35 35 37 37
<< ndifct0 >>
rect 27 19 29 21
rect 38 25 40 27
rect 27 12 29 14
<< ndifct1 >>
rect 7 18 9 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 4 61 6 63
rect 26 61 28 63
rect 37 52 39 54
<< pdifct1 >>
rect 15 60 17 62
<< alu0 >>
rect 3 63 7 68
rect 25 63 29 68
rect 3 61 4 63
rect 6 61 7 63
rect 3 59 7 61
rect 25 61 26 63
rect 28 61 29 63
rect 25 59 29 61
rect 18 54 41 55
rect 18 52 37 54
rect 39 52 41 54
rect 18 51 41 52
rect 18 37 22 51
rect 18 36 30 37
rect 18 34 21 36
rect 23 34 30 36
rect 18 33 30 34
rect 26 29 30 33
rect 26 27 42 29
rect 26 25 38 27
rect 40 25 42 27
rect 36 24 42 25
rect 25 21 31 22
rect 25 19 27 21
rect 29 19 31 21
rect 25 14 31 19
rect 25 12 27 14
rect 29 12 31 14
<< labels >>
rlabel alu0 24 35 24 35 6 an
rlabel alu0 34 27 34 27 6 an
rlabel alu0 29 53 29 53 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 b
rlabel alu1 12 32 12 32 6 b
rlabel alu1 12 56 12 56 6 z
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 44 28 44 6 a
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 36 40 36 40 6 a
<< end >>
