magic
tech scmos
timestamp 1199203121
<< ab >>
rect 0 0 88 80
<< nwell >>
rect -5 36 93 88
<< pwell >>
rect -5 -8 93 36
<< poly >>
rect 32 67 34 72
rect 39 67 41 72
rect 49 67 51 72
rect 56 67 58 72
rect 66 67 68 72
rect 73 67 75 72
rect 9 61 11 65
rect 22 63 24 67
rect 9 39 11 42
rect 22 39 24 42
rect 32 39 34 42
rect 39 39 41 42
rect 49 39 51 42
rect 56 39 58 42
rect 66 39 68 42
rect 9 37 24 39
rect 9 35 11 37
rect 13 35 24 37
rect 9 33 24 35
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 39 37 52 39
rect 56 37 68 39
rect 73 39 75 42
rect 73 37 79 39
rect 39 35 48 37
rect 50 35 52 37
rect 39 33 52 35
rect 59 35 61 37
rect 63 35 65 37
rect 59 33 65 35
rect 73 35 75 37
rect 77 35 79 37
rect 73 33 79 35
rect 10 30 12 33
rect 20 30 22 33
rect 30 30 32 33
rect 40 30 42 33
rect 50 30 52 33
rect 62 30 64 33
rect 10 8 12 13
rect 20 8 22 13
rect 30 8 32 13
rect 40 8 42 13
rect 50 8 52 13
rect 62 8 64 13
<< ndif >>
rect 5 22 10 30
rect 3 20 10 22
rect 3 18 5 20
rect 7 18 10 20
rect 3 16 10 18
rect 5 13 10 16
rect 12 28 20 30
rect 12 26 15 28
rect 17 26 20 28
rect 12 13 20 26
rect 22 20 30 30
rect 22 18 25 20
rect 27 18 30 20
rect 22 13 30 18
rect 32 17 40 30
rect 32 15 35 17
rect 37 15 40 17
rect 32 13 40 15
rect 42 20 50 30
rect 42 18 45 20
rect 47 18 50 20
rect 42 13 50 18
rect 52 13 62 30
rect 64 22 69 30
rect 64 20 71 22
rect 64 18 67 20
rect 69 18 71 20
rect 64 16 71 18
rect 64 13 69 16
rect 54 11 60 13
rect 54 9 56 11
rect 58 9 60 11
rect 54 7 60 9
<< pdif >>
rect 27 63 32 67
rect 14 61 22 63
rect 4 55 9 61
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 59 16 61
rect 18 59 22 61
rect 11 54 22 59
rect 11 52 16 54
rect 18 52 22 54
rect 11 42 22 52
rect 24 53 32 63
rect 24 51 27 53
rect 29 51 32 53
rect 24 46 32 51
rect 24 44 27 46
rect 29 44 32 46
rect 24 42 32 44
rect 34 42 39 67
rect 41 65 49 67
rect 41 63 44 65
rect 46 63 49 65
rect 41 42 49 63
rect 51 42 56 67
rect 58 61 66 67
rect 58 59 61 61
rect 63 59 66 61
rect 58 54 66 59
rect 58 52 61 54
rect 63 52 66 54
rect 58 42 66 52
rect 68 42 73 67
rect 75 65 82 67
rect 75 63 78 65
rect 80 63 82 65
rect 75 58 82 63
rect 75 56 78 58
rect 80 56 82 58
rect 75 42 82 56
<< alu1 >>
rect -2 81 90 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 90 81
rect -2 68 90 79
rect 58 61 64 63
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 58 59 61 61
rect 63 59 64 61
rect 58 54 64 59
rect 25 53 61 54
rect 25 51 27 53
rect 29 52 61 53
rect 63 52 71 54
rect 29 51 71 52
rect 2 47 7 51
rect 25 50 71 51
rect 25 47 30 50
rect 2 46 30 47
rect 2 44 4 46
rect 6 44 27 46
rect 29 44 30 46
rect 2 43 30 44
rect 18 42 30 43
rect 34 42 71 46
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 2 25 6 33
rect 18 29 22 42
rect 34 38 39 42
rect 29 37 39 38
rect 29 35 31 37
rect 33 35 39 37
rect 29 34 39 35
rect 46 37 55 38
rect 46 35 48 37
rect 50 35 55 37
rect 46 34 55 35
rect 73 37 79 38
rect 73 35 75 37
rect 77 35 79 37
rect 13 28 22 29
rect 13 26 15 28
rect 17 26 22 28
rect 49 30 55 34
rect 73 30 79 35
rect 13 25 22 26
rect 49 26 79 30
rect -2 11 90 12
rect -2 9 56 11
rect 58 9 90 11
rect -2 1 90 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 90 1
rect -2 -2 90 -1
<< ptie >>
rect 0 1 88 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 88 1
rect 0 -3 88 -1
<< ntie >>
rect 0 81 88 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 88 81
rect 0 77 88 79
<< nmos >>
rect 10 13 12 30
rect 20 13 22 30
rect 30 13 32 30
rect 40 13 42 30
rect 50 13 52 30
rect 62 13 64 30
<< pmos >>
rect 9 42 11 61
rect 22 42 24 63
rect 32 42 34 67
rect 39 42 41 67
rect 49 42 51 67
rect 56 42 58 67
rect 66 42 68 67
rect 73 42 75 67
<< polyct0 >>
rect 61 35 63 37
<< polyct1 >>
rect 11 35 13 37
rect 31 35 33 37
rect 48 35 50 37
rect 75 35 77 37
<< ndifct0 >>
rect 5 18 7 20
rect 25 18 27 20
rect 35 15 37 17
rect 45 18 47 20
rect 67 18 69 20
<< ndifct1 >>
rect 15 26 17 28
rect 56 9 58 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
<< pdifct0 >>
rect 16 59 18 61
rect 16 52 18 54
rect 44 63 46 65
rect 78 63 80 65
rect 78 56 80 58
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 27 51 29 53
rect 27 44 29 46
rect 61 59 63 61
rect 61 52 63 54
<< alu0 >>
rect 14 61 20 68
rect 43 65 47 68
rect 43 63 44 65
rect 46 63 47 65
rect 77 65 81 68
rect 77 63 78 65
rect 80 63 81 65
rect 43 61 47 63
rect 14 59 16 61
rect 18 59 20 61
rect 14 54 20 59
rect 77 58 81 63
rect 77 56 78 58
rect 80 56 81 58
rect 77 54 81 56
rect 14 52 16 54
rect 18 52 20 54
rect 14 51 20 52
rect 59 37 65 42
rect 59 35 61 37
rect 63 35 65 37
rect 59 34 65 35
rect 26 23 46 27
rect 26 21 30 23
rect 3 20 30 21
rect 3 18 5 20
rect 7 18 25 20
rect 27 18 30 20
rect 42 21 46 23
rect 42 20 71 21
rect 3 17 30 18
rect 34 17 38 19
rect 42 18 45 20
rect 47 18 67 20
rect 69 18 71 20
rect 42 17 71 18
rect 34 15 35 17
rect 37 15 38 17
rect 34 12 38 15
<< labels >>
rlabel alu0 16 19 16 19 6 n1
rlabel alu0 56 19 56 19 6 n1
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 32 4 32 6 b
rlabel alu1 4 52 4 52 6 z
rlabel alu1 20 36 20 36 6 z
rlabel alu1 36 36 36 36 6 a2
rlabel alu1 36 52 36 52 6 z
rlabel pdifct1 28 52 28 52 6 z
rlabel alu1 44 6 44 6 6 vss
rlabel alu1 52 32 52 32 6 a1
rlabel alu1 60 28 60 28 6 a1
rlabel alu1 52 44 52 44 6 a2
rlabel alu1 60 44 60 44 6 a2
rlabel alu1 44 44 44 44 6 a2
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 60 56 60 56 6 z
rlabel alu1 44 74 44 74 6 vdd
rlabel alu1 68 28 68 28 6 a1
rlabel alu1 76 32 76 32 6 a1
rlabel alu1 68 44 68 44 6 a2
rlabel alu1 68 52 68 52 6 z
<< end >>
