magic
tech scmos
timestamp 1199203435
<< ab >>
rect 0 0 144 80
<< nwell >>
rect -5 36 149 88
<< pwell >>
rect -5 -8 149 36
<< poly >>
rect 18 69 20 74
rect 28 69 30 74
rect 38 72 50 74
rect 38 69 40 72
rect 48 69 50 72
rect 69 70 71 74
rect 79 70 81 74
rect 91 70 93 74
rect 101 70 103 74
rect 118 70 120 74
rect 128 70 130 74
rect 2 39 8 41
rect 18 39 20 42
rect 28 39 30 42
rect 38 39 40 42
rect 2 37 4 39
rect 6 37 8 39
rect 16 37 31 39
rect 2 35 11 37
rect 9 30 11 35
rect 16 30 18 37
rect 25 35 27 37
rect 29 35 31 37
rect 25 33 31 35
rect 35 37 41 39
rect 48 38 50 42
rect 69 39 71 42
rect 79 39 81 42
rect 91 39 93 42
rect 101 39 103 42
rect 69 37 87 39
rect 35 35 37 37
rect 39 35 41 37
rect 81 35 83 37
rect 85 35 87 37
rect 35 33 41 35
rect 28 30 30 33
rect 35 30 37 33
rect 45 30 47 34
rect 55 30 57 35
rect 81 33 87 35
rect 91 37 104 39
rect 91 35 99 37
rect 101 35 104 37
rect 91 33 104 35
rect 108 37 114 39
rect 108 35 110 37
rect 112 35 114 37
rect 118 38 120 42
rect 128 39 130 42
rect 118 35 121 38
rect 108 33 114 35
rect 85 30 87 33
rect 92 30 94 33
rect 102 30 104 33
rect 109 30 111 33
rect 119 30 121 35
rect 128 37 135 39
rect 128 35 131 37
rect 133 35 135 37
rect 128 33 135 35
rect 129 30 131 33
rect 9 18 11 23
rect 16 18 18 23
rect 85 12 87 16
rect 92 12 94 16
rect 102 12 104 16
rect 109 12 111 16
rect 28 6 30 11
rect 35 6 37 11
rect 45 8 47 11
rect 55 8 57 11
rect 119 8 121 16
rect 129 8 131 16
rect 45 6 131 8
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 23 9 26
rect 11 23 16 30
rect 18 23 28 30
rect 20 13 28 23
rect 20 11 22 13
rect 24 11 28 13
rect 30 11 35 30
rect 37 21 45 30
rect 37 19 40 21
rect 42 19 45 21
rect 37 11 45 19
rect 47 28 55 30
rect 47 26 50 28
rect 52 26 55 28
rect 47 11 55 26
rect 57 23 62 30
rect 57 21 64 23
rect 57 19 60 21
rect 62 19 64 21
rect 57 17 64 19
rect 78 20 85 30
rect 78 18 80 20
rect 82 18 85 20
rect 57 11 62 17
rect 78 16 85 18
rect 87 16 92 30
rect 94 21 102 30
rect 94 19 97 21
rect 99 19 102 21
rect 94 16 102 19
rect 104 16 109 30
rect 111 20 119 30
rect 111 18 114 20
rect 116 18 119 20
rect 111 16 119 18
rect 121 28 129 30
rect 121 26 124 28
rect 126 26 129 28
rect 121 21 129 26
rect 121 19 124 21
rect 126 19 129 21
rect 121 16 129 19
rect 131 27 138 30
rect 131 25 134 27
rect 136 25 138 27
rect 131 20 138 25
rect 131 18 134 20
rect 136 18 138 20
rect 131 16 138 18
rect 20 9 26 11
<< pdif >>
rect 13 55 18 69
rect 11 53 18 55
rect 11 51 13 53
rect 15 51 18 53
rect 11 46 18 51
rect 11 44 13 46
rect 15 44 18 46
rect 11 42 18 44
rect 20 61 28 69
rect 20 59 23 61
rect 25 59 28 61
rect 20 42 28 59
rect 30 53 38 69
rect 30 51 33 53
rect 35 51 38 53
rect 30 42 38 51
rect 40 46 48 69
rect 40 44 43 46
rect 45 44 48 46
rect 40 42 48 44
rect 50 55 55 69
rect 62 68 69 70
rect 62 66 64 68
rect 66 66 69 68
rect 50 53 57 55
rect 50 51 53 53
rect 55 51 57 53
rect 50 46 57 51
rect 50 44 53 46
rect 55 44 57 46
rect 50 42 57 44
rect 62 42 69 66
rect 71 53 79 70
rect 71 51 74 53
rect 76 51 79 53
rect 71 46 79 51
rect 71 44 74 46
rect 76 44 79 46
rect 71 42 79 44
rect 81 68 91 70
rect 81 66 85 68
rect 87 66 91 68
rect 81 42 91 66
rect 93 53 101 70
rect 93 51 96 53
rect 98 51 101 53
rect 93 42 101 51
rect 103 68 118 70
rect 103 66 106 68
rect 108 66 113 68
rect 115 66 118 68
rect 103 61 118 66
rect 103 59 113 61
rect 115 59 118 61
rect 103 42 118 59
rect 120 46 128 70
rect 120 44 123 46
rect 125 44 128 46
rect 120 42 128 44
rect 130 68 138 70
rect 130 66 134 68
rect 136 66 138 68
rect 130 42 138 66
<< alu1 >>
rect -2 81 146 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 146 81
rect -2 68 146 79
rect 121 58 134 62
rect 10 53 57 54
rect 10 51 13 53
rect 15 51 33 53
rect 35 51 53 53
rect 55 51 57 53
rect 10 50 57 51
rect 10 46 16 50
rect 10 44 13 46
rect 15 44 16 46
rect 10 42 16 44
rect 52 46 57 50
rect 52 44 53 46
rect 55 44 57 46
rect 52 42 57 44
rect 10 31 14 42
rect 2 28 14 31
rect 2 26 4 28
rect 6 26 14 28
rect 81 42 119 46
rect 81 37 87 42
rect 81 35 83 37
rect 85 35 87 37
rect 81 34 87 35
rect 97 37 103 38
rect 97 35 99 37
rect 101 35 103 37
rect 97 30 103 35
rect 130 37 134 58
rect 130 35 131 37
rect 133 35 134 37
rect 130 33 134 35
rect 97 26 111 30
rect 2 25 14 26
rect 9 22 14 25
rect 9 21 64 22
rect 9 19 40 21
rect 42 19 60 21
rect 62 19 64 21
rect 9 18 64 19
rect -2 11 22 12
rect 24 11 146 12
rect -2 1 146 11
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 146 1
rect -2 -2 146 -1
<< ptie >>
rect 0 1 144 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 144 1
rect 0 -3 144 -1
<< ntie >>
rect 0 81 144 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 144 81
rect 0 77 144 79
<< nmos >>
rect 9 23 11 30
rect 16 23 18 30
rect 28 11 30 30
rect 35 11 37 30
rect 45 11 47 30
rect 55 11 57 30
rect 85 16 87 30
rect 92 16 94 30
rect 102 16 104 30
rect 109 16 111 30
rect 119 16 121 30
rect 129 16 131 30
<< pmos >>
rect 18 42 20 69
rect 28 42 30 69
rect 38 42 40 69
rect 48 42 50 69
rect 69 42 71 70
rect 79 42 81 70
rect 91 42 93 70
rect 101 42 103 70
rect 118 42 120 70
rect 128 42 130 70
<< polyct0 >>
rect 4 37 6 39
rect 27 35 29 37
rect 37 35 39 37
rect 110 35 112 37
<< polyct1 >>
rect 83 35 85 37
rect 99 35 101 37
rect 131 35 133 37
<< ndifct0 >>
rect 22 12 24 13
rect 50 26 52 28
rect 80 18 82 20
rect 97 19 99 21
rect 114 18 116 20
rect 124 26 126 28
rect 124 19 126 21
rect 134 25 136 27
rect 134 18 136 20
<< ndifct1 >>
rect 4 26 6 28
rect 22 11 24 12
rect 40 19 42 21
rect 60 19 62 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
<< pdifct0 >>
rect 23 59 25 61
rect 43 44 45 46
rect 64 66 66 68
rect 74 51 76 53
rect 74 44 76 46
rect 85 66 87 68
rect 96 51 98 53
rect 106 66 108 68
rect 113 66 115 68
rect 113 59 115 61
rect 123 44 125 46
rect 134 66 136 68
<< pdifct1 >>
rect 13 51 15 53
rect 13 44 15 46
rect 33 51 35 53
rect 53 51 55 53
rect 53 44 55 46
<< alu0 >>
rect 62 66 64 68
rect 66 66 68 68
rect 62 65 68 66
rect 83 66 85 68
rect 87 66 89 68
rect 83 65 89 66
rect 103 66 106 68
rect 108 66 113 68
rect 115 66 117 68
rect 103 65 117 66
rect 132 66 134 68
rect 136 66 138 68
rect 132 65 138 66
rect 2 61 107 62
rect 2 59 23 61
rect 25 59 107 61
rect 2 58 107 59
rect 111 61 117 65
rect 111 59 113 61
rect 115 59 117 61
rect 111 58 117 59
rect 2 41 6 58
rect 41 46 47 47
rect 26 44 43 46
rect 45 44 47 46
rect 26 42 47 44
rect 2 39 7 41
rect 2 37 4 39
rect 6 37 7 39
rect 2 35 7 37
rect 26 37 30 42
rect 61 38 65 58
rect 103 54 107 58
rect 26 35 27 37
rect 29 35 30 37
rect 26 30 30 35
rect 35 37 65 38
rect 35 35 37 37
rect 39 35 65 37
rect 35 34 65 35
rect 72 53 100 54
rect 72 51 74 53
rect 76 51 96 53
rect 98 51 100 53
rect 72 50 100 51
rect 103 50 126 54
rect 72 46 77 50
rect 122 46 126 50
rect 72 44 74 46
rect 76 44 77 46
rect 72 30 77 44
rect 122 44 123 46
rect 125 44 126 46
rect 108 37 114 42
rect 108 35 110 37
rect 112 35 114 37
rect 108 34 114 35
rect 122 30 126 44
rect 26 28 92 30
rect 26 26 50 28
rect 52 26 92 28
rect 122 28 127 30
rect 122 26 124 28
rect 126 26 127 28
rect 48 25 54 26
rect 88 22 92 26
rect 88 21 101 22
rect 78 20 84 21
rect 78 18 80 20
rect 82 18 84 20
rect 88 19 97 21
rect 99 19 101 21
rect 88 18 101 19
rect 113 20 117 22
rect 113 18 114 20
rect 116 18 117 20
rect 20 13 26 14
rect 20 12 22 13
rect 24 12 26 13
rect 69 12 73 16
rect 78 12 84 18
rect 113 12 117 18
rect 122 21 127 26
rect 122 19 124 21
rect 126 19 127 21
rect 122 17 127 19
rect 133 27 137 29
rect 133 25 134 27
rect 136 25 137 27
rect 133 20 137 25
rect 133 18 134 20
rect 136 18 137 20
rect 133 12 137 18
<< labels >>
rlabel alu0 4 48 4 48 6 bn
rlabel polyct0 28 36 28 36 6 an
rlabel alu0 44 44 44 44 6 an
rlabel alu0 50 36 50 36 6 bn
rlabel alu0 74 40 74 40 6 an
rlabel alu0 94 20 94 20 6 an
rlabel alu0 59 28 59 28 6 an
rlabel alu0 86 52 86 52 6 an
rlabel alu0 54 60 54 60 6 bn
rlabel alu0 124 35 124 35 6 bn
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 12 32 12 32 6 z
rlabel alu1 4 28 4 28 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 72 6 72 6 6 vss
rlabel alu1 100 32 100 32 6 a1
rlabel alu1 84 40 84 40 6 a2
rlabel alu1 100 44 100 44 6 a2
rlabel alu1 92 44 92 44 6 a2
rlabel alu1 72 74 72 74 6 vdd
rlabel alu1 108 28 108 28 6 a1
rlabel alu1 116 44 116 44 6 a2
rlabel alu1 132 44 132 44 6 b
rlabel alu1 108 44 108 44 6 a2
rlabel alu1 124 60 124 60 6 b
<< end >>
