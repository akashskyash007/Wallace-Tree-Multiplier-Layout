magic
tech scmos
timestamp 1199202715
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 30 39
rect 19 35 26 37
rect 28 35 30 37
rect 19 33 30 35
rect 12 30 14 33
rect 19 30 21 33
rect 12 7 14 12
rect 19 7 21 12
<< ndif >>
rect 7 22 12 30
rect 5 20 12 22
rect 5 18 7 20
rect 9 18 12 20
rect 5 16 12 18
rect 7 12 12 16
rect 14 12 19 30
rect 21 23 30 30
rect 21 21 26 23
rect 28 21 30 23
rect 21 16 30 21
rect 21 14 26 16
rect 28 14 30 16
rect 21 12 30 14
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 49 14 55
rect 2 21 6 49
rect 18 41 30 47
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 31 14 35
rect 26 37 30 41
rect 28 35 30 37
rect 26 33 30 35
rect 10 25 22 31
rect 2 20 11 21
rect 2 18 7 20
rect 9 18 11 20
rect 2 17 11 18
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 12 12 14 30
rect 19 12 21 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
<< polyct1 >>
rect 11 35 13 37
rect 26 35 28 37
<< ndifct0 >>
rect 26 21 28 23
rect 26 14 28 16
<< ndifct1 >>
rect 7 18 9 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 59 16 61
rect 14 52 16 54
rect 24 66 26 68
rect 24 59 26 61
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 55 17 59
rect 22 61 28 66
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 14 54 17 55
rect 16 52 17 54
rect 14 50 17 52
rect 24 34 26 41
rect 25 23 29 25
rect 25 21 26 23
rect 28 21 29 23
rect 25 16 29 21
rect 25 14 26 16
rect 28 14 29 16
rect 25 12 29 14
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 32 12 32 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 44 20 44 6 a
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 40 28 40 6 a
<< end >>
