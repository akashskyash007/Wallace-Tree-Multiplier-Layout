magic
tech scmos
timestamp 1199202484
<< ab >>
rect 0 0 144 80
<< nwell >>
rect -5 36 149 88
<< pwell >>
rect -5 -8 149 36
<< poly >>
rect 89 72 135 74
rect 19 66 21 71
rect 29 66 31 71
rect 89 69 91 72
rect 39 67 61 69
rect 9 60 11 65
rect 39 64 41 67
rect 49 64 51 67
rect 59 64 61 67
rect 69 67 91 69
rect 69 64 71 67
rect 79 64 81 67
rect 89 64 91 67
rect 99 64 101 68
rect 113 64 115 68
rect 123 64 125 68
rect 133 66 135 72
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 31 39
rect 39 38 41 42
rect 49 38 51 42
rect 59 39 61 42
rect 9 35 11 37
rect 13 35 19 37
rect 21 35 31 37
rect 9 33 31 35
rect 55 37 61 39
rect 69 38 71 42
rect 79 38 81 42
rect 89 38 91 42
rect 99 39 101 42
rect 113 39 115 42
rect 123 39 125 42
rect 133 39 135 42
rect 55 35 57 37
rect 59 35 61 37
rect 55 34 61 35
rect 99 37 125 39
rect 99 35 107 37
rect 109 35 115 37
rect 117 35 125 37
rect 9 30 11 33
rect 19 30 21 33
rect 29 30 31 33
rect 39 30 41 34
rect 49 30 51 34
rect 55 32 91 34
rect 9 15 11 19
rect 19 14 21 19
rect 29 14 31 19
rect 39 9 41 15
rect 69 29 71 32
rect 79 29 81 32
rect 89 29 91 32
rect 99 33 125 35
rect 129 37 135 39
rect 129 35 131 37
rect 133 35 135 37
rect 129 33 135 35
rect 99 29 101 33
rect 111 29 113 33
rect 121 29 123 33
rect 133 29 135 33
rect 69 13 71 18
rect 79 13 81 18
rect 89 13 91 18
rect 99 13 101 18
rect 111 13 113 18
rect 121 13 123 18
rect 49 9 51 12
rect 133 9 135 14
rect 39 7 135 9
<< ndif >>
rect 2 23 9 30
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 19 19 26
rect 21 23 29 30
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 19 39 26
rect 34 15 39 19
rect 41 28 49 30
rect 41 26 44 28
rect 46 26 49 28
rect 41 15 49 26
rect 44 12 49 15
rect 51 22 56 30
rect 62 27 69 29
rect 62 25 64 27
rect 66 25 69 27
rect 62 23 69 25
rect 51 20 58 22
rect 51 18 54 20
rect 56 18 58 20
rect 64 18 69 23
rect 71 22 79 29
rect 71 20 74 22
rect 76 20 79 22
rect 71 18 79 20
rect 81 27 89 29
rect 81 25 84 27
rect 86 25 89 27
rect 81 18 89 25
rect 91 27 99 29
rect 91 25 94 27
rect 96 25 99 27
rect 91 18 99 25
rect 101 18 111 29
rect 113 22 121 29
rect 113 20 116 22
rect 118 20 121 22
rect 113 18 121 20
rect 123 22 133 29
rect 123 20 127 22
rect 129 20 133 22
rect 123 18 133 20
rect 51 16 58 18
rect 51 12 56 16
rect 103 15 109 18
rect 103 13 105 15
rect 107 13 109 15
rect 125 14 133 18
rect 135 27 142 29
rect 135 25 138 27
rect 140 25 142 27
rect 135 23 142 25
rect 135 14 140 23
rect 103 11 109 13
<< pdif >>
rect 14 60 19 66
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 42 9 56
rect 11 53 19 60
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 56 29 62
rect 21 54 24 56
rect 26 54 29 56
rect 21 42 29 54
rect 31 64 36 66
rect 127 64 133 66
rect 31 61 39 64
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 53 49 64
rect 41 51 44 53
rect 46 51 49 53
rect 41 46 49 51
rect 41 44 44 46
rect 46 44 49 46
rect 41 42 49 44
rect 51 62 59 64
rect 51 60 54 62
rect 56 60 59 62
rect 51 42 59 60
rect 61 46 69 64
rect 61 44 64 46
rect 66 44 69 46
rect 61 42 69 44
rect 71 53 79 64
rect 71 51 74 53
rect 76 51 79 53
rect 71 46 79 51
rect 71 44 74 46
rect 76 44 79 46
rect 71 42 79 44
rect 81 46 89 64
rect 81 44 84 46
rect 86 44 89 46
rect 81 42 89 44
rect 91 53 99 64
rect 91 51 94 53
rect 96 51 99 53
rect 91 46 99 51
rect 91 44 94 46
rect 96 44 99 46
rect 91 42 99 44
rect 101 62 113 64
rect 101 60 108 62
rect 110 60 113 62
rect 101 42 113 60
rect 115 46 123 64
rect 115 44 118 46
rect 120 44 123 46
rect 115 42 123 44
rect 125 62 133 64
rect 125 60 128 62
rect 130 60 133 62
rect 125 42 133 60
rect 135 55 140 66
rect 135 53 142 55
rect 135 51 138 53
rect 140 51 142 53
rect 135 46 142 51
rect 135 44 138 46
rect 140 44 142 46
rect 135 42 142 44
<< alu1 >>
rect -2 81 146 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 146 81
rect -2 68 146 79
rect 2 38 6 47
rect 2 37 23 38
rect 2 35 11 37
rect 13 35 19 37
rect 21 35 23 37
rect 2 34 23 35
rect 2 33 6 34
rect 42 53 47 55
rect 42 51 44 53
rect 46 51 47 53
rect 42 46 47 51
rect 42 44 44 46
rect 46 44 47 46
rect 42 30 47 44
rect 63 46 67 48
rect 63 44 64 46
rect 66 44 67 46
rect 63 30 67 44
rect 82 46 87 48
rect 82 44 84 46
rect 86 44 87 46
rect 82 30 87 44
rect 42 28 88 30
rect 42 26 44 28
rect 46 27 88 28
rect 46 26 64 27
rect 42 24 47 26
rect 63 25 64 26
rect 66 26 84 27
rect 66 25 67 26
rect 63 23 67 25
rect 82 25 84 26
rect 86 25 88 27
rect 82 24 88 25
rect 105 37 119 38
rect 105 35 107 37
rect 109 35 115 37
rect 117 35 119 37
rect 105 34 119 35
rect 130 37 134 47
rect 130 35 131 37
rect 133 35 134 37
rect 105 26 111 34
rect 130 30 134 35
rect 121 26 134 30
rect -2 1 146 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 146 1
rect -2 -2 146 -1
<< ptie >>
rect 0 1 144 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 144 1
rect 0 -3 144 -1
<< ntie >>
rect 0 81 144 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 144 81
rect 0 77 144 79
<< nmos >>
rect 9 19 11 30
rect 19 19 21 30
rect 29 19 31 30
rect 39 15 41 30
rect 49 12 51 30
rect 69 18 71 29
rect 79 18 81 29
rect 89 18 91 29
rect 99 18 101 29
rect 111 18 113 29
rect 121 18 123 29
rect 133 14 135 29
<< pmos >>
rect 9 42 11 60
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 64
rect 49 42 51 64
rect 59 42 61 64
rect 69 42 71 64
rect 79 42 81 64
rect 89 42 91 64
rect 99 42 101 64
rect 113 42 115 64
rect 123 42 125 64
rect 133 42 135 66
<< polyct0 >>
rect 57 35 59 37
<< polyct1 >>
rect 11 35 13 37
rect 19 35 21 37
rect 107 35 109 37
rect 115 35 117 37
rect 131 35 133 37
<< ndifct0 >>
rect 4 21 6 23
rect 14 26 16 28
rect 24 21 26 23
rect 34 26 36 28
rect 54 18 56 20
rect 74 20 76 22
rect 94 25 96 27
rect 116 20 118 22
rect 127 20 129 22
rect 105 13 107 15
rect 138 25 140 27
<< ndifct1 >>
rect 44 26 46 28
rect 64 25 66 27
rect 84 25 86 27
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
<< pdifct0 >>
rect 4 56 6 58
rect 14 51 16 53
rect 14 44 16 46
rect 24 62 26 64
rect 24 54 26 56
rect 34 59 36 61
rect 34 51 36 53
rect 34 44 36 46
rect 54 60 56 62
rect 74 51 76 53
rect 74 44 76 46
rect 94 51 96 53
rect 94 44 96 46
rect 108 60 110 62
rect 118 44 120 46
rect 128 60 130 62
rect 138 51 140 53
rect 138 44 140 46
<< pdifct1 >>
rect 44 51 46 53
rect 44 44 46 46
rect 64 44 66 46
rect 84 44 86 46
<< alu0 >>
rect 3 58 7 68
rect 3 56 4 58
rect 6 56 7 58
rect 3 54 7 56
rect 23 64 27 68
rect 23 62 24 64
rect 26 62 27 64
rect 23 56 27 62
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 23 54 24 56
rect 26 54 27 56
rect 23 52 27 54
rect 33 62 58 63
rect 33 61 54 62
rect 33 59 34 61
rect 36 60 54 61
rect 56 60 58 62
rect 36 59 58 60
rect 63 59 104 63
rect 33 53 37 59
rect 63 55 67 59
rect 100 55 104 59
rect 107 62 111 68
rect 107 60 108 62
rect 110 60 111 62
rect 107 58 111 60
rect 126 62 132 68
rect 126 60 128 62
rect 130 60 132 62
rect 126 59 132 60
rect 13 46 17 51
rect 33 51 34 53
rect 36 51 37 53
rect 33 46 37 51
rect 13 44 14 46
rect 16 44 34 46
rect 36 44 37 46
rect 13 42 37 44
rect 33 31 37 42
rect 13 28 37 31
rect 13 26 14 28
rect 16 27 34 28
rect 16 26 17 27
rect 3 23 7 25
rect 13 24 17 26
rect 33 26 34 27
rect 36 26 37 28
rect 3 21 4 23
rect 6 21 7 23
rect 3 12 7 21
rect 22 23 28 24
rect 22 21 24 23
rect 26 21 28 23
rect 22 12 28 21
rect 33 21 37 26
rect 56 51 67 55
rect 73 53 97 55
rect 73 51 74 53
rect 76 51 94 53
rect 96 51 97 53
rect 100 53 142 55
rect 100 51 138 53
rect 140 51 142 53
rect 56 37 60 51
rect 56 35 57 37
rect 59 35 60 37
rect 56 33 60 35
rect 73 46 77 51
rect 73 44 74 46
rect 76 44 77 46
rect 73 42 77 44
rect 92 47 97 51
rect 92 46 122 47
rect 92 44 94 46
rect 96 44 118 46
rect 120 44 122 46
rect 92 43 122 44
rect 93 27 97 43
rect 93 25 94 27
rect 96 25 97 27
rect 137 46 142 51
rect 137 44 138 46
rect 140 44 142 46
rect 137 42 142 44
rect 138 29 142 42
rect 137 27 142 29
rect 93 23 97 25
rect 137 25 138 27
rect 140 25 142 27
rect 137 23 142 25
rect 72 22 78 23
rect 33 20 58 21
rect 33 18 54 20
rect 56 18 58 20
rect 33 17 58 18
rect 72 20 74 22
rect 76 21 78 22
rect 93 22 120 23
rect 93 21 116 22
rect 76 20 116 21
rect 118 20 120 22
rect 72 19 120 20
rect 125 22 131 23
rect 125 20 127 22
rect 129 20 131 22
rect 72 17 97 19
rect 103 15 109 16
rect 103 13 105 15
rect 107 13 109 15
rect 103 12 109 13
rect 125 12 131 20
<< labels >>
rlabel alu0 15 48 15 48 6 a1n
rlabel alu0 25 29 25 29 6 a1n
rlabel alu0 35 40 35 40 6 a1n
rlabel alu0 45 19 45 19 6 a1n
rlabel alu0 75 48 75 48 6 a0n
rlabel alu0 58 44 58 44 6 sn
rlabel alu0 45 61 45 61 6 a1n
rlabel alu0 84 19 84 19 6 a0n
rlabel alu0 95 36 95 36 6 a0n
rlabel alu0 106 21 106 21 6 a0n
rlabel alu0 107 45 107 45 6 a0n
rlabel alu0 140 39 140 39 6 sn
rlabel polyct1 12 36 12 36 6 a1
rlabel polyct1 20 36 20 36 6 a1
rlabel alu1 4 40 4 40 6 a1
rlabel alu1 52 28 52 28 6 z
rlabel alu1 60 28 60 28 6 z
rlabel alu1 68 28 68 28 6 z
rlabel alu1 44 40 44 40 6 z
rlabel alu1 72 6 72 6 6 vss
rlabel alu1 76 28 76 28 6 z
rlabel alu1 84 36 84 36 6 z
rlabel alu1 72 74 72 74 6 vdd
rlabel alu1 108 32 108 32 6 a0
rlabel alu1 124 28 124 28 6 s
rlabel polyct1 116 36 116 36 6 a0
rlabel alu1 132 40 132 40 6 s
<< end >>
