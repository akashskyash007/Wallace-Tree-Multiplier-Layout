magic
tech scmos
timestamp 1199202444
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 62 11 67
rect 16 62 18 67
rect 26 62 28 67
rect 33 62 35 67
rect 45 58 51 60
rect 45 56 47 58
rect 49 56 51 58
rect 45 54 51 56
rect 45 51 47 54
rect 9 43 11 46
rect 2 41 11 43
rect 2 39 4 41
rect 6 39 8 41
rect 2 37 8 39
rect 16 37 18 46
rect 26 43 28 46
rect 23 41 29 43
rect 23 39 25 41
rect 27 39 29 41
rect 23 37 29 39
rect 6 23 8 37
rect 12 35 18 37
rect 12 33 14 35
rect 16 33 18 35
rect 33 36 35 46
rect 45 42 47 45
rect 45 40 52 42
rect 33 34 46 36
rect 12 31 28 33
rect 16 25 22 27
rect 16 23 18 25
rect 20 23 22 25
rect 6 21 11 23
rect 9 18 11 21
rect 16 21 22 23
rect 16 18 18 21
rect 26 18 28 31
rect 33 32 42 34
rect 44 32 46 34
rect 33 30 46 32
rect 33 18 35 30
rect 50 26 52 40
rect 45 24 52 26
rect 45 21 47 24
rect 45 11 47 15
rect 9 6 11 11
rect 16 6 18 11
rect 26 6 28 11
rect 33 6 35 11
<< ndif >>
rect 37 18 45 21
rect 2 15 9 18
rect 2 13 4 15
rect 6 13 9 15
rect 2 11 9 13
rect 11 11 16 18
rect 18 16 26 18
rect 18 14 21 16
rect 23 14 26 16
rect 18 11 26 14
rect 28 11 33 18
rect 35 15 45 18
rect 47 19 54 21
rect 47 17 50 19
rect 52 17 54 19
rect 47 15 54 17
rect 35 11 43 15
rect 37 7 43 11
rect 37 5 39 7
rect 41 5 43 7
rect 37 3 43 5
<< pdif >>
rect 37 67 43 69
rect 37 65 39 67
rect 41 65 43 67
rect 37 62 43 65
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 46 9 58
rect 11 46 16 62
rect 18 50 26 62
rect 18 48 21 50
rect 23 48 26 50
rect 18 46 26 48
rect 28 46 33 62
rect 35 51 43 62
rect 35 46 45 51
rect 37 45 45 46
rect 47 49 54 51
rect 47 47 50 49
rect 52 47 54 49
rect 47 45 54 47
<< alu1 >>
rect -2 67 58 72
rect -2 65 39 67
rect 41 65 49 67
rect 51 65 58 67
rect -2 64 58 65
rect 45 58 51 59
rect 11 56 47 58
rect 49 56 51 58
rect 11 54 51 56
rect 11 51 15 54
rect 2 46 15 51
rect 19 48 21 50
rect 23 48 38 50
rect 19 46 38 48
rect 2 41 8 46
rect 2 39 4 41
rect 6 39 8 41
rect 2 38 8 39
rect 23 41 30 42
rect 23 39 25 41
rect 27 39 30 41
rect 23 38 30 39
rect 12 35 18 36
rect 12 34 14 35
rect 2 33 14 34
rect 16 33 18 35
rect 2 30 18 33
rect 2 21 6 30
rect 26 26 30 38
rect 16 25 30 26
rect 16 23 18 25
rect 20 23 30 25
rect 16 22 30 23
rect 34 18 38 46
rect 17 16 38 18
rect 17 14 21 16
rect 23 14 38 16
rect 17 13 38 14
rect -2 7 58 8
rect -2 5 39 7
rect 41 5 49 7
rect 51 5 58 7
rect -2 0 58 5
<< ptie >>
rect 47 7 53 9
rect 47 5 49 7
rect 51 5 53 7
rect 47 3 53 5
<< ntie >>
rect 47 67 53 69
rect 47 65 49 67
rect 51 65 53 67
rect 47 63 53 65
<< nmos >>
rect 9 11 11 18
rect 16 11 18 18
rect 26 11 28 18
rect 33 11 35 18
rect 45 15 47 21
<< pmos >>
rect 9 46 11 62
rect 16 46 18 62
rect 26 46 28 62
rect 33 46 35 62
rect 45 45 47 51
<< polyct0 >>
rect 42 32 44 34
<< polyct1 >>
rect 47 56 49 58
rect 4 39 6 41
rect 25 39 27 41
rect 14 33 16 35
rect 18 23 20 25
<< ndifct0 >>
rect 4 13 6 15
rect 50 17 52 19
<< ndifct1 >>
rect 21 14 23 16
rect 39 5 41 7
<< ntiect1 >>
rect 49 65 51 67
<< ptiect1 >>
rect 49 5 51 7
<< pdifct0 >>
rect 4 58 6 60
rect 50 47 52 49
<< pdifct1 >>
rect 39 65 41 67
rect 21 48 23 50
<< alu0 >>
rect 3 60 7 64
rect 3 58 4 60
rect 6 58 7 60
rect 3 56 7 58
rect 19 50 25 51
rect 49 49 53 51
rect 49 47 50 49
rect 52 47 53 49
rect 49 36 53 47
rect 41 34 53 36
rect 41 32 42 34
rect 44 32 53 34
rect 41 30 53 32
rect 3 15 7 17
rect 3 13 4 15
rect 6 13 7 15
rect 49 19 53 30
rect 49 17 50 19
rect 52 17 53 19
rect 49 15 53 17
rect 3 8 7 13
<< labels >>
rlabel alu0 47 33 47 33 6 sn
rlabel alu0 51 33 51 33 6 sn
rlabel alu1 4 24 4 24 6 a0
rlabel alu1 4 48 4 48 6 s
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 32 12 32 6 a0
rlabel alu1 20 24 20 24 6 a1
rlabel alu1 12 48 12 48 6 s
rlabel alu1 20 56 20 56 6 s
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 16 28 16 6 z
rlabel alu1 28 32 28 32 6 a1
rlabel alu1 36 28 36 28 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 56 36 56 6 s
rlabel alu1 28 56 28 56 6 s
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 56 44 56 6 s
<< end >>
