magic
tech scmos
timestamp 1199475729
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< alu1 >>
rect -2 97 72 102
rect -2 95 47 97
rect 49 95 55 97
rect 57 95 72 97
rect -2 88 72 95
rect -2 9 72 12
rect -2 7 15 9
rect 17 7 23 9
rect 25 7 72 9
rect -2 -2 72 7
<< alu2 >>
rect 7 97 63 102
rect 7 95 15 97
rect 17 95 23 97
rect 25 95 47 97
rect 49 95 55 97
rect 57 95 63 97
rect 7 88 63 95
rect 7 9 63 12
rect 7 7 15 9
rect 17 7 23 9
rect 25 7 47 9
rect 49 7 55 9
rect 57 7 63 9
rect 7 -2 63 7
<< alu3 >>
rect 8 97 32 102
rect 8 95 15 97
rect 17 95 23 97
rect 25 95 32 97
rect 8 -2 32 95
rect 38 9 62 102
rect 38 7 47 9
rect 49 7 55 9
rect 57 7 62 9
rect 38 -2 62 7
<< via1 >>
rect 47 95 49 97
rect 55 95 57 97
rect 15 7 17 9
rect 23 7 25 9
<< via2 >>
rect 15 95 17 97
rect 23 95 25 97
rect 47 7 49 9
rect 55 7 57 9
<< labels >>
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 35 94 35 94 6 vdd
rlabel alu2 35 6 35 6 6 vss
rlabel alu2 35 94 35 94 6 vdd
rlabel alu3 20 50 20 50 6 vdd
rlabel alu3 50 50 50 50 6 vss
<< end >>
