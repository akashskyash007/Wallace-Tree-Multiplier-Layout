magic
tech scmos
timestamp 1199201954
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 31 60 33 65
rect 41 60 43 65
rect 53 60 55 65
rect 9 50 11 55
rect 9 35 11 38
rect 31 35 33 44
rect 41 35 43 44
rect 53 41 55 44
rect 53 39 62 41
rect 53 37 58 39
rect 60 37 62 39
rect 53 35 62 37
rect 9 33 19 35
rect 13 31 15 33
rect 17 31 19 33
rect 13 29 19 31
rect 31 33 37 35
rect 31 31 33 33
rect 35 31 37 33
rect 31 29 37 31
rect 41 33 47 35
rect 41 31 43 33
rect 45 31 47 33
rect 41 29 47 31
rect 13 26 15 29
rect 13 15 15 20
rect 31 19 33 29
rect 41 19 43 29
rect 53 24 55 35
rect 48 22 55 24
rect 48 19 50 22
rect 31 8 33 13
rect 41 7 43 12
rect 48 7 50 12
<< ndif >>
rect 6 24 13 26
rect 6 22 8 24
rect 10 22 13 24
rect 6 20 13 22
rect 15 24 23 26
rect 15 22 19 24
rect 21 22 23 24
rect 15 20 23 22
rect 17 19 23 20
rect 17 17 31 19
rect 17 15 19 17
rect 21 15 26 17
rect 28 15 31 17
rect 17 13 31 15
rect 33 17 41 19
rect 33 15 36 17
rect 38 15 41 17
rect 33 13 41 15
rect 36 12 41 13
rect 43 12 48 19
rect 50 16 57 19
rect 50 14 53 16
rect 55 14 57 16
rect 50 12 57 14
<< pdif >>
rect 45 67 51 69
rect 45 65 47 67
rect 49 65 51 67
rect 45 60 51 65
rect 26 57 31 60
rect 24 55 31 57
rect 24 53 26 55
rect 28 53 31 55
rect 4 44 9 50
rect 2 42 9 44
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 48 18 50
rect 11 46 14 48
rect 16 46 18 48
rect 11 38 18 46
rect 24 48 31 53
rect 24 46 26 48
rect 28 46 31 48
rect 24 44 31 46
rect 33 58 41 60
rect 33 56 36 58
rect 38 56 41 58
rect 33 44 41 56
rect 43 44 53 60
rect 55 58 62 60
rect 55 56 58 58
rect 60 56 62 58
rect 55 54 62 56
rect 55 44 60 54
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 13 67
rect 15 65 47 67
rect 49 65 66 67
rect -2 64 66 65
rect 2 42 7 44
rect 2 40 4 42
rect 6 40 7 42
rect 2 38 7 40
rect 2 27 6 38
rect 34 45 46 51
rect 50 45 62 51
rect 34 35 38 45
rect 57 39 62 45
rect 57 37 58 39
rect 60 37 62 39
rect 57 35 62 37
rect 2 24 14 27
rect 32 33 38 35
rect 32 31 33 33
rect 35 31 38 33
rect 32 29 38 31
rect 42 33 46 35
rect 42 31 43 33
rect 45 31 46 33
rect 42 26 46 31
rect 2 22 8 24
rect 10 22 14 24
rect 2 21 14 22
rect 42 22 55 26
rect 2 13 6 21
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 13 7
rect 15 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 17 9
rect 3 5 5 7
rect 7 5 13 7
rect 15 5 17 7
rect 3 3 17 5
<< ntie >>
rect 3 67 17 69
rect 3 65 5 67
rect 7 65 13 67
rect 15 65 17 67
rect 3 63 17 65
<< nmos >>
rect 13 20 15 26
rect 31 13 33 19
rect 41 12 43 19
rect 48 12 50 19
<< pmos >>
rect 9 38 11 50
rect 31 44 33 60
rect 41 44 43 60
rect 53 44 55 60
<< polyct0 >>
rect 15 31 17 33
<< polyct1 >>
rect 58 37 60 39
rect 33 31 35 33
rect 43 31 45 33
<< ndifct0 >>
rect 19 22 21 24
rect 19 15 21 17
rect 26 15 28 17
rect 36 15 38 17
rect 53 14 55 16
<< ndifct1 >>
rect 8 22 10 24
<< ntiect1 >>
rect 5 65 7 67
rect 13 65 15 67
<< ptiect1 >>
rect 5 5 7 7
rect 13 5 15 7
<< pdifct0 >>
rect 26 53 28 55
rect 14 46 16 48
rect 26 46 28 48
rect 36 56 38 58
rect 58 56 60 58
<< pdifct1 >>
rect 47 65 49 67
rect 4 40 6 42
<< alu0 >>
rect 13 48 17 64
rect 34 58 62 59
rect 13 46 14 48
rect 16 46 17 48
rect 13 44 17 46
rect 25 55 29 57
rect 34 56 36 58
rect 38 56 58 58
rect 60 56 62 58
rect 34 55 62 56
rect 25 53 26 55
rect 28 53 29 55
rect 25 48 29 53
rect 25 46 26 48
rect 28 46 29 48
rect 25 34 29 46
rect 13 33 29 34
rect 13 31 15 33
rect 17 31 29 33
rect 13 30 29 31
rect 25 26 29 30
rect 18 24 22 26
rect 18 22 19 24
rect 21 22 22 24
rect 25 22 39 26
rect 18 18 22 22
rect 18 17 30 18
rect 18 15 19 17
rect 21 15 26 17
rect 28 15 30 17
rect 18 14 30 15
rect 35 17 39 22
rect 35 15 36 17
rect 38 15 39 17
rect 18 8 22 14
rect 35 13 39 15
rect 52 16 56 18
rect 52 14 53 16
rect 55 14 56 16
rect 52 8 56 14
<< labels >>
rlabel alu0 48 57 48 57 6 n1
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel polyct1 44 32 44 32 6 a2
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 48 44 48 6 b
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 24 52 24 6 a2
rlabel alu1 52 48 52 48 6 a1
rlabel alu1 60 44 60 44 6 a1
<< end >>
