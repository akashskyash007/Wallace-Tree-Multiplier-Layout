magic
tech scmos
timestamp 1199201822
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 63 11 68
rect 21 63 23 68
rect 41 63 43 68
rect 51 63 53 68
rect 61 63 63 68
rect 9 48 11 51
rect 9 46 15 48
rect 9 44 11 46
rect 13 44 15 46
rect 9 42 15 44
rect 9 22 11 42
rect 21 38 23 51
rect 41 39 43 47
rect 51 39 53 47
rect 61 44 63 47
rect 60 42 70 44
rect 60 40 66 42
rect 68 40 70 42
rect 16 36 24 38
rect 16 34 18 36
rect 20 34 24 36
rect 16 32 24 34
rect 33 37 43 39
rect 33 35 35 37
rect 37 35 43 37
rect 49 37 55 39
rect 49 35 51 37
rect 53 35 55 37
rect 33 33 45 35
rect 49 33 55 35
rect 22 29 24 32
rect 43 30 45 33
rect 53 30 55 33
rect 60 38 70 40
rect 60 30 62 38
rect 22 18 24 23
rect 9 11 11 16
rect 43 19 45 24
rect 53 18 55 23
rect 60 18 62 23
<< ndif >>
rect 13 23 22 29
rect 24 27 31 29
rect 24 25 27 27
rect 29 25 31 27
rect 24 23 31 25
rect 35 24 43 30
rect 45 28 53 30
rect 45 26 48 28
rect 50 26 53 28
rect 45 24 53 26
rect 13 22 20 23
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 20 22
rect 13 11 20 16
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
rect 35 11 41 24
rect 48 23 53 24
rect 55 23 60 30
rect 62 27 69 30
rect 62 25 65 27
rect 67 25 69 27
rect 62 23 69 25
rect 35 9 37 11
rect 39 9 41 11
rect 35 7 41 9
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 63 19 69
rect 4 57 9 63
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 51 9 53
rect 11 51 21 63
rect 23 57 28 63
rect 23 55 30 57
rect 23 53 26 55
rect 28 53 30 55
rect 36 53 41 63
rect 23 51 30 53
rect 34 51 41 53
rect 34 49 36 51
rect 38 49 41 51
rect 34 47 41 49
rect 43 61 51 63
rect 43 59 46 61
rect 48 59 51 61
rect 43 54 51 59
rect 43 52 46 54
rect 48 52 51 54
rect 43 47 51 52
rect 53 61 61 63
rect 53 59 56 61
rect 58 59 61 61
rect 53 47 61 59
rect 63 61 70 63
rect 63 59 66 61
rect 68 59 70 61
rect 63 54 70 59
rect 63 52 66 54
rect 68 52 70 54
rect 63 50 70 52
rect 63 47 68 50
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 71 74 79
rect -2 69 15 71
rect 17 69 74 71
rect -2 68 74 69
rect 10 57 22 63
rect 10 46 14 57
rect 10 44 11 46
rect 13 44 14 46
rect 10 41 14 44
rect 18 37 22 47
rect 10 36 22 37
rect 10 34 18 36
rect 20 34 22 36
rect 10 33 22 34
rect 34 51 39 56
rect 34 49 36 51
rect 38 49 39 51
rect 34 47 39 49
rect 34 43 46 47
rect 10 25 14 33
rect 42 29 46 43
rect 57 42 70 47
rect 65 40 66 42
rect 68 40 70 42
rect 42 28 52 29
rect 42 26 48 28
rect 50 26 52 28
rect 42 25 52 26
rect 65 33 70 40
rect -2 11 74 12
rect -2 9 15 11
rect 17 9 37 11
rect 39 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 22 23 24 29
rect 43 24 45 30
rect 9 16 11 22
rect 53 23 55 30
rect 60 23 62 30
<< pmos >>
rect 9 51 11 63
rect 21 51 23 63
rect 41 47 43 63
rect 51 47 53 63
rect 61 47 63 63
<< polyct0 >>
rect 35 35 37 37
rect 51 35 53 37
<< polyct1 >>
rect 11 44 13 46
rect 66 40 68 42
rect 18 34 20 36
<< ndifct0 >>
rect 27 25 29 27
rect 4 18 6 20
rect 65 25 67 27
<< ndifct1 >>
rect 48 26 50 28
rect 15 9 17 11
rect 37 9 39 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 53 6 55
rect 26 53 28 55
rect 46 59 48 61
rect 46 52 48 54
rect 56 59 58 61
rect 66 59 68 61
rect 66 52 68 54
<< pdifct1 >>
rect 15 69 17 71
rect 36 49 38 51
<< alu0 >>
rect 44 61 50 62
rect 44 59 46 61
rect 48 59 50 61
rect 2 55 7 57
rect 2 53 4 55
rect 6 53 7 55
rect 2 51 7 53
rect 2 21 6 51
rect 25 55 29 57
rect 25 53 26 55
rect 28 53 29 55
rect 25 38 29 53
rect 44 55 50 59
rect 54 61 60 68
rect 54 59 56 61
rect 58 59 60 61
rect 54 58 60 59
rect 64 61 70 62
rect 64 59 66 61
rect 68 59 70 61
rect 64 55 70 59
rect 44 54 70 55
rect 44 52 46 54
rect 48 52 66 54
rect 68 52 70 54
rect 44 51 70 52
rect 25 37 39 38
rect 25 35 35 37
rect 37 35 39 37
rect 25 34 39 35
rect 25 27 31 34
rect 25 25 27 27
rect 29 25 31 27
rect 49 37 60 38
rect 49 35 51 37
rect 53 35 60 37
rect 49 34 60 35
rect 25 24 31 25
rect 56 21 60 34
rect 2 20 60 21
rect 2 18 4 20
rect 6 18 60 20
rect 2 17 60 18
rect 64 27 68 29
rect 64 25 65 27
rect 67 25 68 27
rect 64 12 68 25
<< labels >>
rlabel alu0 4 54 4 54 6 a2n
rlabel alu0 27 40 27 40 6 bn
rlabel alu0 32 36 32 36 6 bn
rlabel alu0 47 56 47 56 6 n1
rlabel alu0 31 19 31 19 6 a2n
rlabel alu0 54 36 54 36 6 a2n
rlabel alu0 57 53 57 53 6 n1
rlabel alu0 67 56 67 56 6 n1
rlabel alu1 12 28 12 28 6 b
rlabel alu1 12 52 12 52 6 a2
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 60 20 60 6 a2
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 44 36 44 36 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 44 60 44 6 a1
rlabel alu1 68 40 68 40 6 a1
<< end >>
