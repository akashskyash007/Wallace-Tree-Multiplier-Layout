magic
tech scmos
timestamp 1199470706
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 11 83 13 88
rect 23 83 25 88
rect 35 83 37 88
rect 57 82 64 84
rect 57 80 60 82
rect 62 80 64 82
rect 57 78 64 80
rect 57 75 59 78
rect 11 47 13 63
rect 23 54 25 63
rect 35 60 37 63
rect 35 58 47 60
rect 23 52 41 54
rect 23 51 27 52
rect 11 45 21 47
rect 11 44 17 45
rect 13 43 17 44
rect 19 43 21 45
rect 13 41 21 43
rect 13 26 15 41
rect 25 31 27 51
rect 35 50 37 52
rect 39 50 41 52
rect 35 48 41 50
rect 45 43 47 58
rect 45 41 51 43
rect 45 39 47 41
rect 49 39 51 41
rect 45 37 51 39
rect 21 29 27 31
rect 21 26 23 29
rect 33 26 35 31
rect 45 26 47 37
rect 57 26 59 55
rect 13 12 15 17
rect 21 12 23 17
rect 33 5 35 17
rect 45 12 47 17
rect 57 5 59 17
rect 33 3 59 5
<< ndif >>
rect 4 21 13 26
rect 4 19 7 21
rect 9 19 13 21
rect 4 17 13 19
rect 15 17 21 26
rect 23 21 33 26
rect 23 19 27 21
rect 29 19 33 21
rect 23 17 33 19
rect 35 21 45 26
rect 35 19 39 21
rect 41 19 45 21
rect 35 17 45 19
rect 47 17 57 26
rect 59 23 64 26
rect 59 21 67 23
rect 59 19 63 21
rect 65 19 67 21
rect 59 17 67 19
rect 49 11 55 17
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
<< pdif >>
rect 39 91 55 93
rect 39 89 41 91
rect 43 89 51 91
rect 53 89 55 91
rect 39 83 55 89
rect 3 81 11 83
rect 3 79 5 81
rect 7 79 11 81
rect 3 77 11 79
rect 6 63 11 77
rect 13 71 23 83
rect 13 69 17 71
rect 19 69 23 71
rect 13 63 23 69
rect 25 71 35 83
rect 25 69 29 71
rect 31 69 35 71
rect 25 63 35 69
rect 37 81 55 83
rect 37 79 51 81
rect 53 79 55 81
rect 37 75 55 79
rect 37 63 57 75
rect 50 55 57 63
rect 59 61 64 75
rect 59 59 67 61
rect 59 57 63 59
rect 65 57 67 59
rect 59 55 67 57
<< alu1 >>
rect -2 95 72 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 72 95
rect -2 91 72 93
rect -2 89 41 91
rect 43 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 3 81 40 82
rect 3 79 5 81
rect 7 79 40 81
rect 3 78 40 79
rect 8 71 23 73
rect 8 69 17 71
rect 19 69 23 71
rect 8 68 23 69
rect 28 71 32 73
rect 28 69 29 71
rect 31 69 32 71
rect 8 33 12 68
rect 28 47 32 69
rect 36 52 40 78
rect 50 81 54 88
rect 50 79 51 81
rect 53 79 54 81
rect 50 77 54 79
rect 58 82 64 83
rect 58 80 60 82
rect 62 80 64 82
rect 58 73 64 80
rect 48 67 64 73
rect 48 57 52 67
rect 62 59 66 61
rect 62 57 63 59
rect 65 57 66 59
rect 62 52 66 57
rect 36 50 37 52
rect 39 50 66 52
rect 36 48 66 50
rect 16 45 32 47
rect 16 43 17 45
rect 19 43 32 45
rect 16 41 32 43
rect 8 27 22 33
rect 28 32 32 41
rect 37 41 52 43
rect 37 39 47 41
rect 49 39 52 41
rect 37 38 52 39
rect 28 28 42 32
rect 6 21 10 23
rect 6 19 7 21
rect 9 19 10 21
rect 6 12 10 19
rect 18 22 22 27
rect 18 21 33 22
rect 18 19 27 21
rect 29 19 33 21
rect 18 17 33 19
rect 38 21 42 28
rect 38 19 39 21
rect 41 19 42 21
rect 38 17 42 19
rect 48 17 52 38
rect 62 21 66 48
rect 62 19 63 21
rect 65 19 66 21
rect 62 17 66 19
rect -2 11 72 12
rect -2 9 51 11
rect 53 9 72 11
rect -2 7 72 9
rect -2 5 10 7
rect 12 5 19 7
rect 21 5 72 7
rect -2 0 72 5
<< ptie >>
rect 8 7 23 9
rect 8 5 10 7
rect 12 5 19 7
rect 21 5 23 7
rect 8 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 13 17 15 26
rect 21 17 23 26
rect 33 17 35 26
rect 45 17 47 26
rect 57 17 59 26
<< pmos >>
rect 11 63 13 83
rect 23 63 25 83
rect 35 63 37 83
rect 57 55 59 75
<< polyct1 >>
rect 60 80 62 82
rect 17 43 19 45
rect 37 50 39 52
rect 47 39 49 41
<< ndifct1 >>
rect 7 19 9 21
rect 27 19 29 21
rect 39 19 41 21
rect 63 19 65 21
rect 51 9 53 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 10 5 12 7
rect 19 5 21 7
<< pdifct1 >>
rect 41 89 43 91
rect 51 89 53 91
rect 5 79 7 81
rect 17 69 19 71
rect 29 69 31 71
rect 51 79 53 81
rect 63 57 65 59
<< labels >>
rlabel polyct1 18 44 18 44 6 an
rlabel pdifct1 6 80 6 80 6 bn
rlabel ndifct1 40 20 40 20 6 an
rlabel polyct1 38 51 38 51 6 bn
rlabel pdifct1 30 70 30 70 6 an
rlabel ndifct1 64 20 64 20 6 bn
rlabel pdifct1 64 58 64 58 6 bn
rlabel alu1 10 50 10 50 6 z
rlabel alu1 30 20 30 20 6 z
rlabel alu1 20 25 20 25 6 z
rlabel alu1 20 70 20 70 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 50 30 50 30 6 a
rlabel alu1 40 40 40 40 6 a
rlabel alu1 50 65 50 65 6 b
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 75 60 75 6 b
<< end >>
