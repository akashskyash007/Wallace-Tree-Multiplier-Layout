magic
tech scmos
timestamp 1199203533
<< ab >>
rect 0 0 96 72
<< nwell >>
rect -5 32 101 77
<< pwell >>
rect -5 -5 101 32
<< poly >>
rect 12 66 14 70
rect 19 66 21 70
rect 31 66 33 70
rect 38 66 40 70
rect 48 66 50 70
rect 58 66 60 70
rect 68 66 70 70
rect 75 66 77 70
rect 85 66 87 70
rect 12 35 14 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 9 26 11 29
rect 19 26 21 38
rect 31 35 33 46
rect 38 43 40 46
rect 48 43 50 46
rect 58 43 60 46
rect 68 43 70 46
rect 38 41 43 43
rect 48 41 61 43
rect 41 37 43 41
rect 55 39 57 41
rect 59 39 61 41
rect 55 37 61 39
rect 65 41 70 43
rect 41 35 51 37
rect 31 33 37 35
rect 31 31 33 33
rect 35 31 37 33
rect 49 31 51 35
rect 65 31 67 41
rect 75 35 77 46
rect 85 35 87 38
rect 31 29 44 31
rect 49 29 67 31
rect 71 33 77 35
rect 71 31 73 33
rect 75 31 77 33
rect 71 29 77 31
rect 81 33 87 35
rect 81 31 83 33
rect 85 31 87 33
rect 81 29 87 31
rect 42 26 44 29
rect 52 26 54 29
rect 28 16 34 18
rect 28 14 30 16
rect 32 14 34 16
rect 28 12 34 14
rect 61 25 67 29
rect 61 23 63 25
rect 65 23 67 25
rect 84 24 86 29
rect 61 21 67 23
rect 9 7 11 12
rect 19 9 21 12
rect 28 9 30 12
rect 19 7 30 9
rect 42 9 44 14
rect 52 9 54 14
rect 84 6 86 11
<< ndif >>
rect 4 18 9 26
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 12 19 22
rect 21 24 28 26
rect 21 22 24 24
rect 26 22 28 24
rect 21 20 28 22
rect 21 12 26 20
rect 36 14 42 26
rect 44 24 52 26
rect 44 22 47 24
rect 49 22 52 24
rect 44 14 52 22
rect 54 18 59 26
rect 77 22 84 24
rect 77 20 79 22
rect 81 20 84 22
rect 77 18 84 20
rect 54 14 62 18
rect 36 10 40 14
rect 34 7 40 10
rect 34 5 36 7
rect 38 5 40 7
rect 34 3 40 5
rect 56 7 62 14
rect 56 5 58 7
rect 60 5 62 7
rect 56 3 62 5
rect 79 11 84 18
rect 86 15 94 24
rect 86 13 89 15
rect 91 13 94 15
rect 86 11 94 13
<< pdif >>
rect 7 58 12 66
rect 5 56 12 58
rect 5 54 7 56
rect 9 54 12 56
rect 5 49 12 54
rect 5 47 7 49
rect 9 47 12 49
rect 5 45 12 47
rect 7 38 12 45
rect 14 38 19 66
rect 21 64 31 66
rect 21 62 25 64
rect 27 62 31 64
rect 21 46 31 62
rect 33 46 38 66
rect 40 50 48 66
rect 40 48 43 50
rect 45 48 48 50
rect 40 46 48 48
rect 50 57 58 66
rect 50 55 53 57
rect 55 55 58 57
rect 50 46 58 55
rect 60 57 68 66
rect 60 55 63 57
rect 65 55 68 57
rect 60 50 68 55
rect 60 48 63 50
rect 65 48 68 50
rect 60 46 68 48
rect 70 46 75 66
rect 77 64 85 66
rect 77 62 80 64
rect 82 62 85 64
rect 77 57 85 62
rect 77 55 80 57
rect 82 55 85 57
rect 77 46 85 55
rect 21 38 26 46
rect 80 38 85 46
rect 87 59 92 66
rect 87 57 94 59
rect 87 55 90 57
rect 92 55 94 57
rect 87 50 94 55
rect 87 48 90 50
rect 92 48 94 50
rect 87 46 94 48
rect 87 38 92 46
<< alu1 >>
rect -2 64 98 72
rect 2 50 10 51
rect 25 57 57 58
rect 25 55 53 57
rect 55 55 57 57
rect 25 54 57 55
rect 25 50 30 54
rect 2 49 30 50
rect 2 47 7 49
rect 9 47 30 49
rect 2 46 30 47
rect 2 25 6 46
rect 42 34 46 43
rect 73 42 79 50
rect 55 41 86 42
rect 55 39 57 41
rect 59 39 86 41
rect 55 38 86 39
rect 31 33 77 34
rect 31 31 33 33
rect 35 31 73 33
rect 75 31 77 33
rect 31 30 77 31
rect 82 33 86 38
rect 82 31 83 33
rect 85 31 86 33
rect 82 29 86 31
rect 57 25 71 26
rect 2 24 18 25
rect 2 22 14 24
rect 16 22 18 24
rect 2 21 18 22
rect 57 23 63 25
rect 65 23 71 25
rect 57 22 71 23
rect -2 7 98 8
rect -2 5 36 7
rect 38 5 58 7
rect 60 5 69 7
rect 71 5 98 7
rect -2 0 98 5
<< ptie >>
rect 67 7 73 18
rect 67 5 69 7
rect 71 5 73 7
rect 67 3 73 5
<< nmos >>
rect 9 12 11 26
rect 19 12 21 26
rect 42 14 44 26
rect 52 14 54 26
rect 84 11 86 24
<< pmos >>
rect 12 38 14 66
rect 19 38 21 66
rect 31 46 33 66
rect 38 46 40 66
rect 48 46 50 66
rect 58 46 60 66
rect 68 46 70 66
rect 75 46 77 66
rect 85 38 87 66
<< polyct0 >>
rect 11 31 13 33
rect 30 14 32 16
<< polyct1 >>
rect 57 39 59 41
rect 33 31 35 33
rect 73 31 75 33
rect 83 31 85 33
rect 63 23 65 25
<< ndifct0 >>
rect 4 14 6 16
rect 24 22 26 24
rect 47 22 49 24
rect 79 20 81 22
rect 89 13 91 15
<< ndifct1 >>
rect 14 22 16 24
rect 36 5 38 7
rect 58 5 60 7
<< ptiect1 >>
rect 69 5 71 7
<< pdifct0 >>
rect 7 54 9 56
rect 25 62 27 64
rect 43 48 45 50
rect 63 55 65 57
rect 63 48 65 50
rect 80 62 82 64
rect 80 55 82 57
rect 90 55 92 57
rect 90 48 92 50
<< pdifct1 >>
rect 7 47 9 49
rect 53 55 55 57
<< alu0 >>
rect 23 62 25 64
rect 27 62 29 64
rect 23 61 29 62
rect 78 62 80 64
rect 82 62 84 64
rect 6 56 10 58
rect 6 54 7 56
rect 9 54 10 56
rect 6 51 10 54
rect 62 57 67 59
rect 62 55 63 57
rect 65 55 67 57
rect 30 46 31 54
rect 62 51 67 55
rect 78 57 84 62
rect 78 55 80 57
rect 82 55 84 57
rect 78 54 84 55
rect 89 57 94 59
rect 89 55 90 57
rect 92 55 94 57
rect 34 50 67 51
rect 89 50 94 55
rect 34 48 43 50
rect 45 48 63 50
rect 65 48 67 50
rect 34 47 67 48
rect 34 42 38 47
rect 22 38 38 42
rect 22 34 26 38
rect 89 48 90 50
rect 92 48 94 50
rect 89 46 94 48
rect 9 33 26 34
rect 9 31 11 33
rect 13 31 26 33
rect 9 30 26 31
rect 22 25 26 30
rect 90 25 94 46
rect 22 24 51 25
rect 22 22 24 24
rect 26 22 47 24
rect 49 22 51 24
rect 78 22 94 25
rect 22 21 51 22
rect 78 20 79 22
rect 81 21 94 22
rect 81 20 82 21
rect 78 17 82 20
rect 2 16 82 17
rect 2 14 4 16
rect 6 14 30 16
rect 32 14 82 16
rect 2 13 82 14
rect 88 15 92 17
rect 88 13 89 15
rect 91 13 92 15
rect 88 8 92 13
<< labels >>
rlabel alu0 17 32 17 32 6 an
rlabel alu0 36 23 36 23 6 an
rlabel alu0 50 49 50 49 6 an
rlabel alu0 64 53 64 53 6 an
rlabel alu0 42 15 42 15 6 bn
rlabel alu0 80 19 80 19 6 bn
rlabel alu0 92 40 92 40 6 bn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 36 32 36 32 6 a1
rlabel alu1 44 36 44 36 6 a1
rlabel alu1 28 52 28 52 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 48 4 48 4 6 vss
rlabel alu1 52 32 52 32 6 a1
rlabel alu1 60 32 60 32 6 a1
rlabel alu1 68 32 68 32 6 a1
rlabel alu1 68 24 68 24 6 a2
rlabel alu1 60 24 60 24 6 a2
rlabel alu1 60 40 60 40 6 b
rlabel alu1 68 40 68 40 6 b
rlabel alu1 52 56 52 56 6 z
rlabel alu1 48 68 48 68 6 vdd
rlabel polyct1 84 32 84 32 6 b
rlabel alu1 76 44 76 44 6 b
<< end >>
