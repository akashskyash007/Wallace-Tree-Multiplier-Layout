magic
tech scmos
timestamp 1199543756
<< ab >>
rect 0 0 120 100
<< nwell >>
rect -5 48 125 105
<< pwell >>
rect -5 -5 125 48
<< poly >>
rect 13 94 15 98
rect 25 94 27 98
rect 37 85 39 89
rect 49 85 51 89
rect 61 85 63 89
rect 73 85 75 89
rect 87 85 89 89
rect 97 85 99 89
rect 107 85 109 89
rect 13 43 15 55
rect 25 43 27 55
rect 37 43 39 63
rect 49 43 51 63
rect 61 43 63 63
rect 73 43 75 61
rect 13 41 33 43
rect 13 39 29 41
rect 31 39 33 41
rect 13 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 67 41 75 43
rect 67 39 69 41
rect 71 39 75 41
rect 87 53 89 56
rect 97 53 99 56
rect 87 51 93 53
rect 87 49 89 51
rect 91 49 93 51
rect 87 47 93 49
rect 97 51 103 53
rect 97 49 99 51
rect 101 49 103 51
rect 97 47 103 49
rect 87 39 89 47
rect 97 39 99 47
rect 67 37 75 39
rect 83 37 89 39
rect 95 37 99 39
rect 107 43 109 55
rect 107 41 113 43
rect 107 39 109 41
rect 111 39 113 41
rect 107 37 113 39
rect 13 34 15 37
rect 25 34 27 37
rect 39 33 41 37
rect 49 33 51 37
rect 59 33 61 37
rect 71 29 73 37
rect 83 25 85 37
rect 95 25 97 37
rect 107 25 109 37
rect 13 10 15 14
rect 25 10 27 14
rect 39 13 41 17
rect 49 13 51 17
rect 59 13 61 17
rect 71 13 73 17
rect 83 13 85 17
rect 95 13 97 17
rect 107 13 109 17
<< ndif >>
rect 5 31 13 34
rect 5 29 7 31
rect 9 29 13 31
rect 5 21 13 29
rect 5 19 7 21
rect 9 19 13 21
rect 5 14 13 19
rect 15 31 25 34
rect 15 29 19 31
rect 21 29 25 31
rect 15 14 25 29
rect 27 33 37 34
rect 27 17 39 33
rect 41 17 49 33
rect 51 17 59 33
rect 61 29 66 33
rect 61 21 71 29
rect 61 19 65 21
rect 67 19 71 21
rect 61 17 71 19
rect 73 25 80 29
rect 73 21 83 25
rect 73 19 77 21
rect 79 19 83 21
rect 73 17 83 19
rect 85 17 95 25
rect 97 21 107 25
rect 97 19 101 21
rect 103 19 107 21
rect 97 17 107 19
rect 109 21 117 25
rect 109 19 113 21
rect 115 19 117 21
rect 109 17 117 19
rect 27 14 37 17
rect 31 11 37 14
rect 87 11 93 17
rect 31 9 33 11
rect 35 9 37 11
rect 31 7 37 9
rect 87 9 89 11
rect 91 9 93 11
rect 87 7 93 9
<< pdif >>
rect 5 91 13 94
rect 5 89 7 91
rect 9 89 13 91
rect 5 81 13 89
rect 5 79 7 81
rect 9 79 13 81
rect 5 71 13 79
rect 5 69 7 71
rect 9 69 13 71
rect 5 61 13 69
rect 5 59 7 61
rect 9 59 13 61
rect 5 55 13 59
rect 15 81 25 94
rect 15 79 19 81
rect 21 79 25 81
rect 15 71 25 79
rect 15 69 19 71
rect 21 69 25 71
rect 15 61 25 69
rect 15 59 19 61
rect 21 59 25 61
rect 15 55 25 59
rect 27 85 34 94
rect 53 91 59 93
rect 53 89 55 91
rect 57 89 59 91
rect 53 85 59 89
rect 27 81 37 85
rect 27 79 31 81
rect 33 79 37 81
rect 27 63 37 79
rect 39 81 49 85
rect 39 79 43 81
rect 45 79 49 81
rect 39 63 49 79
rect 51 63 61 85
rect 63 81 73 85
rect 63 79 67 81
rect 69 79 73 81
rect 63 63 73 79
rect 27 55 34 63
rect 66 61 73 63
rect 75 71 87 85
rect 75 69 79 71
rect 81 69 87 71
rect 75 61 87 69
rect 77 59 79 61
rect 81 59 87 61
rect 77 56 87 59
rect 89 56 97 85
rect 99 56 107 85
rect 102 55 107 56
rect 109 81 117 85
rect 109 79 113 81
rect 115 79 117 81
rect 109 55 117 79
<< alu1 >>
rect -2 95 122 100
rect -2 93 67 95
rect 69 93 79 95
rect 81 93 91 95
rect 93 93 103 95
rect 105 93 122 95
rect -2 91 122 93
rect -2 89 7 91
rect 9 89 55 91
rect 57 89 122 91
rect -2 88 122 89
rect 6 81 10 88
rect 6 79 7 81
rect 9 79 10 81
rect 6 71 10 79
rect 6 69 7 71
rect 9 69 10 71
rect 6 61 10 69
rect 6 59 7 61
rect 9 59 10 61
rect 6 57 10 59
rect 18 81 22 83
rect 18 79 19 81
rect 21 79 22 81
rect 18 71 22 79
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 77 34 79
rect 41 81 117 82
rect 41 79 43 81
rect 45 79 67 81
rect 69 79 113 81
rect 115 79 117 81
rect 41 78 117 79
rect 18 69 19 71
rect 21 69 22 71
rect 18 61 22 69
rect 18 59 19 61
rect 21 59 22 61
rect 6 31 10 33
rect 6 29 7 31
rect 9 29 10 31
rect 6 21 10 29
rect 6 19 7 21
rect 9 19 10 21
rect 6 12 10 19
rect 18 31 22 59
rect 18 29 19 31
rect 21 29 22 31
rect 18 17 22 29
rect 28 41 32 43
rect 28 39 29 41
rect 31 39 32 41
rect 28 22 32 39
rect 38 41 42 73
rect 38 39 39 41
rect 41 39 42 41
rect 38 27 42 39
rect 48 41 52 73
rect 48 39 49 41
rect 51 39 52 41
rect 48 27 52 39
rect 58 41 62 73
rect 58 39 59 41
rect 61 39 62 41
rect 58 37 62 39
rect 68 41 72 73
rect 68 39 69 41
rect 71 39 72 41
rect 68 37 72 39
rect 78 71 82 73
rect 78 69 79 71
rect 81 69 82 71
rect 78 61 82 69
rect 78 59 79 61
rect 81 59 82 61
rect 78 32 82 59
rect 64 28 82 32
rect 88 51 92 73
rect 88 49 89 51
rect 91 49 92 51
rect 64 22 68 28
rect 88 27 92 49
rect 98 51 102 73
rect 98 49 99 51
rect 101 49 102 51
rect 98 27 102 49
rect 108 41 112 73
rect 108 39 109 41
rect 111 39 112 41
rect 108 27 112 39
rect 28 21 68 22
rect 28 19 65 21
rect 67 19 68 21
rect 28 18 68 19
rect 75 21 105 22
rect 75 19 77 21
rect 79 19 101 21
rect 103 19 105 21
rect 75 18 105 19
rect 112 21 116 23
rect 112 19 113 21
rect 115 19 116 21
rect 64 17 68 18
rect 112 12 116 19
rect -2 11 122 12
rect -2 9 33 11
rect 35 9 89 11
rect 91 9 122 11
rect -2 7 45 9
rect 47 7 55 9
rect 57 7 65 9
rect 67 7 76 9
rect 78 7 103 9
rect 105 7 111 9
rect 113 7 122 9
rect -2 0 122 7
<< ptie >>
rect 43 9 80 11
rect 43 7 45 9
rect 47 7 55 9
rect 57 7 65 9
rect 67 7 76 9
rect 78 7 80 9
rect 101 9 115 11
rect 101 7 103 9
rect 105 7 111 9
rect 113 7 115 9
rect 43 5 80 7
rect 101 5 115 7
<< ntie >>
rect 65 95 107 97
rect 65 93 67 95
rect 69 93 79 95
rect 81 93 91 95
rect 93 93 103 95
rect 105 93 107 95
rect 65 91 107 93
<< nmos >>
rect 13 14 15 34
rect 25 14 27 34
rect 39 17 41 33
rect 49 17 51 33
rect 59 17 61 33
rect 71 17 73 29
rect 83 17 85 25
rect 95 17 97 25
rect 107 17 109 25
<< pmos >>
rect 13 55 15 94
rect 25 55 27 94
rect 37 63 39 85
rect 49 63 51 85
rect 61 63 63 85
rect 73 61 75 85
rect 87 56 89 85
rect 97 56 99 85
rect 107 55 109 85
<< polyct1 >>
rect 29 39 31 41
rect 39 39 41 41
rect 49 39 51 41
rect 59 39 61 41
rect 69 39 71 41
rect 89 49 91 51
rect 99 49 101 51
rect 109 39 111 41
<< ndifct1 >>
rect 7 29 9 31
rect 7 19 9 21
rect 19 29 21 31
rect 65 19 67 21
rect 77 19 79 21
rect 101 19 103 21
rect 113 19 115 21
rect 33 9 35 11
rect 89 9 91 11
<< ntiect1 >>
rect 67 93 69 95
rect 79 93 81 95
rect 91 93 93 95
rect 103 93 105 95
<< ptiect1 >>
rect 45 7 47 9
rect 55 7 57 9
rect 65 7 67 9
rect 76 7 78 9
rect 103 7 105 9
rect 111 7 113 9
<< pdifct1 >>
rect 7 89 9 91
rect 7 79 9 81
rect 7 69 9 71
rect 7 59 9 61
rect 19 79 21 81
rect 19 69 21 71
rect 19 59 21 61
rect 55 89 57 91
rect 31 79 33 81
rect 43 79 45 81
rect 67 79 69 81
rect 79 69 81 71
rect 79 59 81 61
rect 113 79 115 81
<< labels >>
rlabel alu1 20 50 20 50 6 q
rlabel alu1 50 50 50 50 6 i1
rlabel alu1 40 50 40 50 6 i0
rlabel alu1 60 6 60 6 6 vss
rlabel alu1 60 55 60 55 6 i2
rlabel alu1 70 55 70 55 6 i6
rlabel alu1 60 94 60 94 6 vdd
rlabel polyct1 100 50 100 50 6 i4
rlabel alu1 110 50 110 50 6 i5
rlabel polyct1 90 50 90 50 6 i3
<< end >>
