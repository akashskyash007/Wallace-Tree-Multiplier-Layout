magic
tech scmos
timestamp 1199544222
<< ab >>
rect 0 0 120 100
<< nwell >>
rect -5 48 125 105
<< pwell >>
rect -5 -5 125 48
<< poly >>
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 59 94 61 98
rect 11 76 13 80
rect 11 53 13 56
rect 23 53 25 56
rect 11 51 25 53
rect 35 53 37 56
rect 95 94 97 98
rect 107 94 109 98
rect 71 76 73 80
rect 35 51 43 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 3 41 9 43
rect 47 41 49 55
rect 59 43 61 55
rect 71 53 73 56
rect 67 51 73 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 95 43 97 55
rect 107 43 109 55
rect 3 39 5 41
rect 7 39 49 41
rect 3 37 9 39
rect 17 31 23 33
rect 17 29 19 31
rect 21 29 23 31
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 11 27 25 29
rect 11 24 13 27
rect 23 24 25 27
rect 35 27 43 29
rect 35 24 37 27
rect 47 25 49 39
rect 57 41 63 43
rect 77 41 83 43
rect 57 39 59 41
rect 61 39 79 41
rect 81 39 83 41
rect 57 37 63 39
rect 77 37 83 39
rect 87 41 109 43
rect 87 39 89 41
rect 91 39 109 41
rect 87 37 109 39
rect 67 31 73 33
rect 67 29 69 31
rect 71 29 73 31
rect 59 27 73 29
rect 11 10 13 14
rect 59 24 61 27
rect 71 24 73 27
rect 95 25 97 37
rect 107 25 109 37
rect 71 10 73 14
rect 23 2 25 6
rect 35 2 37 6
rect 47 2 49 6
rect 59 2 61 6
rect 95 2 97 6
rect 107 2 109 6
<< ndif >>
rect 42 24 47 25
rect 3 21 11 24
rect 3 19 5 21
rect 7 19 11 21
rect 3 14 11 19
rect 13 14 23 24
rect 15 11 23 14
rect 15 9 17 11
rect 19 9 23 11
rect 15 6 23 9
rect 25 6 35 24
rect 37 21 47 24
rect 37 19 41 21
rect 43 19 47 21
rect 37 6 47 19
rect 49 24 54 25
rect 75 31 83 33
rect 75 29 79 31
rect 81 29 83 31
rect 75 27 83 29
rect 75 24 81 27
rect 49 6 59 24
rect 61 14 71 24
rect 73 14 81 24
rect 90 21 95 25
rect 61 11 69 14
rect 61 9 65 11
rect 67 9 69 11
rect 87 11 95 21
rect 61 6 69 9
rect 87 9 89 11
rect 91 9 95 11
rect 87 6 95 9
rect 97 21 107 25
rect 97 19 101 21
rect 103 19 107 21
rect 97 6 107 19
rect 109 21 117 25
rect 109 19 113 21
rect 115 19 117 21
rect 109 11 117 19
rect 109 9 113 11
rect 115 9 117 11
rect 109 6 117 9
<< pdif >>
rect 15 91 23 94
rect 15 89 17 91
rect 19 89 23 91
rect 15 76 23 89
rect 3 71 11 76
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 56 11 59
rect 13 56 23 76
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 56 35 69
rect 37 71 47 94
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 42 55 47 56
rect 49 81 59 94
rect 49 79 53 81
rect 55 79 59 81
rect 49 71 59 79
rect 49 69 53 71
rect 55 69 59 71
rect 49 61 59 69
rect 49 59 53 61
rect 55 59 59 61
rect 49 55 59 59
rect 61 91 69 94
rect 61 89 65 91
rect 67 89 69 91
rect 61 76 69 89
rect 87 91 95 94
rect 87 89 89 91
rect 91 89 95 91
rect 87 81 95 89
rect 87 79 89 81
rect 91 79 95 81
rect 61 56 71 76
rect 73 61 81 76
rect 87 71 95 79
rect 87 69 89 71
rect 91 69 95 71
rect 87 67 95 69
rect 73 59 83 61
rect 73 57 79 59
rect 81 57 83 59
rect 73 56 83 57
rect 61 55 66 56
rect 77 55 83 56
rect 90 55 95 67
rect 97 81 107 94
rect 97 79 101 81
rect 103 79 107 81
rect 97 71 107 79
rect 97 69 101 71
rect 103 69 107 71
rect 97 61 107 69
rect 97 59 101 61
rect 103 59 107 61
rect 97 55 107 59
rect 109 91 117 94
rect 109 89 113 91
rect 115 89 117 91
rect 109 81 117 89
rect 109 79 113 81
rect 115 79 117 81
rect 109 71 117 79
rect 109 69 113 71
rect 115 69 117 71
rect 109 61 117 69
rect 109 59 113 61
rect 115 59 117 61
rect 109 55 117 59
<< alu1 >>
rect -2 95 122 100
rect -2 93 5 95
rect 7 93 77 95
rect 79 93 122 95
rect -2 91 122 93
rect -2 89 17 91
rect 19 89 65 91
rect 67 89 89 91
rect 91 89 113 91
rect 115 89 122 91
rect -2 88 122 89
rect 4 71 8 73
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 4 59 5 61
rect 7 59 8 61
rect 4 41 8 59
rect 4 39 5 41
rect 7 39 8 41
rect 4 21 8 39
rect 4 19 5 21
rect 7 19 8 21
rect 4 17 8 19
rect 18 51 22 83
rect 28 82 32 83
rect 52 82 56 83
rect 28 81 56 82
rect 28 79 29 81
rect 31 79 53 81
rect 55 79 56 81
rect 28 78 56 79
rect 28 71 32 78
rect 28 69 29 71
rect 31 69 32 71
rect 28 67 32 69
rect 40 71 44 73
rect 40 69 41 71
rect 43 69 44 71
rect 40 62 44 69
rect 18 49 19 51
rect 21 49 22 51
rect 18 31 22 49
rect 18 29 19 31
rect 21 29 22 31
rect 18 17 22 29
rect 28 58 44 62
rect 52 71 56 78
rect 52 69 53 71
rect 55 69 56 71
rect 52 61 56 69
rect 52 59 53 61
rect 55 59 56 61
rect 28 22 32 58
rect 52 57 56 59
rect 68 52 72 83
rect 88 81 92 88
rect 88 79 89 81
rect 91 79 92 81
rect 88 71 92 79
rect 88 69 89 71
rect 91 69 92 71
rect 88 67 92 69
rect 98 82 102 83
rect 98 81 105 82
rect 98 79 101 81
rect 103 79 105 81
rect 98 78 105 79
rect 112 81 116 88
rect 112 79 113 81
rect 115 79 116 81
rect 98 72 102 78
rect 98 71 105 72
rect 98 69 101 71
rect 103 69 105 71
rect 98 68 105 69
rect 112 71 116 79
rect 112 69 113 71
rect 115 69 116 71
rect 98 62 102 68
rect 98 61 105 62
rect 37 51 72 52
rect 37 49 39 51
rect 41 49 69 51
rect 71 49 72 51
rect 37 48 72 49
rect 48 41 63 42
rect 48 39 59 41
rect 61 39 63 41
rect 48 38 63 39
rect 48 32 52 38
rect 37 31 52 32
rect 37 29 39 31
rect 41 29 52 31
rect 37 28 52 29
rect 68 31 72 48
rect 68 29 69 31
rect 71 29 72 31
rect 68 27 72 29
rect 78 59 82 61
rect 78 57 79 59
rect 81 57 82 59
rect 78 41 82 57
rect 98 59 101 61
rect 103 59 105 61
rect 98 58 105 59
rect 112 61 116 69
rect 112 59 113 61
rect 115 59 116 61
rect 78 39 79 41
rect 81 39 82 41
rect 78 31 82 39
rect 78 29 79 31
rect 81 29 82 31
rect 78 27 82 29
rect 88 41 92 43
rect 88 39 89 41
rect 91 39 92 41
rect 88 22 92 39
rect 28 21 92 22
rect 28 19 41 21
rect 43 19 92 21
rect 28 18 92 19
rect 98 22 102 58
rect 112 57 116 59
rect 98 21 105 22
rect 98 19 101 21
rect 103 19 105 21
rect 98 18 105 19
rect 112 21 116 23
rect 112 19 113 21
rect 115 19 116 21
rect 98 17 102 18
rect 112 12 116 19
rect -2 11 122 12
rect -2 9 17 11
rect 19 9 65 11
rect 67 9 89 11
rect 91 9 113 11
rect 115 9 122 11
rect -2 0 122 9
<< ntie >>
rect 3 95 9 97
rect 3 93 5 95
rect 7 93 9 95
rect 75 95 81 97
rect 3 86 9 93
rect 75 93 77 95
rect 79 93 81 95
rect 75 86 81 93
<< nmos >>
rect 11 14 13 24
rect 23 6 25 24
rect 35 6 37 24
rect 47 6 49 25
rect 59 6 61 24
rect 71 14 73 24
rect 95 6 97 25
rect 107 6 109 25
<< pmos >>
rect 11 56 13 76
rect 23 56 25 94
rect 35 56 37 94
rect 47 55 49 94
rect 59 55 61 94
rect 71 56 73 76
rect 95 55 97 94
rect 107 55 109 94
<< polyct1 >>
rect 19 49 21 51
rect 39 49 41 51
rect 69 49 71 51
rect 5 39 7 41
rect 19 29 21 31
rect 39 29 41 31
rect 59 39 61 41
rect 79 39 81 41
rect 89 39 91 41
rect 69 29 71 31
<< ndifct1 >>
rect 5 19 7 21
rect 17 9 19 11
rect 41 19 43 21
rect 79 29 81 31
rect 65 9 67 11
rect 89 9 91 11
rect 101 19 103 21
rect 113 19 115 21
rect 113 9 115 11
<< ntiect1 >>
rect 5 93 7 95
rect 77 93 79 95
<< pdifct1 >>
rect 17 89 19 91
rect 5 69 7 71
rect 5 59 7 61
rect 29 79 31 81
rect 29 69 31 71
rect 41 69 43 71
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
rect 65 89 67 91
rect 89 89 91 91
rect 89 79 91 81
rect 89 69 91 71
rect 79 57 81 59
rect 101 79 103 81
rect 101 69 103 71
rect 101 59 103 61
rect 113 89 115 91
rect 113 79 115 81
rect 113 69 115 71
rect 113 59 115 61
<< labels >>
rlabel polyct1 20 50 20 50 6 i0
rlabel polyct1 40 50 40 50 6 i1
rlabel alu1 50 50 50 50 6 i1
rlabel alu1 60 6 60 6 6 vss
rlabel alu1 60 50 60 50 6 i1
rlabel alu1 70 55 70 55 6 i1
rlabel alu1 60 94 60 94 6 vdd
rlabel alu1 100 50 100 50 6 q
<< end >>
