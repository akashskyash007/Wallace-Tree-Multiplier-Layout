magic
tech scmos
timestamp 1635951023
<< ab >>
rect -290 77 -258 149
rect -254 77 -230 149
rect -226 77 -186 149
rect -131 77 -91 149
rect -87 77 -47 148
rect -43 77 -3 149
rect 10 77 50 149
rect 54 77 94 149
rect 97 77 137 149
rect -390 5 -262 77
rect -259 5 -131 77
rect -127 5 1 77
rect 5 5 69 77
rect -380 -66 -356 5
rect -354 -66 -290 5
rect -286 -66 -262 5
rect -258 -66 -194 5
rect -452 -140 -428 -68
rect -424 -139 -384 -67
rect -312 -138 -272 -66
rect -153 -67 -129 5
rect -126 -67 -62 5
rect 7 -67 47 5
rect -161 -139 -121 -67
rect -117 -139 -77 -67
rect -543 -212 -415 -140
rect -411 -212 -283 -140
rect -274 -211 -146 -139
rect -504 -284 -480 -212
rect -478 -284 -414 -212
rect -411 -284 -387 -212
rect -384 -284 -320 -212
rect -238 -283 -214 -211
rect -210 -283 -146 -211
rect -143 -211 -79 -139
rect -143 -283 -103 -211
rect -580 -355 -540 -284
rect -507 -355 -475 -284
rect -383 -355 -351 -284
rect -237 -353 -205 -283
rect -789 -498 -725 -426
rect -721 -427 -593 -355
rect -589 -427 -461 -355
rect -457 -427 -329 -355
rect -263 -425 -199 -353
rect -721 -498 -697 -427
rect -693 -499 -629 -427
rect -589 -499 -565 -427
rect -561 -499 -497 -427
rect -457 -498 -433 -427
rect -432 -498 -368 -427
rect -263 -496 -223 -425
<< nwell >>
rect -295 82 -181 117
rect -136 116 -86 117
rect -48 116 142 117
rect -136 82 142 116
rect -395 72 142 82
rect -395 37 74 72
rect -385 -55 -189 -26
rect -395 -62 -189 -55
rect -158 -62 -57 -27
rect -429 -63 -189 -62
rect -457 -71 -189 -63
rect -457 -107 -379 -71
rect -457 -108 -423 -107
rect -317 -106 -267 -71
rect -166 -72 -57 -62
rect 2 -72 52 -27
rect -166 -107 -72 -72
rect -278 -172 -74 -171
rect -548 -216 -74 -172
rect -548 -217 -278 -216
rect -509 -252 -315 -217
rect -585 -350 -535 -316
rect -243 -251 -98 -216
rect -512 -344 -470 -316
rect -512 -350 -445 -344
rect -388 -350 -346 -316
rect -242 -348 -200 -315
rect -726 -395 -324 -350
rect -268 -393 -194 -348
rect -794 -459 -692 -458
rect -794 -503 -624 -459
rect -698 -504 -624 -503
rect -594 -504 -492 -459
rect -462 -503 -363 -458
rect -268 -501 -218 -456
<< pwell >>
rect -295 117 -181 154
rect -136 153 -86 154
rect -48 153 142 154
rect -136 117 142 153
rect -86 116 -48 117
rect -395 0 74 37
rect -385 -26 -189 0
rect -158 -27 -57 0
rect -423 -108 -379 -107
rect -457 -135 -379 -108
rect -317 -107 -267 -106
rect 2 -27 52 0
rect -317 -135 -72 -107
rect -548 -144 -72 -135
rect -548 -171 -74 -144
rect -548 -172 -278 -171
rect -509 -279 -315 -252
rect -585 -316 -535 -279
rect -512 -289 -315 -279
rect -243 -288 -98 -251
rect -512 -316 -470 -289
rect -388 -316 -346 -289
rect -242 -315 -200 -288
rect -726 -421 -324 -395
rect -794 -432 -324 -421
rect -268 -430 -194 -393
rect -794 -458 -624 -432
rect -692 -459 -624 -458
rect -594 -459 -492 -432
rect -462 -458 -363 -432
rect -268 -456 -218 -430
<< poly >>
rect -281 142 -279 147
rect -274 142 -272 147
rect -245 132 -243 137
rect -217 134 -215 138
rect -204 136 -202 141
rect -197 136 -195 141
rect -281 120 -279 130
rect -274 127 -272 130
rect -274 125 -264 127
rect -270 123 -268 125
rect -266 123 -264 125
rect -122 134 -120 138
rect -109 136 -107 141
rect -102 136 -100 141
rect -78 133 -76 137
rect -65 135 -63 140
rect -58 135 -56 140
rect -270 121 -264 123
rect -281 118 -275 120
rect -281 116 -279 118
rect -277 116 -275 118
rect -281 114 -275 116
rect -280 106 -278 114
rect -270 106 -268 121
rect -245 120 -243 123
rect -217 120 -215 125
rect -204 120 -202 125
rect -245 118 -239 120
rect -245 116 -243 118
rect -241 116 -239 118
rect -245 114 -239 116
rect -217 118 -211 120
rect -217 116 -215 118
rect -213 116 -211 118
rect -217 114 -211 116
rect -207 118 -201 120
rect -207 116 -205 118
rect -203 116 -201 118
rect -207 114 -201 116
rect -245 111 -243 114
rect -217 110 -215 114
rect -280 87 -278 92
rect -270 88 -268 92
rect -245 88 -243 93
rect -207 103 -205 114
rect -197 112 -195 125
rect -122 120 -120 125
rect -109 120 -107 125
rect -122 118 -116 120
rect -122 116 -120 118
rect -118 116 -116 118
rect -122 114 -116 116
rect -112 118 -106 120
rect -112 116 -110 118
rect -108 116 -106 118
rect -112 114 -106 116
rect -197 110 -191 112
rect -122 110 -120 114
rect -197 108 -195 110
rect -193 108 -191 110
rect -197 106 -191 108
rect -197 103 -195 106
rect -217 88 -215 92
rect -112 103 -110 114
rect -102 112 -100 125
rect -34 134 -32 138
rect -21 136 -19 141
rect -14 136 -12 141
rect 19 134 21 138
rect 32 136 34 141
rect 39 136 41 141
rect 63 134 65 138
rect 76 136 78 141
rect 83 136 85 141
rect 106 134 108 138
rect 119 136 121 141
rect 126 136 128 141
rect -78 119 -76 124
rect -65 119 -63 124
rect -78 117 -72 119
rect -78 115 -76 117
rect -74 115 -72 117
rect -78 113 -72 115
rect -68 117 -62 119
rect -68 115 -66 117
rect -64 115 -62 117
rect -68 113 -62 115
rect -102 110 -96 112
rect -102 108 -100 110
rect -98 108 -96 110
rect -78 109 -76 113
rect -102 106 -96 108
rect -102 103 -100 106
rect -207 85 -205 90
rect -197 85 -195 90
rect -122 88 -120 92
rect -68 102 -66 113
rect -58 111 -56 124
rect -34 120 -32 125
rect -21 120 -19 125
rect -34 118 -28 120
rect -34 116 -32 118
rect -30 116 -28 118
rect -34 114 -28 116
rect -24 118 -18 120
rect -24 116 -22 118
rect -20 116 -18 118
rect -24 114 -18 116
rect -58 109 -52 111
rect -34 110 -32 114
rect -58 107 -56 109
rect -54 107 -52 109
rect -58 105 -52 107
rect -58 102 -56 105
rect -112 85 -110 90
rect -102 85 -100 90
rect -78 87 -76 91
rect -24 103 -22 114
rect -14 112 -12 125
rect 19 120 21 125
rect 32 120 34 125
rect 19 118 25 120
rect 19 116 21 118
rect 23 116 25 118
rect 19 114 25 116
rect 29 118 35 120
rect 29 116 31 118
rect 33 116 35 118
rect 29 114 35 116
rect -14 110 -8 112
rect 19 110 21 114
rect -14 108 -12 110
rect -10 108 -8 110
rect -14 106 -8 108
rect -14 103 -12 106
rect -68 84 -66 89
rect -58 84 -56 89
rect -34 88 -32 92
rect 29 103 31 114
rect 39 112 41 125
rect 63 120 65 125
rect 76 120 78 125
rect 63 118 69 120
rect 63 116 65 118
rect 67 116 69 118
rect 63 114 69 116
rect 73 118 79 120
rect 73 116 75 118
rect 77 116 79 118
rect 73 114 79 116
rect 39 110 45 112
rect 63 110 65 114
rect 39 108 41 110
rect 43 108 45 110
rect 39 106 45 108
rect 39 103 41 106
rect -24 85 -22 90
rect -14 85 -12 90
rect 19 88 21 92
rect 73 103 75 114
rect 83 112 85 125
rect 106 120 108 125
rect 119 120 121 125
rect 106 118 112 120
rect 106 116 108 118
rect 110 116 112 118
rect 106 114 112 116
rect 116 118 122 120
rect 116 116 118 118
rect 120 116 122 118
rect 116 114 122 116
rect 83 110 89 112
rect 106 110 108 114
rect 83 108 85 110
rect 87 108 89 110
rect 83 106 89 108
rect 83 103 85 106
rect 29 85 31 90
rect 39 85 41 90
rect 63 88 65 92
rect 116 103 118 114
rect 126 112 128 125
rect 126 110 132 112
rect 126 108 128 110
rect 130 108 132 110
rect 126 106 132 108
rect 126 103 128 106
rect 73 85 75 90
rect 83 85 85 90
rect 106 88 108 92
rect 116 85 118 90
rect 126 85 128 90
rect -381 71 -379 75
rect -371 71 -369 75
rect -361 71 -359 75
rect -351 71 -349 75
rect -341 71 -339 75
rect -321 71 -319 75
rect -311 71 -309 75
rect -301 71 -299 75
rect -351 54 -349 57
rect -341 54 -339 57
rect -351 52 -339 54
rect -345 50 -343 52
rect -341 50 -339 52
rect -345 48 -339 50
rect -250 71 -248 75
rect -240 71 -238 75
rect -230 71 -228 75
rect -220 71 -218 75
rect -210 71 -208 75
rect -190 71 -188 75
rect -180 71 -178 75
rect -170 71 -168 75
rect -290 64 -288 68
rect -280 64 -278 68
rect -290 47 -288 50
rect -280 47 -278 50
rect -290 45 -264 47
rect -381 40 -379 43
rect -371 40 -369 43
rect -361 40 -359 43
rect -321 40 -319 43
rect -311 40 -309 43
rect -381 38 -375 40
rect -381 36 -379 38
rect -377 36 -375 38
rect -381 34 -375 36
rect -371 38 -365 40
rect -361 38 -325 40
rect -371 36 -369 38
rect -367 36 -365 38
rect -371 34 -365 36
rect -380 25 -378 34
rect -371 30 -369 34
rect -353 30 -351 38
rect -331 36 -329 38
rect -327 36 -325 38
rect -331 34 -325 36
rect -321 38 -315 40
rect -321 36 -319 38
rect -317 36 -315 38
rect -321 34 -315 36
rect -311 38 -305 40
rect -311 36 -309 38
rect -307 36 -305 38
rect -301 39 -299 43
rect -301 37 -287 39
rect -311 34 -305 36
rect -293 35 -291 37
rect -289 35 -287 37
rect -341 32 -335 34
rect -341 30 -339 32
rect -337 30 -335 32
rect -373 28 -369 30
rect -373 25 -371 28
rect -363 25 -361 30
rect -341 28 -335 30
rect -341 25 -339 28
rect -318 25 -316 34
rect -311 25 -309 34
rect -293 33 -287 35
rect -291 30 -289 33
rect -280 31 -278 45
rect -270 43 -268 45
rect -266 43 -264 45
rect -220 54 -218 57
rect -210 54 -208 57
rect -220 52 -208 54
rect -214 50 -212 52
rect -210 50 -208 52
rect -214 48 -208 50
rect -118 71 -116 75
rect -108 71 -106 75
rect -98 71 -96 75
rect -88 71 -86 75
rect -78 71 -76 75
rect -58 71 -56 75
rect -48 71 -46 75
rect -38 71 -36 75
rect -159 64 -157 68
rect -149 64 -147 68
rect -159 47 -157 50
rect -149 47 -147 50
rect -159 45 -133 47
rect -270 41 -264 43
rect -250 40 -248 43
rect -240 40 -238 43
rect -230 40 -228 43
rect -190 40 -188 43
rect -180 40 -178 43
rect -250 38 -244 40
rect -250 36 -248 38
rect -246 36 -244 38
rect -250 34 -244 36
rect -240 38 -234 40
rect -230 38 -194 40
rect -240 36 -238 38
rect -236 36 -234 38
rect -240 34 -234 36
rect -301 25 -299 30
rect -353 13 -351 17
rect -380 7 -378 12
rect -373 7 -371 12
rect -363 9 -361 12
rect -341 9 -339 14
rect -363 7 -339 9
rect -249 25 -247 34
rect -240 30 -238 34
rect -222 30 -220 38
rect -200 36 -198 38
rect -196 36 -194 38
rect -200 34 -194 36
rect -190 38 -184 40
rect -190 36 -188 38
rect -186 36 -184 38
rect -190 34 -184 36
rect -180 38 -174 40
rect -180 36 -178 38
rect -176 36 -174 38
rect -170 39 -168 43
rect -170 37 -156 39
rect -180 34 -174 36
rect -162 35 -160 37
rect -158 35 -156 37
rect -210 32 -204 34
rect -210 30 -208 32
rect -206 30 -204 32
rect -242 28 -238 30
rect -242 25 -240 28
rect -232 25 -230 30
rect -291 13 -289 17
rect -318 7 -316 12
rect -311 7 -309 12
rect -301 9 -299 12
rect -280 9 -278 20
rect -301 7 -278 9
rect -210 28 -204 30
rect -210 25 -208 28
rect -187 25 -185 34
rect -180 25 -178 34
rect -162 33 -156 35
rect -160 30 -158 33
rect -149 31 -147 45
rect -139 43 -137 45
rect -135 43 -133 45
rect -88 54 -86 57
rect -78 54 -76 57
rect -88 52 -76 54
rect -82 50 -80 52
rect -78 50 -76 52
rect -82 48 -76 50
rect 22 71 24 75
rect -27 64 -25 68
rect -17 64 -15 68
rect -27 47 -25 50
rect -17 47 -15 50
rect -27 45 -1 47
rect -139 41 -133 43
rect -118 40 -116 43
rect -108 40 -106 43
rect -98 40 -96 43
rect -58 40 -56 43
rect -48 40 -46 43
rect -118 38 -112 40
rect -118 36 -116 38
rect -114 36 -112 38
rect -118 34 -112 36
rect -108 38 -102 40
rect -98 38 -62 40
rect -108 36 -106 38
rect -104 36 -102 38
rect -108 34 -102 36
rect -170 25 -168 30
rect -222 13 -220 17
rect -249 7 -247 12
rect -242 7 -240 12
rect -232 9 -230 12
rect -210 9 -208 14
rect -232 7 -208 9
rect -117 25 -115 34
rect -108 30 -106 34
rect -90 30 -88 38
rect -68 36 -66 38
rect -64 36 -62 38
rect -68 34 -62 36
rect -58 38 -52 40
rect -58 36 -56 38
rect -54 36 -52 38
rect -58 34 -52 36
rect -48 38 -42 40
rect -48 36 -46 38
rect -44 36 -42 38
rect -38 39 -36 43
rect -38 37 -24 39
rect -48 34 -42 36
rect -30 35 -28 37
rect -26 35 -24 37
rect -78 32 -72 34
rect -78 30 -76 32
rect -74 30 -72 32
rect -110 28 -106 30
rect -110 25 -108 28
rect -100 25 -98 30
rect -160 13 -158 17
rect -187 7 -185 12
rect -180 7 -178 12
rect -170 9 -168 12
rect -149 9 -147 20
rect -170 7 -147 9
rect -78 28 -72 30
rect -78 25 -76 28
rect -55 25 -53 34
rect -48 25 -46 34
rect -30 33 -24 35
rect -28 30 -26 33
rect -17 31 -15 45
rect -7 43 -5 45
rect -3 43 -1 45
rect -7 41 -1 43
rect 7 46 13 48
rect 7 44 9 46
rect 11 44 13 46
rect 58 71 60 75
rect 38 62 40 66
rect 48 62 50 66
rect 7 42 13 44
rect 11 41 13 42
rect 22 41 24 44
rect 38 41 40 44
rect 11 39 24 41
rect 30 39 40 41
rect 48 40 50 44
rect 58 41 60 44
rect 14 31 16 39
rect 30 35 32 39
rect 23 33 32 35
rect 44 38 50 40
rect 44 36 46 38
rect 48 36 50 38
rect 44 34 50 36
rect 54 39 60 41
rect 54 37 56 39
rect 58 37 60 39
rect 54 35 60 37
rect 23 31 25 33
rect 27 31 32 33
rect -38 25 -36 30
rect -90 13 -88 17
rect -117 7 -115 12
rect -110 7 -108 12
rect -100 9 -98 12
rect -78 9 -76 14
rect -100 7 -76 9
rect 23 29 32 31
rect 48 31 50 34
rect 30 26 32 29
rect 40 26 42 30
rect 48 29 52 31
rect 50 26 52 29
rect 57 26 59 35
rect -28 13 -26 17
rect -55 7 -53 12
rect -48 7 -46 12
rect -38 9 -36 12
rect -17 9 -15 20
rect 14 19 16 22
rect 14 17 19 19
rect -38 7 -15 9
rect 17 9 19 17
rect 30 13 32 17
rect 40 9 42 17
rect 50 9 52 14
rect 57 9 59 14
rect 17 7 42 9
rect -345 -6 -343 -1
rect -326 1 -304 3
rect -371 -11 -369 -6
rect -333 -8 -331 -3
rect -326 -8 -324 1
rect -316 -8 -314 -3
rect -306 -8 -304 1
rect -249 -6 -247 -1
rect -230 1 -208 3
rect -371 -23 -369 -20
rect -345 -23 -343 -18
rect -277 -11 -275 -6
rect -237 -8 -235 -3
rect -230 -8 -228 1
rect -220 -8 -218 -3
rect -210 -8 -208 1
rect -117 -7 -115 -2
rect -98 0 -76 2
rect -333 -23 -331 -20
rect -326 -23 -324 -20
rect -316 -23 -314 -20
rect -306 -23 -304 -20
rect -277 -23 -275 -20
rect -249 -23 -247 -18
rect -144 -12 -142 -7
rect -237 -23 -235 -20
rect -230 -23 -228 -20
rect -220 -23 -218 -20
rect -210 -23 -208 -20
rect -105 -9 -103 -4
rect -98 -9 -96 0
rect -88 -9 -86 -4
rect -78 -9 -76 0
rect -371 -25 -365 -23
rect -371 -27 -369 -25
rect -367 -27 -365 -25
rect -371 -29 -365 -27
rect -345 -25 -330 -23
rect -345 -27 -343 -25
rect -341 -27 -330 -25
rect -326 -26 -323 -23
rect -345 -29 -330 -27
rect -371 -32 -369 -29
rect -342 -32 -340 -29
rect -332 -32 -330 -29
rect -325 -32 -323 -26
rect -319 -25 -313 -23
rect -319 -27 -317 -25
rect -315 -27 -313 -25
rect -319 -29 -313 -27
rect -306 -25 -299 -23
rect -306 -27 -303 -25
rect -301 -27 -299 -25
rect -306 -29 -299 -27
rect -277 -25 -271 -23
rect -277 -27 -275 -25
rect -273 -27 -271 -25
rect -277 -29 -271 -27
rect -249 -25 -234 -23
rect -249 -27 -247 -25
rect -245 -27 -234 -25
rect -230 -26 -227 -23
rect -249 -29 -234 -27
rect -315 -32 -313 -29
rect -305 -32 -303 -29
rect -277 -32 -275 -29
rect -246 -32 -244 -29
rect -236 -32 -234 -29
rect -229 -32 -227 -26
rect -223 -25 -217 -23
rect -223 -27 -221 -25
rect -219 -27 -217 -25
rect -223 -29 -217 -27
rect -210 -25 -203 -23
rect -210 -27 -207 -25
rect -205 -27 -203 -25
rect -210 -29 -203 -27
rect -144 -24 -142 -21
rect -117 -24 -115 -19
rect 16 -10 18 -6
rect 29 -8 31 -3
rect 36 -8 38 -3
rect -105 -24 -103 -21
rect -98 -24 -96 -21
rect -88 -24 -86 -21
rect -78 -24 -76 -21
rect 16 -24 18 -19
rect 29 -24 31 -19
rect -144 -26 -138 -24
rect -144 -28 -142 -26
rect -140 -28 -138 -26
rect -219 -32 -217 -29
rect -209 -32 -207 -29
rect -144 -30 -138 -28
rect -117 -26 -102 -24
rect -117 -28 -115 -26
rect -113 -28 -102 -26
rect -98 -27 -95 -24
rect -117 -30 -102 -28
rect -371 -55 -369 -50
rect -277 -55 -275 -50
rect -144 -33 -142 -30
rect -114 -33 -112 -30
rect -104 -33 -102 -30
rect -97 -33 -95 -27
rect -91 -26 -85 -24
rect -91 -28 -89 -26
rect -87 -28 -85 -26
rect -91 -30 -85 -28
rect -78 -26 -71 -24
rect -78 -28 -75 -26
rect -73 -28 -71 -26
rect -78 -30 -71 -28
rect 16 -26 22 -24
rect 16 -28 18 -26
rect 20 -28 22 -26
rect 16 -30 22 -28
rect 26 -26 32 -24
rect 26 -28 28 -26
rect 30 -28 32 -26
rect 26 -30 32 -28
rect -87 -33 -85 -30
rect -77 -33 -75 -30
rect -144 -56 -142 -51
rect -342 -64 -340 -59
rect -332 -64 -330 -59
rect -325 -64 -323 -59
rect -315 -64 -313 -59
rect -305 -64 -303 -59
rect -246 -64 -244 -59
rect -236 -64 -234 -59
rect -229 -64 -227 -59
rect -219 -64 -217 -59
rect -209 -64 -207 -59
rect 16 -34 18 -30
rect 26 -41 28 -30
rect 36 -32 38 -19
rect 36 -34 42 -32
rect 36 -36 38 -34
rect 40 -36 42 -34
rect 36 -38 42 -36
rect 36 -41 38 -38
rect 16 -56 18 -52
rect 26 -59 28 -54
rect 36 -59 38 -54
rect -114 -65 -112 -60
rect -104 -65 -102 -60
rect -97 -65 -95 -60
rect -87 -65 -85 -60
rect -77 -65 -75 -60
rect -443 -84 -441 -79
rect -415 -82 -413 -78
rect -405 -80 -403 -75
rect -395 -80 -393 -75
rect -303 -81 -301 -77
rect -293 -79 -291 -74
rect -283 -79 -281 -74
rect -443 -105 -441 -102
rect -415 -104 -413 -100
rect -405 -104 -403 -93
rect -395 -96 -393 -93
rect -395 -98 -389 -96
rect -395 -100 -393 -98
rect -391 -100 -389 -98
rect -152 -82 -150 -78
rect -142 -80 -140 -75
rect -132 -80 -130 -75
rect -395 -102 -389 -100
rect -443 -107 -437 -105
rect -443 -109 -441 -107
rect -439 -109 -437 -107
rect -443 -111 -437 -109
rect -415 -106 -409 -104
rect -415 -108 -413 -106
rect -411 -108 -409 -106
rect -415 -110 -409 -108
rect -405 -106 -399 -104
rect -405 -108 -403 -106
rect -401 -108 -399 -106
rect -405 -110 -399 -108
rect -443 -114 -441 -111
rect -415 -115 -413 -110
rect -402 -115 -400 -110
rect -395 -115 -393 -102
rect -303 -103 -301 -99
rect -293 -103 -291 -92
rect -283 -95 -281 -92
rect -283 -97 -277 -95
rect -283 -99 -281 -97
rect -279 -99 -277 -97
rect -283 -101 -277 -99
rect -108 -82 -106 -78
rect -98 -80 -96 -75
rect -88 -80 -86 -75
rect -303 -105 -297 -103
rect -303 -107 -301 -105
rect -299 -107 -297 -105
rect -303 -109 -297 -107
rect -293 -105 -287 -103
rect -293 -107 -291 -105
rect -289 -107 -287 -105
rect -293 -109 -287 -107
rect -303 -114 -301 -109
rect -290 -114 -288 -109
rect -283 -114 -281 -101
rect -152 -104 -150 -100
rect -142 -104 -140 -93
rect -132 -96 -130 -93
rect -132 -98 -126 -96
rect -132 -100 -130 -98
rect -128 -100 -126 -98
rect -132 -102 -126 -100
rect -152 -106 -146 -104
rect -152 -108 -150 -106
rect -148 -108 -146 -106
rect -152 -110 -146 -108
rect -142 -106 -136 -104
rect -142 -108 -140 -106
rect -138 -108 -136 -106
rect -142 -110 -136 -108
rect -443 -128 -441 -123
rect -415 -128 -413 -124
rect -402 -131 -400 -126
rect -395 -131 -393 -126
rect -303 -127 -301 -123
rect -152 -115 -150 -110
rect -139 -115 -137 -110
rect -132 -115 -130 -102
rect -108 -104 -106 -100
rect -98 -104 -96 -93
rect -88 -96 -86 -93
rect -88 -98 -82 -96
rect -88 -100 -86 -98
rect -84 -100 -82 -98
rect -88 -102 -82 -100
rect -108 -106 -102 -104
rect -108 -108 -106 -106
rect -104 -108 -102 -106
rect -108 -110 -102 -108
rect -98 -106 -92 -104
rect -98 -108 -96 -106
rect -94 -108 -92 -106
rect -98 -110 -92 -108
rect -108 -115 -106 -110
rect -95 -115 -93 -110
rect -88 -115 -86 -102
rect -290 -130 -288 -125
rect -283 -130 -281 -125
rect -152 -128 -150 -124
rect -139 -131 -137 -126
rect -132 -131 -130 -126
rect -108 -128 -106 -124
rect -95 -131 -93 -126
rect -88 -131 -86 -126
rect -533 -147 -531 -142
rect -526 -147 -524 -142
rect -516 -144 -492 -142
rect -516 -147 -514 -144
rect -506 -152 -504 -148
rect -494 -149 -492 -144
rect -471 -147 -469 -142
rect -464 -147 -462 -142
rect -454 -144 -431 -142
rect -454 -147 -452 -144
rect -533 -169 -531 -160
rect -526 -163 -524 -160
rect -526 -165 -522 -163
rect -516 -165 -514 -160
rect -444 -152 -442 -148
rect -494 -163 -492 -160
rect -494 -165 -488 -163
rect -524 -169 -522 -165
rect -534 -171 -528 -169
rect -534 -173 -532 -171
rect -530 -173 -528 -171
rect -534 -175 -528 -173
rect -524 -171 -518 -169
rect -524 -173 -522 -171
rect -520 -173 -518 -171
rect -506 -173 -504 -165
rect -494 -167 -492 -165
rect -490 -167 -488 -165
rect -494 -169 -488 -167
rect -471 -169 -469 -160
rect -464 -169 -462 -160
rect -454 -165 -452 -160
rect -433 -155 -431 -144
rect -401 -147 -399 -142
rect -394 -147 -392 -142
rect -384 -144 -360 -142
rect -384 -147 -382 -144
rect -444 -168 -442 -165
rect -374 -152 -372 -148
rect -362 -149 -360 -144
rect -339 -147 -337 -142
rect -332 -147 -330 -142
rect -322 -144 -299 -142
rect -322 -147 -320 -144
rect -484 -171 -478 -169
rect -484 -173 -482 -171
rect -480 -173 -478 -171
rect -524 -175 -518 -173
rect -514 -175 -478 -173
rect -474 -171 -468 -169
rect -474 -173 -472 -171
rect -470 -173 -468 -171
rect -474 -175 -468 -173
rect -464 -171 -458 -169
rect -464 -173 -462 -171
rect -460 -173 -458 -171
rect -446 -170 -440 -168
rect -446 -172 -444 -170
rect -442 -172 -440 -170
rect -464 -175 -458 -173
rect -454 -174 -440 -172
rect -534 -178 -532 -175
rect -524 -178 -522 -175
rect -514 -178 -512 -175
rect -474 -178 -472 -175
rect -464 -178 -462 -175
rect -454 -178 -452 -174
rect -498 -185 -492 -183
rect -498 -187 -496 -185
rect -494 -187 -492 -185
rect -504 -189 -492 -187
rect -504 -192 -502 -189
rect -494 -192 -492 -189
rect -433 -180 -431 -166
rect -401 -169 -399 -160
rect -394 -163 -392 -160
rect -394 -165 -390 -163
rect -384 -165 -382 -160
rect -312 -152 -310 -148
rect -362 -163 -360 -160
rect -362 -165 -356 -163
rect -392 -169 -390 -165
rect -402 -171 -396 -169
rect -402 -173 -400 -171
rect -398 -173 -396 -171
rect -402 -175 -396 -173
rect -392 -171 -386 -169
rect -392 -173 -390 -171
rect -388 -173 -386 -171
rect -374 -173 -372 -165
rect -362 -167 -360 -165
rect -358 -167 -356 -165
rect -362 -169 -356 -167
rect -339 -169 -337 -160
rect -332 -169 -330 -160
rect -322 -165 -320 -160
rect -301 -155 -299 -144
rect -264 -146 -262 -141
rect -257 -146 -255 -141
rect -247 -143 -223 -141
rect -247 -146 -245 -143
rect -312 -168 -310 -165
rect -237 -151 -235 -147
rect -225 -148 -223 -143
rect -202 -146 -200 -141
rect -195 -146 -193 -141
rect -185 -143 -162 -141
rect -185 -146 -183 -143
rect -352 -171 -346 -169
rect -352 -173 -350 -171
rect -348 -173 -346 -171
rect -392 -175 -386 -173
rect -382 -175 -346 -173
rect -342 -171 -336 -169
rect -342 -173 -340 -171
rect -338 -173 -336 -171
rect -342 -175 -336 -173
rect -332 -171 -326 -169
rect -332 -173 -330 -171
rect -328 -173 -326 -171
rect -314 -170 -308 -168
rect -314 -172 -312 -170
rect -310 -172 -308 -170
rect -332 -175 -326 -173
rect -322 -174 -308 -172
rect -423 -178 -417 -176
rect -402 -178 -400 -175
rect -392 -178 -390 -175
rect -382 -178 -380 -175
rect -342 -178 -340 -175
rect -332 -178 -330 -175
rect -322 -178 -320 -174
rect -423 -180 -421 -178
rect -419 -180 -417 -178
rect -443 -182 -417 -180
rect -443 -185 -441 -182
rect -433 -185 -431 -182
rect -443 -203 -441 -199
rect -433 -203 -431 -199
rect -534 -210 -532 -206
rect -524 -210 -522 -206
rect -514 -210 -512 -206
rect -504 -210 -502 -206
rect -494 -210 -492 -206
rect -474 -210 -472 -206
rect -464 -210 -462 -206
rect -454 -210 -452 -206
rect -366 -185 -360 -183
rect -366 -187 -364 -185
rect -362 -187 -360 -185
rect -372 -189 -360 -187
rect -372 -192 -370 -189
rect -362 -192 -360 -189
rect -301 -180 -299 -166
rect -264 -168 -262 -159
rect -257 -162 -255 -159
rect -257 -164 -253 -162
rect -247 -164 -245 -159
rect -175 -151 -173 -147
rect -225 -162 -223 -159
rect -225 -164 -219 -162
rect -255 -168 -253 -164
rect -265 -170 -259 -168
rect -265 -172 -263 -170
rect -261 -172 -259 -170
rect -265 -174 -259 -172
rect -255 -170 -249 -168
rect -255 -172 -253 -170
rect -251 -172 -249 -170
rect -237 -172 -235 -164
rect -225 -166 -223 -164
rect -221 -166 -219 -164
rect -225 -168 -219 -166
rect -202 -168 -200 -159
rect -195 -168 -193 -159
rect -185 -164 -183 -159
rect -164 -154 -162 -143
rect -116 -143 -91 -141
rect -133 -148 -131 -143
rect -126 -148 -124 -143
rect -175 -167 -173 -164
rect -116 -151 -114 -143
rect -106 -151 -104 -147
rect -93 -151 -91 -143
rect -93 -153 -88 -151
rect -90 -156 -88 -153
rect -215 -170 -209 -168
rect -215 -172 -213 -170
rect -211 -172 -209 -170
rect -255 -174 -249 -172
rect -245 -174 -209 -172
rect -205 -170 -199 -168
rect -205 -172 -203 -170
rect -201 -172 -199 -170
rect -205 -174 -199 -172
rect -195 -170 -189 -168
rect -195 -172 -193 -170
rect -191 -172 -189 -170
rect -177 -169 -171 -167
rect -177 -171 -175 -169
rect -173 -171 -171 -169
rect -195 -174 -189 -172
rect -185 -173 -171 -171
rect -291 -178 -285 -176
rect -265 -177 -263 -174
rect -255 -177 -253 -174
rect -245 -177 -243 -174
rect -205 -177 -203 -174
rect -195 -177 -193 -174
rect -185 -177 -183 -173
rect -291 -180 -289 -178
rect -287 -180 -285 -178
rect -311 -182 -285 -180
rect -311 -185 -309 -182
rect -301 -185 -299 -182
rect -311 -203 -309 -199
rect -301 -203 -299 -199
rect -229 -184 -223 -182
rect -229 -186 -227 -184
rect -225 -186 -223 -184
rect -235 -188 -223 -186
rect -235 -191 -233 -188
rect -225 -191 -223 -188
rect -164 -179 -162 -165
rect -133 -169 -131 -160
rect -126 -163 -124 -160
rect -126 -165 -122 -163
rect -116 -164 -114 -160
rect -106 -163 -104 -160
rect -124 -168 -122 -165
rect -106 -165 -97 -163
rect -106 -167 -101 -165
rect -99 -167 -97 -165
rect -134 -171 -128 -169
rect -134 -173 -132 -171
rect -130 -173 -128 -171
rect -134 -175 -128 -173
rect -124 -170 -118 -168
rect -124 -172 -122 -170
rect -120 -172 -118 -170
rect -124 -174 -118 -172
rect -106 -169 -97 -167
rect -106 -173 -104 -169
rect -90 -173 -88 -165
rect -154 -177 -148 -175
rect -154 -179 -152 -177
rect -150 -179 -148 -177
rect -134 -178 -132 -175
rect -124 -178 -122 -174
rect -114 -175 -104 -173
rect -98 -175 -85 -173
rect -114 -178 -112 -175
rect -98 -178 -96 -175
rect -87 -176 -85 -175
rect -87 -178 -81 -176
rect -174 -181 -148 -179
rect -174 -184 -172 -181
rect -164 -184 -162 -181
rect -174 -202 -172 -198
rect -164 -202 -162 -198
rect -402 -210 -400 -206
rect -392 -210 -390 -206
rect -382 -210 -380 -206
rect -372 -210 -370 -206
rect -362 -210 -360 -206
rect -342 -210 -340 -206
rect -332 -210 -330 -206
rect -322 -210 -320 -206
rect -265 -209 -263 -205
rect -255 -209 -253 -205
rect -245 -209 -243 -205
rect -235 -209 -233 -205
rect -225 -209 -223 -205
rect -205 -209 -203 -205
rect -195 -209 -193 -205
rect -185 -209 -183 -205
rect -124 -200 -122 -196
rect -114 -200 -112 -196
rect -134 -209 -132 -205
rect -87 -180 -85 -178
rect -83 -180 -81 -178
rect -87 -182 -81 -180
rect -98 -209 -96 -205
rect -466 -219 -464 -214
rect -456 -219 -454 -214
rect -449 -219 -447 -214
rect -439 -219 -437 -214
rect -429 -219 -427 -214
rect -372 -219 -370 -214
rect -362 -219 -360 -214
rect -355 -219 -353 -214
rect -345 -219 -343 -214
rect -335 -219 -333 -214
rect -198 -218 -196 -213
rect -188 -218 -186 -213
rect -181 -218 -179 -213
rect -171 -218 -169 -213
rect -161 -218 -159 -213
rect -495 -228 -493 -223
rect -402 -228 -400 -223
rect -229 -227 -227 -222
rect -134 -226 -132 -222
rect -124 -224 -122 -219
rect -114 -224 -112 -219
rect -495 -249 -493 -246
rect -466 -249 -464 -246
rect -456 -249 -454 -246
rect -495 -251 -489 -249
rect -495 -253 -493 -251
rect -491 -253 -489 -251
rect -495 -255 -489 -253
rect -469 -251 -454 -249
rect -469 -253 -467 -251
rect -465 -253 -454 -251
rect -449 -252 -447 -246
rect -439 -249 -437 -246
rect -429 -249 -427 -246
rect -402 -249 -400 -246
rect -372 -249 -370 -246
rect -362 -249 -360 -246
rect -469 -255 -454 -253
rect -450 -255 -447 -252
rect -443 -251 -437 -249
rect -443 -253 -441 -251
rect -439 -253 -437 -251
rect -443 -255 -437 -253
rect -430 -251 -423 -249
rect -430 -253 -427 -251
rect -425 -253 -423 -251
rect -430 -255 -423 -253
rect -402 -251 -396 -249
rect -402 -253 -400 -251
rect -398 -253 -396 -251
rect -402 -255 -396 -253
rect -375 -251 -360 -249
rect -375 -253 -373 -251
rect -371 -253 -360 -251
rect -355 -252 -353 -246
rect -345 -249 -343 -246
rect -335 -249 -333 -246
rect -229 -248 -227 -245
rect -198 -248 -196 -245
rect -188 -248 -186 -245
rect -375 -255 -360 -253
rect -356 -255 -353 -252
rect -349 -251 -343 -249
rect -349 -253 -347 -251
rect -345 -253 -343 -251
rect -349 -255 -343 -253
rect -336 -251 -329 -249
rect -336 -253 -333 -251
rect -331 -253 -329 -251
rect -336 -255 -329 -253
rect -229 -250 -223 -248
rect -229 -252 -227 -250
rect -225 -252 -223 -250
rect -229 -254 -223 -252
rect -201 -250 -186 -248
rect -201 -252 -199 -250
rect -197 -252 -186 -250
rect -181 -251 -179 -245
rect -171 -248 -169 -245
rect -161 -248 -159 -245
rect -134 -248 -132 -244
rect -124 -248 -122 -237
rect -114 -240 -112 -237
rect -114 -242 -108 -240
rect -114 -244 -112 -242
rect -110 -244 -108 -242
rect -114 -246 -108 -244
rect -201 -254 -186 -252
rect -182 -254 -179 -251
rect -175 -250 -169 -248
rect -175 -252 -173 -250
rect -171 -252 -169 -250
rect -175 -254 -169 -252
rect -162 -250 -155 -248
rect -162 -252 -159 -250
rect -157 -252 -155 -250
rect -162 -254 -155 -252
rect -134 -250 -128 -248
rect -134 -252 -132 -250
rect -130 -252 -128 -250
rect -134 -254 -128 -252
rect -124 -250 -118 -248
rect -124 -252 -122 -250
rect -120 -252 -118 -250
rect -124 -254 -118 -252
rect -495 -258 -493 -255
rect -469 -260 -467 -255
rect -457 -258 -455 -255
rect -450 -258 -448 -255
rect -440 -258 -438 -255
rect -430 -258 -428 -255
rect -402 -258 -400 -255
rect -495 -272 -493 -267
rect -375 -260 -373 -255
rect -363 -258 -361 -255
rect -356 -258 -354 -255
rect -346 -258 -344 -255
rect -336 -258 -334 -255
rect -229 -257 -227 -254
rect -469 -277 -467 -272
rect -457 -275 -455 -270
rect -450 -279 -448 -270
rect -440 -275 -438 -270
rect -430 -279 -428 -270
rect -402 -272 -400 -267
rect -201 -259 -199 -254
rect -189 -257 -187 -254
rect -182 -257 -180 -254
rect -172 -257 -170 -254
rect -162 -257 -160 -254
rect -450 -281 -428 -279
rect -375 -277 -373 -272
rect -363 -275 -361 -270
rect -356 -279 -354 -270
rect -346 -275 -344 -270
rect -336 -279 -334 -270
rect -229 -271 -227 -266
rect -134 -259 -132 -254
rect -121 -259 -119 -254
rect -114 -259 -112 -246
rect -356 -281 -334 -279
rect -201 -276 -199 -271
rect -189 -274 -187 -269
rect -182 -278 -180 -269
rect -172 -274 -170 -269
rect -162 -278 -160 -269
rect -134 -272 -132 -268
rect -182 -280 -160 -278
rect -121 -275 -119 -270
rect -114 -275 -112 -270
rect -498 -291 -496 -286
rect -491 -291 -489 -286
rect -374 -291 -372 -286
rect -367 -291 -365 -286
rect -228 -290 -226 -285
rect -221 -290 -219 -285
rect -571 -299 -569 -295
rect -558 -297 -556 -292
rect -551 -297 -549 -292
rect -571 -313 -569 -308
rect -558 -313 -556 -308
rect -571 -315 -565 -313
rect -571 -317 -569 -315
rect -567 -317 -565 -315
rect -571 -319 -565 -317
rect -561 -315 -555 -313
rect -561 -317 -559 -315
rect -557 -317 -555 -315
rect -561 -319 -555 -317
rect -571 -323 -569 -319
rect -561 -330 -559 -319
rect -551 -321 -549 -308
rect -498 -313 -496 -303
rect -491 -306 -489 -303
rect -491 -308 -481 -306
rect -487 -310 -485 -308
rect -483 -310 -481 -308
rect -487 -312 -481 -310
rect -498 -315 -492 -313
rect -498 -317 -496 -315
rect -494 -317 -492 -315
rect -498 -319 -492 -317
rect -551 -323 -545 -321
rect -551 -325 -549 -323
rect -547 -325 -545 -323
rect -551 -327 -545 -325
rect -497 -327 -495 -319
rect -487 -327 -485 -312
rect -374 -313 -372 -303
rect -367 -306 -365 -303
rect -367 -308 -357 -306
rect -363 -310 -361 -308
rect -359 -310 -357 -308
rect -363 -312 -357 -310
rect -228 -312 -226 -302
rect -221 -305 -219 -302
rect -221 -307 -211 -305
rect -217 -309 -215 -307
rect -213 -309 -211 -307
rect -217 -311 -211 -309
rect -374 -315 -368 -313
rect -374 -317 -372 -315
rect -370 -317 -368 -315
rect -374 -319 -368 -317
rect -373 -327 -371 -319
rect -363 -327 -361 -312
rect -228 -314 -222 -312
rect -228 -316 -226 -314
rect -224 -316 -222 -314
rect -228 -318 -222 -316
rect -227 -326 -225 -318
rect -217 -326 -215 -311
rect -551 -330 -549 -327
rect -571 -345 -569 -341
rect -561 -348 -559 -343
rect -551 -348 -549 -343
rect -497 -346 -495 -341
rect -487 -345 -485 -341
rect -373 -346 -371 -341
rect -363 -345 -361 -341
rect -227 -345 -225 -340
rect -217 -344 -215 -340
rect -712 -361 -710 -357
rect -702 -361 -700 -357
rect -692 -361 -690 -357
rect -682 -361 -680 -357
rect -672 -361 -670 -357
rect -652 -361 -650 -357
rect -642 -361 -640 -357
rect -632 -361 -630 -357
rect -682 -378 -680 -375
rect -672 -378 -670 -375
rect -682 -380 -670 -378
rect -676 -382 -674 -380
rect -672 -382 -670 -380
rect -676 -384 -670 -382
rect -580 -361 -578 -357
rect -570 -361 -568 -357
rect -560 -361 -558 -357
rect -550 -361 -548 -357
rect -540 -361 -538 -357
rect -520 -361 -518 -357
rect -510 -361 -508 -357
rect -500 -361 -498 -357
rect -621 -368 -619 -364
rect -611 -368 -609 -364
rect -621 -385 -619 -382
rect -611 -385 -609 -382
rect -621 -387 -595 -385
rect -712 -392 -710 -389
rect -702 -392 -700 -389
rect -692 -392 -690 -389
rect -652 -392 -650 -389
rect -642 -392 -640 -389
rect -712 -394 -706 -392
rect -712 -396 -710 -394
rect -708 -396 -706 -394
rect -712 -398 -706 -396
rect -702 -394 -696 -392
rect -692 -394 -656 -392
rect -702 -396 -700 -394
rect -698 -396 -696 -394
rect -702 -398 -696 -396
rect -711 -407 -709 -398
rect -702 -402 -700 -398
rect -684 -402 -682 -394
rect -662 -396 -660 -394
rect -658 -396 -656 -394
rect -662 -398 -656 -396
rect -652 -394 -646 -392
rect -652 -396 -650 -394
rect -648 -396 -646 -394
rect -652 -398 -646 -396
rect -642 -394 -636 -392
rect -642 -396 -640 -394
rect -638 -396 -636 -394
rect -632 -393 -630 -389
rect -632 -395 -618 -393
rect -642 -398 -636 -396
rect -624 -397 -622 -395
rect -620 -397 -618 -395
rect -672 -400 -666 -398
rect -672 -402 -670 -400
rect -668 -402 -666 -400
rect -704 -404 -700 -402
rect -704 -407 -702 -404
rect -694 -407 -692 -402
rect -672 -404 -666 -402
rect -672 -407 -670 -404
rect -649 -407 -647 -398
rect -642 -407 -640 -398
rect -624 -399 -618 -397
rect -622 -402 -620 -399
rect -611 -401 -609 -387
rect -601 -389 -599 -387
rect -597 -389 -595 -387
rect -550 -378 -548 -375
rect -540 -378 -538 -375
rect -550 -380 -538 -378
rect -544 -382 -542 -380
rect -540 -382 -538 -380
rect -544 -384 -538 -382
rect -448 -361 -446 -357
rect -438 -361 -436 -357
rect -428 -361 -426 -357
rect -418 -361 -416 -357
rect -408 -361 -406 -357
rect -388 -361 -386 -357
rect -378 -361 -376 -357
rect -368 -361 -366 -357
rect -246 -359 -244 -355
rect -489 -368 -487 -364
rect -479 -368 -477 -364
rect -489 -385 -487 -382
rect -479 -385 -477 -382
rect -489 -387 -463 -385
rect -601 -391 -595 -389
rect -580 -392 -578 -389
rect -570 -392 -568 -389
rect -560 -392 -558 -389
rect -520 -392 -518 -389
rect -510 -392 -508 -389
rect -580 -394 -574 -392
rect -580 -396 -578 -394
rect -576 -396 -574 -394
rect -580 -398 -574 -396
rect -570 -394 -564 -392
rect -560 -394 -524 -392
rect -570 -396 -568 -394
rect -566 -396 -564 -394
rect -570 -398 -564 -396
rect -632 -407 -630 -402
rect -684 -419 -682 -415
rect -711 -425 -709 -420
rect -704 -425 -702 -420
rect -694 -423 -692 -420
rect -672 -423 -670 -418
rect -694 -425 -670 -423
rect -579 -407 -577 -398
rect -570 -402 -568 -398
rect -552 -402 -550 -394
rect -530 -396 -528 -394
rect -526 -396 -524 -394
rect -530 -398 -524 -396
rect -520 -394 -514 -392
rect -520 -396 -518 -394
rect -516 -396 -514 -394
rect -520 -398 -514 -396
rect -510 -394 -504 -392
rect -510 -396 -508 -394
rect -506 -396 -504 -394
rect -500 -393 -498 -389
rect -500 -395 -486 -393
rect -510 -398 -504 -396
rect -492 -397 -490 -395
rect -488 -397 -486 -395
rect -540 -400 -534 -398
rect -540 -402 -538 -400
rect -536 -402 -534 -400
rect -572 -404 -568 -402
rect -572 -407 -570 -404
rect -562 -407 -560 -402
rect -622 -419 -620 -415
rect -649 -425 -647 -420
rect -642 -425 -640 -420
rect -632 -423 -630 -420
rect -611 -423 -609 -412
rect -632 -425 -609 -423
rect -540 -404 -534 -402
rect -540 -407 -538 -404
rect -517 -407 -515 -398
rect -510 -407 -508 -398
rect -492 -399 -486 -397
rect -490 -402 -488 -399
rect -479 -401 -477 -387
rect -469 -389 -467 -387
rect -465 -389 -463 -387
rect -418 -378 -416 -375
rect -408 -378 -406 -375
rect -418 -380 -406 -378
rect -412 -382 -410 -380
rect -408 -382 -406 -380
rect -412 -384 -406 -382
rect -357 -368 -355 -364
rect -347 -368 -345 -364
rect -357 -385 -355 -382
rect -347 -385 -345 -382
rect -261 -384 -255 -382
rect -357 -387 -331 -385
rect -469 -391 -463 -389
rect -448 -392 -446 -389
rect -438 -392 -436 -389
rect -428 -392 -426 -389
rect -388 -392 -386 -389
rect -378 -392 -376 -389
rect -448 -394 -442 -392
rect -448 -396 -446 -394
rect -444 -396 -442 -394
rect -448 -398 -442 -396
rect -438 -394 -432 -392
rect -428 -394 -392 -392
rect -438 -396 -436 -394
rect -434 -396 -432 -394
rect -438 -398 -432 -396
rect -500 -407 -498 -402
rect -552 -419 -550 -415
rect -579 -425 -577 -420
rect -572 -425 -570 -420
rect -562 -423 -560 -420
rect -540 -423 -538 -418
rect -562 -425 -538 -423
rect -447 -407 -445 -398
rect -438 -402 -436 -398
rect -420 -402 -418 -394
rect -398 -396 -396 -394
rect -394 -396 -392 -394
rect -398 -398 -392 -396
rect -388 -394 -382 -392
rect -388 -396 -386 -394
rect -384 -396 -382 -394
rect -388 -398 -382 -396
rect -378 -394 -372 -392
rect -378 -396 -376 -394
rect -374 -396 -372 -394
rect -368 -393 -366 -389
rect -368 -395 -354 -393
rect -378 -398 -372 -396
rect -360 -397 -358 -395
rect -356 -397 -354 -395
rect -408 -400 -402 -398
rect -408 -402 -406 -400
rect -404 -402 -402 -400
rect -440 -404 -436 -402
rect -440 -407 -438 -404
rect -430 -407 -428 -402
rect -490 -419 -488 -415
rect -517 -425 -515 -420
rect -510 -425 -508 -420
rect -500 -423 -498 -420
rect -479 -423 -477 -412
rect -500 -425 -477 -423
rect -408 -404 -402 -402
rect -408 -407 -406 -404
rect -385 -407 -383 -398
rect -378 -407 -376 -398
rect -360 -399 -354 -397
rect -358 -402 -356 -399
rect -347 -401 -345 -387
rect -337 -389 -335 -387
rect -333 -389 -331 -387
rect -261 -386 -259 -384
rect -257 -386 -255 -384
rect -210 -359 -208 -355
rect -230 -368 -228 -364
rect -220 -368 -218 -364
rect -261 -388 -255 -386
rect -337 -391 -331 -389
rect -257 -389 -255 -388
rect -246 -389 -244 -386
rect -230 -389 -228 -386
rect -257 -391 -244 -389
rect -238 -391 -228 -389
rect -220 -390 -218 -386
rect -210 -389 -208 -386
rect -254 -399 -252 -391
rect -238 -395 -236 -391
rect -245 -397 -236 -395
rect -224 -392 -218 -390
rect -224 -394 -222 -392
rect -220 -394 -218 -392
rect -224 -396 -218 -394
rect -214 -391 -208 -389
rect -214 -393 -212 -391
rect -210 -393 -208 -391
rect -214 -395 -208 -393
rect -245 -399 -243 -397
rect -241 -399 -236 -397
rect -368 -407 -366 -402
rect -420 -419 -418 -415
rect -447 -425 -445 -420
rect -440 -425 -438 -420
rect -430 -423 -428 -420
rect -408 -423 -406 -418
rect -430 -425 -406 -423
rect -245 -401 -236 -399
rect -220 -399 -218 -396
rect -238 -404 -236 -401
rect -228 -404 -226 -400
rect -220 -401 -216 -399
rect -218 -404 -216 -401
rect -211 -404 -209 -395
rect -254 -411 -252 -408
rect -358 -419 -356 -415
rect -385 -425 -383 -420
rect -378 -425 -376 -420
rect -368 -423 -366 -420
rect -347 -423 -345 -412
rect -254 -413 -249 -411
rect -368 -425 -345 -423
rect -251 -421 -249 -413
rect -238 -417 -236 -413
rect -228 -421 -226 -413
rect -218 -421 -216 -416
rect -211 -421 -209 -416
rect -251 -423 -226 -421
rect -762 -430 -737 -428
rect -779 -435 -777 -430
rect -772 -435 -770 -430
rect -762 -438 -760 -430
rect -752 -438 -750 -434
rect -739 -438 -737 -430
rect -739 -440 -734 -438
rect -736 -443 -734 -440
rect -712 -443 -710 -438
rect -684 -439 -682 -434
rect -665 -432 -643 -430
rect -779 -456 -777 -447
rect -772 -450 -770 -447
rect -772 -452 -768 -450
rect -762 -451 -760 -447
rect -752 -450 -750 -447
rect -770 -455 -768 -452
rect -752 -452 -743 -450
rect -672 -441 -670 -436
rect -665 -441 -663 -432
rect -655 -441 -653 -436
rect -645 -441 -643 -432
rect -552 -439 -550 -434
rect -533 -432 -511 -430
rect -752 -454 -747 -452
rect -745 -454 -743 -452
rect -780 -458 -774 -456
rect -780 -460 -778 -458
rect -776 -460 -774 -458
rect -780 -462 -774 -460
rect -770 -457 -764 -455
rect -770 -459 -768 -457
rect -766 -459 -764 -457
rect -770 -461 -764 -459
rect -752 -456 -743 -454
rect -752 -460 -750 -456
rect -736 -460 -734 -452
rect -712 -455 -710 -452
rect -712 -457 -706 -455
rect -712 -459 -710 -457
rect -708 -459 -706 -457
rect -780 -465 -778 -462
rect -770 -465 -768 -461
rect -760 -462 -750 -460
rect -744 -462 -731 -460
rect -760 -465 -758 -462
rect -744 -465 -742 -462
rect -733 -463 -731 -462
rect -712 -461 -706 -459
rect -684 -456 -682 -451
rect -580 -444 -578 -439
rect -540 -441 -538 -436
rect -533 -441 -531 -432
rect -523 -441 -521 -436
rect -513 -441 -511 -432
rect -423 -438 -421 -433
rect -404 -431 -382 -429
rect -672 -456 -670 -453
rect -665 -456 -663 -453
rect -655 -456 -653 -453
rect -645 -456 -643 -453
rect -580 -456 -578 -453
rect -552 -456 -550 -451
rect -448 -443 -446 -438
rect -411 -440 -409 -435
rect -404 -440 -402 -431
rect -394 -440 -392 -435
rect -384 -440 -382 -431
rect -254 -439 -252 -435
rect -241 -437 -239 -432
rect -234 -437 -232 -432
rect -540 -456 -538 -453
rect -533 -456 -531 -453
rect -523 -456 -521 -453
rect -513 -456 -511 -453
rect -448 -455 -446 -452
rect -423 -455 -421 -450
rect -411 -455 -409 -452
rect -404 -455 -402 -452
rect -394 -455 -392 -452
rect -384 -455 -382 -452
rect -254 -453 -252 -448
rect -241 -453 -239 -448
rect -254 -455 -248 -453
rect -684 -458 -669 -456
rect -684 -460 -682 -458
rect -680 -460 -669 -458
rect -665 -459 -662 -456
rect -733 -465 -727 -463
rect -712 -464 -710 -461
rect -684 -462 -669 -460
rect -770 -487 -768 -483
rect -760 -487 -758 -483
rect -780 -496 -778 -492
rect -733 -467 -731 -465
rect -729 -467 -727 -465
rect -733 -469 -727 -467
rect -681 -465 -679 -462
rect -671 -465 -669 -462
rect -664 -465 -662 -459
rect -658 -458 -652 -456
rect -658 -460 -656 -458
rect -654 -460 -652 -458
rect -658 -462 -652 -460
rect -645 -458 -638 -456
rect -645 -460 -642 -458
rect -640 -460 -638 -458
rect -645 -462 -638 -460
rect -580 -458 -574 -456
rect -580 -460 -578 -458
rect -576 -460 -574 -458
rect -580 -462 -574 -460
rect -552 -458 -537 -456
rect -552 -460 -550 -458
rect -548 -460 -537 -458
rect -533 -459 -530 -456
rect -552 -462 -537 -460
rect -654 -465 -652 -462
rect -644 -465 -642 -462
rect -580 -465 -578 -462
rect -549 -465 -547 -462
rect -539 -465 -537 -462
rect -532 -465 -530 -459
rect -526 -458 -520 -456
rect -526 -460 -524 -458
rect -522 -460 -520 -458
rect -526 -462 -520 -460
rect -513 -458 -506 -456
rect -513 -460 -510 -458
rect -508 -460 -506 -458
rect -513 -462 -506 -460
rect -448 -457 -442 -455
rect -448 -459 -446 -457
rect -444 -459 -442 -457
rect -448 -461 -442 -459
rect -423 -457 -408 -455
rect -423 -459 -421 -457
rect -419 -459 -408 -457
rect -404 -458 -401 -455
rect -423 -461 -408 -459
rect -522 -465 -520 -462
rect -512 -465 -510 -462
rect -448 -464 -446 -461
rect -420 -464 -418 -461
rect -410 -464 -408 -461
rect -403 -464 -401 -458
rect -397 -457 -391 -455
rect -397 -459 -395 -457
rect -393 -459 -391 -457
rect -397 -461 -391 -459
rect -384 -457 -377 -455
rect -384 -459 -381 -457
rect -379 -459 -377 -457
rect -384 -461 -377 -459
rect -254 -457 -252 -455
rect -250 -457 -248 -455
rect -254 -459 -248 -457
rect -244 -455 -238 -453
rect -244 -457 -242 -455
rect -240 -457 -238 -455
rect -244 -459 -238 -457
rect -393 -464 -391 -461
rect -383 -464 -381 -461
rect -254 -463 -252 -459
rect -712 -487 -710 -482
rect -744 -496 -742 -492
rect -580 -488 -578 -483
rect -448 -487 -446 -482
rect -244 -470 -242 -459
rect -234 -461 -232 -448
rect -234 -463 -228 -461
rect -234 -465 -232 -463
rect -230 -465 -228 -463
rect -234 -467 -228 -465
rect -234 -470 -232 -467
rect -254 -485 -252 -481
rect -244 -488 -242 -483
rect -234 -488 -232 -483
rect -681 -497 -679 -492
rect -671 -497 -669 -492
rect -664 -497 -662 -492
rect -654 -497 -652 -492
rect -644 -497 -642 -492
rect -549 -497 -547 -492
rect -539 -497 -537 -492
rect -532 -497 -530 -492
rect -522 -497 -520 -492
rect -512 -497 -510 -492
rect -420 -496 -418 -491
rect -410 -496 -408 -491
rect -403 -496 -401 -491
rect -393 -496 -391 -491
rect -383 -496 -381 -491
<< ndif >>
rect -286 136 -281 142
rect -288 134 -281 136
rect -288 132 -286 134
rect -284 132 -281 134
rect -288 130 -281 132
rect -279 130 -274 142
rect -272 140 -260 142
rect -213 144 -206 146
rect -213 142 -211 144
rect -209 142 -206 144
rect -272 138 -264 140
rect -262 138 -260 140
rect -272 130 -260 138
rect -213 136 -206 142
rect -118 144 -111 146
rect -118 142 -116 144
rect -114 142 -111 144
rect -213 134 -204 136
rect -224 132 -217 134
rect -250 129 -245 132
rect -252 127 -245 129
rect -252 125 -250 127
rect -248 125 -245 127
rect -252 123 -245 125
rect -243 130 -232 132
rect -243 128 -236 130
rect -234 128 -232 130
rect -224 130 -222 132
rect -220 130 -217 132
rect -224 128 -217 130
rect -243 123 -232 128
rect -222 125 -217 128
rect -215 125 -204 134
rect -202 125 -197 136
rect -195 134 -188 136
rect -118 136 -111 142
rect -74 143 -67 145
rect -74 141 -72 143
rect -70 141 -67 143
rect -118 134 -109 136
rect -195 132 -192 134
rect -190 132 -188 134
rect -195 130 -188 132
rect -129 132 -122 134
rect -129 130 -127 132
rect -125 130 -122 132
rect -195 125 -190 130
rect -129 128 -122 130
rect -127 125 -122 128
rect -120 125 -109 134
rect -107 125 -102 136
rect -100 134 -93 136
rect -100 132 -97 134
rect -95 132 -93 134
rect -74 135 -67 141
rect -30 144 -23 146
rect -30 142 -28 144
rect -26 142 -23 144
rect -74 133 -65 135
rect -100 130 -93 132
rect -85 131 -78 133
rect -100 125 -95 130
rect -85 129 -83 131
rect -81 129 -78 131
rect -85 127 -78 129
rect -83 124 -78 127
rect -76 124 -65 133
rect -63 124 -58 135
rect -56 133 -49 135
rect -30 136 -23 142
rect 23 144 30 146
rect 23 142 25 144
rect 27 142 30 144
rect -30 134 -21 136
rect -56 131 -53 133
rect -51 131 -49 133
rect -56 129 -49 131
rect -41 132 -34 134
rect -41 130 -39 132
rect -37 130 -34 132
rect -56 124 -51 129
rect -41 128 -34 130
rect -39 125 -34 128
rect -32 125 -21 134
rect -19 125 -14 136
rect -12 134 -5 136
rect 23 136 30 142
rect 67 144 74 146
rect 67 142 69 144
rect 71 142 74 144
rect 23 134 32 136
rect -12 132 -9 134
rect -7 132 -5 134
rect -12 130 -5 132
rect 12 132 19 134
rect 12 130 14 132
rect 16 130 19 132
rect -12 125 -7 130
rect 12 128 19 130
rect 14 125 19 128
rect 21 125 32 134
rect 34 125 39 136
rect 41 134 48 136
rect 67 136 74 142
rect 110 144 117 146
rect 110 142 112 144
rect 114 142 117 144
rect 67 134 76 136
rect 41 132 44 134
rect 46 132 48 134
rect 41 130 48 132
rect 56 132 63 134
rect 56 130 58 132
rect 60 130 63 132
rect 41 125 46 130
rect 56 128 63 130
rect 58 125 63 128
rect 65 125 76 134
rect 78 125 83 136
rect 85 134 92 136
rect 110 136 117 142
rect 110 134 119 136
rect 85 132 88 134
rect 90 132 92 134
rect 85 130 92 132
rect 99 132 106 134
rect 99 130 101 132
rect 103 130 106 132
rect 85 125 90 130
rect 99 128 106 130
rect 101 125 106 128
rect 108 125 119 134
rect 121 125 126 136
rect 128 134 135 136
rect 128 132 131 134
rect 133 132 135 134
rect 128 130 135 132
rect 128 125 133 130
rect -358 25 -353 30
rect -388 12 -380 25
rect -378 12 -373 25
rect -371 22 -363 25
rect -371 20 -368 22
rect -366 20 -363 22
rect -371 12 -363 20
rect -361 23 -353 25
rect -361 21 -358 23
rect -356 21 -353 23
rect -361 17 -353 21
rect -351 25 -343 30
rect -285 30 -280 31
rect -296 25 -291 30
rect -351 17 -341 25
rect -361 12 -356 17
rect -349 15 -341 17
rect -349 13 -347 15
rect -345 14 -341 15
rect -339 23 -332 25
rect -339 21 -336 23
rect -334 21 -332 23
rect -339 19 -332 21
rect -339 14 -334 19
rect -345 13 -343 14
rect -388 10 -386 12
rect -384 10 -382 12
rect -388 8 -382 10
rect -349 11 -343 13
rect -326 12 -318 25
rect -316 12 -311 25
rect -309 22 -301 25
rect -309 20 -306 22
rect -304 20 -301 22
rect -309 12 -301 20
rect -299 23 -291 25
rect -299 21 -296 23
rect -294 21 -291 23
rect -299 17 -291 21
rect -289 21 -280 30
rect -289 19 -286 21
rect -284 20 -280 21
rect -278 29 -271 31
rect -278 27 -275 29
rect -273 27 -271 29
rect -278 25 -271 27
rect -227 25 -222 30
rect -278 20 -273 25
rect -284 19 -282 20
rect -289 17 -282 19
rect -299 12 -294 17
rect -326 10 -324 12
rect -322 10 -320 12
rect -326 8 -320 10
rect -257 12 -249 25
rect -247 12 -242 25
rect -240 22 -232 25
rect -240 20 -237 22
rect -235 20 -232 22
rect -240 12 -232 20
rect -230 23 -222 25
rect -230 21 -227 23
rect -225 21 -222 23
rect -230 17 -222 21
rect -220 25 -212 30
rect -154 30 -149 31
rect -165 25 -160 30
rect -220 17 -210 25
rect -230 12 -225 17
rect -218 15 -210 17
rect -218 13 -216 15
rect -214 14 -210 15
rect -208 23 -201 25
rect -208 21 -205 23
rect -203 21 -201 23
rect -208 19 -201 21
rect -208 14 -203 19
rect -214 13 -212 14
rect -257 10 -255 12
rect -253 10 -251 12
rect -257 8 -251 10
rect -218 11 -212 13
rect -195 12 -187 25
rect -185 12 -180 25
rect -178 22 -170 25
rect -178 20 -175 22
rect -173 20 -170 22
rect -178 12 -170 20
rect -168 23 -160 25
rect -168 21 -165 23
rect -163 21 -160 23
rect -168 17 -160 21
rect -158 21 -149 30
rect -158 19 -155 21
rect -153 20 -149 21
rect -147 29 -140 31
rect -147 27 -144 29
rect -142 27 -140 29
rect -147 25 -140 27
rect -95 25 -90 30
rect -147 20 -142 25
rect -153 19 -151 20
rect -158 17 -151 19
rect -168 12 -163 17
rect -195 10 -193 12
rect -191 10 -189 12
rect -195 8 -189 10
rect -125 12 -117 25
rect -115 12 -110 25
rect -108 22 -100 25
rect -108 20 -105 22
rect -103 20 -100 22
rect -108 12 -100 20
rect -98 23 -90 25
rect -98 21 -95 23
rect -93 21 -90 23
rect -98 17 -90 21
rect -88 25 -80 30
rect -22 30 -17 31
rect -33 25 -28 30
rect -88 17 -78 25
rect -98 12 -93 17
rect -86 15 -78 17
rect -86 13 -84 15
rect -82 14 -78 15
rect -76 23 -69 25
rect -76 21 -73 23
rect -71 21 -69 23
rect -76 19 -69 21
rect -76 14 -71 19
rect -82 13 -80 14
rect -125 10 -123 12
rect -121 10 -119 12
rect -125 8 -119 10
rect -86 11 -80 13
rect -63 12 -55 25
rect -53 12 -48 25
rect -46 22 -38 25
rect -46 20 -43 22
rect -41 20 -38 22
rect -46 12 -38 20
rect -36 23 -28 25
rect -36 21 -33 23
rect -31 21 -28 23
rect -36 17 -28 21
rect -26 21 -17 30
rect -26 19 -23 21
rect -21 20 -17 21
rect -15 29 -8 31
rect -15 27 -12 29
rect -10 27 -8 29
rect -15 25 -8 27
rect 7 29 14 31
rect 7 27 9 29
rect 11 27 14 29
rect 7 25 14 27
rect -15 20 -10 25
rect 9 22 14 25
rect 16 26 21 31
rect 16 22 30 26
rect -21 19 -19 20
rect -26 17 -19 19
rect -36 12 -31 17
rect -63 10 -61 12
rect -59 10 -57 12
rect -63 8 -57 10
rect 21 21 30 22
rect 21 19 23 21
rect 25 19 30 21
rect 21 17 30 19
rect 32 24 40 26
rect 32 22 35 24
rect 37 22 40 24
rect 32 17 40 22
rect 42 22 50 26
rect 42 20 45 22
rect 47 20 50 22
rect 42 17 50 20
rect 45 14 50 17
rect 52 14 57 26
rect 59 14 67 26
rect 61 12 67 14
rect 61 10 63 12
rect 65 10 67 12
rect 61 8 67 10
rect -341 1 -335 3
rect -341 -1 -339 1
rect -337 -1 -335 1
rect -341 -6 -335 -1
rect -352 -8 -345 -6
rect -352 -10 -350 -8
rect -348 -10 -345 -8
rect -376 -14 -371 -11
rect -378 -16 -371 -14
rect -378 -18 -376 -16
rect -374 -18 -371 -16
rect -378 -20 -371 -18
rect -369 -13 -358 -11
rect -352 -12 -345 -10
rect -369 -15 -362 -13
rect -360 -15 -358 -13
rect -369 -20 -358 -15
rect -350 -18 -345 -12
rect -343 -8 -335 -6
rect -245 1 -239 3
rect -245 -1 -243 1
rect -241 -1 -239 1
rect -245 -6 -239 -1
rect -343 -18 -333 -8
rect -341 -20 -333 -18
rect -331 -20 -326 -8
rect -324 -16 -316 -8
rect -324 -18 -321 -16
rect -319 -18 -316 -16
rect -324 -20 -316 -18
rect -314 -10 -306 -8
rect -314 -12 -311 -10
rect -309 -12 -306 -10
rect -314 -20 -306 -12
rect -304 -10 -296 -8
rect -304 -12 -301 -10
rect -299 -12 -296 -10
rect -256 -8 -249 -6
rect -256 -10 -254 -8
rect -252 -10 -249 -8
rect -304 -20 -296 -12
rect -282 -14 -277 -11
rect -284 -16 -277 -14
rect -284 -18 -282 -16
rect -280 -18 -277 -16
rect -284 -20 -277 -18
rect -275 -13 -264 -11
rect -256 -12 -249 -10
rect -275 -15 -268 -13
rect -266 -15 -264 -13
rect -275 -20 -264 -15
rect -254 -18 -249 -12
rect -247 -8 -239 -6
rect -113 0 -107 2
rect -113 -2 -111 0
rect -109 -2 -107 0
rect -113 -7 -107 -2
rect -247 -18 -237 -8
rect -245 -20 -237 -18
rect -235 -20 -230 -8
rect -228 -16 -220 -8
rect -228 -18 -225 -16
rect -223 -18 -220 -16
rect -228 -20 -220 -18
rect -218 -10 -210 -8
rect -218 -12 -215 -10
rect -213 -12 -210 -10
rect -218 -20 -210 -12
rect -208 -10 -200 -8
rect -208 -12 -205 -10
rect -203 -12 -200 -10
rect -124 -9 -117 -7
rect -124 -11 -122 -9
rect -120 -11 -117 -9
rect -208 -20 -200 -12
rect -149 -15 -144 -12
rect -151 -17 -144 -15
rect -151 -19 -149 -17
rect -147 -19 -144 -17
rect -151 -21 -144 -19
rect -142 -14 -131 -12
rect -124 -13 -117 -11
rect -142 -16 -135 -14
rect -133 -16 -131 -14
rect -142 -21 -131 -16
rect -122 -19 -117 -13
rect -115 -9 -107 -7
rect 20 0 27 2
rect 20 -2 22 0
rect 24 -2 27 0
rect -115 -19 -105 -9
rect -113 -21 -105 -19
rect -103 -21 -98 -9
rect -96 -17 -88 -9
rect -96 -19 -93 -17
rect -91 -19 -88 -17
rect -96 -21 -88 -19
rect -86 -11 -78 -9
rect -86 -13 -83 -11
rect -81 -13 -78 -11
rect -86 -21 -78 -13
rect -76 -11 -68 -9
rect 20 -8 27 -2
rect 20 -10 29 -8
rect -76 -13 -73 -11
rect -71 -13 -68 -11
rect -76 -21 -68 -13
rect 9 -12 16 -10
rect 9 -14 11 -12
rect 13 -14 16 -12
rect 9 -16 16 -14
rect 11 -19 16 -16
rect 18 -19 29 -10
rect 31 -19 36 -8
rect 38 -10 45 -8
rect 38 -12 41 -10
rect 43 -12 45 -10
rect 38 -14 45 -12
rect 38 -19 43 -14
rect -450 -116 -443 -114
rect -450 -118 -448 -116
rect -446 -118 -443 -116
rect -450 -120 -443 -118
rect -448 -123 -443 -120
rect -441 -119 -430 -114
rect -420 -118 -415 -115
rect -441 -121 -434 -119
rect -432 -121 -430 -119
rect -441 -123 -430 -121
rect -422 -120 -415 -118
rect -422 -122 -420 -120
rect -418 -122 -415 -120
rect -422 -124 -415 -122
rect -413 -124 -402 -115
rect -411 -126 -402 -124
rect -400 -126 -395 -115
rect -393 -120 -388 -115
rect -308 -117 -303 -114
rect -310 -119 -303 -117
rect -393 -122 -386 -120
rect -393 -124 -390 -122
rect -388 -124 -386 -122
rect -310 -121 -308 -119
rect -306 -121 -303 -119
rect -310 -123 -303 -121
rect -301 -123 -290 -114
rect -393 -126 -386 -124
rect -411 -132 -404 -126
rect -299 -125 -290 -123
rect -288 -125 -283 -114
rect -281 -119 -276 -114
rect -157 -118 -152 -115
rect -281 -121 -274 -119
rect -281 -123 -278 -121
rect -276 -123 -274 -121
rect -281 -125 -274 -123
rect -159 -120 -152 -118
rect -159 -122 -157 -120
rect -155 -122 -152 -120
rect -159 -124 -152 -122
rect -150 -124 -139 -115
rect -411 -134 -409 -132
rect -407 -134 -404 -132
rect -411 -136 -404 -134
rect -299 -131 -292 -125
rect -148 -126 -139 -124
rect -137 -126 -132 -115
rect -130 -120 -125 -115
rect -113 -118 -108 -115
rect -115 -120 -108 -118
rect -130 -122 -123 -120
rect -130 -124 -127 -122
rect -125 -124 -123 -122
rect -115 -122 -113 -120
rect -111 -122 -108 -120
rect -115 -124 -108 -122
rect -106 -124 -95 -115
rect -130 -126 -123 -124
rect -299 -133 -297 -131
rect -295 -133 -292 -131
rect -299 -135 -292 -133
rect -148 -132 -141 -126
rect -104 -126 -95 -124
rect -93 -126 -88 -115
rect -86 -120 -81 -115
rect -86 -122 -79 -120
rect -86 -124 -83 -122
rect -81 -124 -79 -122
rect -86 -126 -79 -124
rect -148 -134 -146 -132
rect -144 -134 -141 -132
rect -148 -136 -141 -134
rect -104 -132 -97 -126
rect -104 -134 -102 -132
rect -100 -134 -97 -132
rect -104 -136 -97 -134
rect -541 -145 -535 -143
rect -541 -147 -539 -145
rect -537 -147 -535 -145
rect -541 -160 -533 -147
rect -531 -160 -526 -147
rect -524 -155 -516 -147
rect -524 -157 -521 -155
rect -519 -157 -516 -155
rect -524 -160 -516 -157
rect -514 -152 -509 -147
rect -502 -148 -496 -146
rect -502 -150 -500 -148
rect -498 -149 -496 -148
rect -479 -145 -473 -143
rect -479 -147 -477 -145
rect -475 -147 -473 -145
rect -498 -150 -494 -149
rect -502 -152 -494 -150
rect -514 -156 -506 -152
rect -514 -158 -511 -156
rect -509 -158 -506 -156
rect -514 -160 -506 -158
rect -511 -165 -506 -160
rect -504 -160 -494 -152
rect -492 -154 -487 -149
rect -492 -156 -485 -154
rect -492 -158 -489 -156
rect -487 -158 -485 -156
rect -492 -160 -485 -158
rect -479 -160 -471 -147
rect -469 -160 -464 -147
rect -462 -155 -454 -147
rect -462 -157 -459 -155
rect -457 -157 -454 -155
rect -462 -160 -454 -157
rect -452 -152 -447 -147
rect -452 -156 -444 -152
rect -452 -158 -449 -156
rect -447 -158 -444 -156
rect -452 -160 -444 -158
rect -504 -165 -496 -160
rect -449 -165 -444 -160
rect -442 -154 -435 -152
rect -442 -156 -439 -154
rect -437 -155 -435 -154
rect -409 -145 -403 -143
rect -409 -147 -407 -145
rect -405 -147 -403 -145
rect -437 -156 -433 -155
rect -442 -165 -433 -156
rect -438 -166 -433 -165
rect -431 -160 -426 -155
rect -409 -160 -401 -147
rect -399 -160 -394 -147
rect -392 -155 -384 -147
rect -392 -157 -389 -155
rect -387 -157 -384 -155
rect -392 -160 -384 -157
rect -382 -152 -377 -147
rect -370 -148 -364 -146
rect -370 -150 -368 -148
rect -366 -149 -364 -148
rect -347 -145 -341 -143
rect -347 -147 -345 -145
rect -343 -147 -341 -145
rect -366 -150 -362 -149
rect -370 -152 -362 -150
rect -382 -156 -374 -152
rect -382 -158 -379 -156
rect -377 -158 -374 -156
rect -382 -160 -374 -158
rect -431 -162 -424 -160
rect -431 -164 -428 -162
rect -426 -164 -424 -162
rect -431 -166 -424 -164
rect -379 -165 -374 -160
rect -372 -160 -362 -152
rect -360 -154 -355 -149
rect -360 -156 -353 -154
rect -360 -158 -357 -156
rect -355 -158 -353 -156
rect -360 -160 -353 -158
rect -347 -160 -339 -147
rect -337 -160 -332 -147
rect -330 -155 -322 -147
rect -330 -157 -327 -155
rect -325 -157 -322 -155
rect -330 -160 -322 -157
rect -320 -152 -315 -147
rect -320 -156 -312 -152
rect -320 -158 -317 -156
rect -315 -158 -312 -156
rect -320 -160 -312 -158
rect -372 -165 -364 -160
rect -317 -165 -312 -160
rect -310 -154 -303 -152
rect -310 -156 -307 -154
rect -305 -155 -303 -154
rect -272 -144 -266 -142
rect -272 -146 -270 -144
rect -268 -146 -266 -144
rect -305 -156 -301 -155
rect -310 -165 -301 -156
rect -306 -166 -301 -165
rect -299 -160 -294 -155
rect -272 -159 -264 -146
rect -262 -159 -257 -146
rect -255 -154 -247 -146
rect -255 -156 -252 -154
rect -250 -156 -247 -154
rect -255 -159 -247 -156
rect -245 -151 -240 -146
rect -233 -147 -227 -145
rect -233 -149 -231 -147
rect -229 -148 -227 -147
rect -210 -144 -204 -142
rect -210 -146 -208 -144
rect -206 -146 -204 -144
rect -229 -149 -225 -148
rect -233 -151 -225 -149
rect -245 -155 -237 -151
rect -245 -157 -242 -155
rect -240 -157 -237 -155
rect -245 -159 -237 -157
rect -299 -162 -292 -160
rect -299 -164 -296 -162
rect -294 -164 -292 -162
rect -299 -166 -292 -164
rect -242 -164 -237 -159
rect -235 -159 -225 -151
rect -223 -153 -218 -148
rect -223 -155 -216 -153
rect -223 -157 -220 -155
rect -218 -157 -216 -155
rect -223 -159 -216 -157
rect -210 -159 -202 -146
rect -200 -159 -195 -146
rect -193 -154 -185 -146
rect -193 -156 -190 -154
rect -188 -156 -185 -154
rect -193 -159 -185 -156
rect -183 -151 -178 -146
rect -183 -155 -175 -151
rect -183 -157 -180 -155
rect -178 -157 -175 -155
rect -183 -159 -175 -157
rect -235 -164 -227 -159
rect -180 -164 -175 -159
rect -173 -153 -166 -151
rect -173 -155 -170 -153
rect -168 -154 -166 -153
rect -141 -144 -135 -142
rect -141 -146 -139 -144
rect -137 -146 -135 -144
rect -141 -148 -135 -146
rect -168 -155 -164 -154
rect -173 -164 -164 -155
rect -169 -165 -164 -164
rect -162 -159 -157 -154
rect -162 -161 -155 -159
rect -141 -160 -133 -148
rect -131 -160 -126 -148
rect -124 -151 -119 -148
rect -124 -154 -116 -151
rect -124 -156 -121 -154
rect -119 -156 -116 -154
rect -124 -160 -116 -156
rect -114 -156 -106 -151
rect -114 -158 -111 -156
rect -109 -158 -106 -156
rect -114 -160 -106 -158
rect -104 -153 -95 -151
rect -104 -155 -99 -153
rect -97 -155 -95 -153
rect -104 -156 -95 -155
rect -104 -160 -90 -156
rect -162 -163 -159 -161
rect -157 -163 -155 -161
rect -162 -165 -155 -163
rect -95 -165 -90 -160
rect -88 -159 -83 -156
rect -88 -161 -81 -159
rect -88 -163 -85 -161
rect -83 -163 -81 -161
rect -88 -165 -81 -163
rect -502 -260 -495 -258
rect -502 -262 -500 -260
rect -498 -262 -495 -260
rect -502 -264 -495 -262
rect -500 -267 -495 -264
rect -493 -263 -482 -258
rect -465 -260 -457 -258
rect -493 -265 -486 -263
rect -484 -265 -482 -263
rect -493 -267 -482 -265
rect -474 -266 -469 -260
rect -476 -268 -469 -266
rect -476 -270 -474 -268
rect -472 -270 -469 -268
rect -476 -272 -469 -270
rect -467 -270 -457 -260
rect -455 -270 -450 -258
rect -448 -260 -440 -258
rect -448 -262 -445 -260
rect -443 -262 -440 -260
rect -448 -270 -440 -262
rect -438 -266 -430 -258
rect -438 -268 -435 -266
rect -433 -268 -430 -266
rect -438 -270 -430 -268
rect -428 -266 -420 -258
rect -409 -260 -402 -258
rect -409 -262 -407 -260
rect -405 -262 -402 -260
rect -409 -264 -402 -262
rect -428 -268 -425 -266
rect -423 -268 -420 -266
rect -407 -267 -402 -264
rect -400 -263 -389 -258
rect -371 -260 -363 -258
rect -400 -265 -393 -263
rect -391 -265 -389 -263
rect -400 -267 -389 -265
rect -380 -266 -375 -260
rect -428 -270 -420 -268
rect -467 -272 -459 -270
rect -465 -277 -459 -272
rect -465 -279 -463 -277
rect -461 -279 -459 -277
rect -465 -281 -459 -279
rect -382 -268 -375 -266
rect -382 -270 -380 -268
rect -378 -270 -375 -268
rect -382 -272 -375 -270
rect -373 -270 -363 -260
rect -361 -270 -356 -258
rect -354 -260 -346 -258
rect -354 -262 -351 -260
rect -349 -262 -346 -260
rect -354 -270 -346 -262
rect -344 -266 -336 -258
rect -344 -268 -341 -266
rect -339 -268 -336 -266
rect -344 -270 -336 -268
rect -334 -266 -326 -258
rect -236 -259 -229 -257
rect -236 -261 -234 -259
rect -232 -261 -229 -259
rect -236 -263 -229 -261
rect -234 -266 -229 -263
rect -227 -262 -216 -257
rect -197 -259 -189 -257
rect -227 -264 -220 -262
rect -218 -264 -216 -262
rect -227 -266 -216 -264
rect -206 -265 -201 -259
rect -334 -268 -331 -266
rect -329 -268 -326 -266
rect -334 -270 -326 -268
rect -373 -272 -365 -270
rect -371 -277 -365 -272
rect -371 -279 -369 -277
rect -367 -279 -365 -277
rect -371 -281 -365 -279
rect -208 -267 -201 -265
rect -208 -269 -206 -267
rect -204 -269 -201 -267
rect -208 -271 -201 -269
rect -199 -269 -189 -259
rect -187 -269 -182 -257
rect -180 -259 -172 -257
rect -180 -261 -177 -259
rect -175 -261 -172 -259
rect -180 -269 -172 -261
rect -170 -265 -162 -257
rect -170 -267 -167 -265
rect -165 -267 -162 -265
rect -170 -269 -162 -267
rect -160 -265 -152 -257
rect -139 -262 -134 -259
rect -160 -267 -157 -265
rect -155 -267 -152 -265
rect -160 -269 -152 -267
rect -141 -264 -134 -262
rect -141 -266 -139 -264
rect -137 -266 -134 -264
rect -141 -268 -134 -266
rect -132 -268 -121 -259
rect -199 -271 -191 -269
rect -197 -276 -191 -271
rect -197 -278 -195 -276
rect -193 -278 -191 -276
rect -197 -280 -191 -278
rect -130 -270 -121 -268
rect -119 -270 -114 -259
rect -112 -264 -107 -259
rect -112 -266 -105 -264
rect -112 -268 -109 -266
rect -107 -268 -105 -266
rect -112 -270 -105 -268
rect -130 -276 -123 -270
rect -130 -278 -128 -276
rect -126 -278 -123 -276
rect -130 -280 -123 -278
rect -567 -289 -560 -287
rect -567 -291 -565 -289
rect -563 -291 -560 -289
rect -567 -297 -560 -291
rect -503 -297 -498 -291
rect -567 -299 -558 -297
rect -578 -301 -571 -299
rect -578 -303 -576 -301
rect -574 -303 -571 -301
rect -578 -305 -571 -303
rect -576 -308 -571 -305
rect -569 -308 -558 -299
rect -556 -308 -551 -297
rect -549 -299 -542 -297
rect -549 -301 -546 -299
rect -544 -301 -542 -299
rect -549 -303 -542 -301
rect -505 -299 -498 -297
rect -505 -301 -503 -299
rect -501 -301 -498 -299
rect -505 -303 -498 -301
rect -496 -303 -491 -291
rect -489 -293 -477 -291
rect -489 -295 -481 -293
rect -479 -295 -477 -293
rect -489 -303 -477 -295
rect -379 -297 -374 -291
rect -381 -299 -374 -297
rect -381 -301 -379 -299
rect -377 -301 -374 -299
rect -381 -303 -374 -301
rect -372 -303 -367 -291
rect -365 -293 -353 -291
rect -365 -295 -357 -293
rect -355 -295 -353 -293
rect -365 -303 -353 -295
rect -233 -296 -228 -290
rect -235 -298 -228 -296
rect -235 -300 -233 -298
rect -231 -300 -228 -298
rect -235 -302 -228 -300
rect -226 -302 -221 -290
rect -219 -292 -207 -290
rect -219 -294 -211 -292
rect -209 -294 -207 -292
rect -219 -302 -207 -294
rect -549 -308 -544 -303
rect -689 -407 -684 -402
rect -719 -420 -711 -407
rect -709 -420 -704 -407
rect -702 -410 -694 -407
rect -702 -412 -699 -410
rect -697 -412 -694 -410
rect -702 -420 -694 -412
rect -692 -409 -684 -407
rect -692 -411 -689 -409
rect -687 -411 -684 -409
rect -692 -415 -684 -411
rect -682 -407 -674 -402
rect -616 -402 -611 -401
rect -627 -407 -622 -402
rect -682 -415 -672 -407
rect -692 -420 -687 -415
rect -680 -417 -672 -415
rect -680 -419 -678 -417
rect -676 -418 -672 -417
rect -670 -409 -663 -407
rect -670 -411 -667 -409
rect -665 -411 -663 -409
rect -670 -413 -663 -411
rect -670 -418 -665 -413
rect -676 -419 -674 -418
rect -719 -422 -717 -420
rect -715 -422 -713 -420
rect -719 -424 -713 -422
rect -680 -421 -674 -419
rect -657 -420 -649 -407
rect -647 -420 -642 -407
rect -640 -410 -632 -407
rect -640 -412 -637 -410
rect -635 -412 -632 -410
rect -640 -420 -632 -412
rect -630 -409 -622 -407
rect -630 -411 -627 -409
rect -625 -411 -622 -409
rect -630 -415 -622 -411
rect -620 -411 -611 -402
rect -620 -413 -617 -411
rect -615 -412 -611 -411
rect -609 -403 -602 -401
rect -609 -405 -606 -403
rect -604 -405 -602 -403
rect -609 -407 -602 -405
rect -557 -407 -552 -402
rect -609 -412 -604 -407
rect -615 -413 -613 -412
rect -620 -415 -613 -413
rect -630 -420 -625 -415
rect -657 -422 -655 -420
rect -653 -422 -651 -420
rect -657 -424 -651 -422
rect -587 -420 -579 -407
rect -577 -420 -572 -407
rect -570 -410 -562 -407
rect -570 -412 -567 -410
rect -565 -412 -562 -410
rect -570 -420 -562 -412
rect -560 -409 -552 -407
rect -560 -411 -557 -409
rect -555 -411 -552 -409
rect -560 -415 -552 -411
rect -550 -407 -542 -402
rect -484 -402 -479 -401
rect -495 -407 -490 -402
rect -550 -415 -540 -407
rect -560 -420 -555 -415
rect -548 -417 -540 -415
rect -548 -419 -546 -417
rect -544 -418 -540 -417
rect -538 -409 -531 -407
rect -538 -411 -535 -409
rect -533 -411 -531 -409
rect -538 -413 -531 -411
rect -538 -418 -533 -413
rect -544 -419 -542 -418
rect -587 -422 -585 -420
rect -583 -422 -581 -420
rect -587 -424 -581 -422
rect -548 -421 -542 -419
rect -525 -420 -517 -407
rect -515 -420 -510 -407
rect -508 -410 -500 -407
rect -508 -412 -505 -410
rect -503 -412 -500 -410
rect -508 -420 -500 -412
rect -498 -409 -490 -407
rect -498 -411 -495 -409
rect -493 -411 -490 -409
rect -498 -415 -490 -411
rect -488 -411 -479 -402
rect -488 -413 -485 -411
rect -483 -412 -479 -411
rect -477 -403 -470 -401
rect -477 -405 -474 -403
rect -472 -405 -470 -403
rect -477 -407 -470 -405
rect -425 -407 -420 -402
rect -477 -412 -472 -407
rect -483 -413 -481 -412
rect -488 -415 -481 -413
rect -498 -420 -493 -415
rect -525 -422 -523 -420
rect -521 -422 -519 -420
rect -525 -424 -519 -422
rect -455 -420 -447 -407
rect -445 -420 -440 -407
rect -438 -410 -430 -407
rect -438 -412 -435 -410
rect -433 -412 -430 -410
rect -438 -420 -430 -412
rect -428 -409 -420 -407
rect -428 -411 -425 -409
rect -423 -411 -420 -409
rect -428 -415 -420 -411
rect -418 -407 -410 -402
rect -261 -401 -254 -399
rect -352 -402 -347 -401
rect -363 -407 -358 -402
rect -418 -415 -408 -407
rect -428 -420 -423 -415
rect -416 -417 -408 -415
rect -416 -419 -414 -417
rect -412 -418 -408 -417
rect -406 -409 -399 -407
rect -406 -411 -403 -409
rect -401 -411 -399 -409
rect -406 -413 -399 -411
rect -406 -418 -401 -413
rect -412 -419 -410 -418
rect -455 -422 -453 -420
rect -451 -422 -449 -420
rect -455 -424 -449 -422
rect -416 -421 -410 -419
rect -393 -420 -385 -407
rect -383 -420 -378 -407
rect -376 -410 -368 -407
rect -376 -412 -373 -410
rect -371 -412 -368 -410
rect -376 -420 -368 -412
rect -366 -409 -358 -407
rect -366 -411 -363 -409
rect -361 -411 -358 -409
rect -366 -415 -358 -411
rect -356 -411 -347 -402
rect -356 -413 -353 -411
rect -351 -412 -347 -411
rect -345 -403 -338 -401
rect -345 -405 -342 -403
rect -340 -405 -338 -403
rect -261 -403 -259 -401
rect -257 -403 -254 -401
rect -261 -405 -254 -403
rect -345 -407 -338 -405
rect -345 -412 -340 -407
rect -259 -408 -254 -405
rect -252 -404 -247 -399
rect -252 -408 -238 -404
rect -247 -409 -238 -408
rect -247 -411 -245 -409
rect -243 -411 -238 -409
rect -351 -413 -349 -412
rect -356 -415 -349 -413
rect -366 -420 -361 -415
rect -393 -422 -391 -420
rect -389 -422 -387 -420
rect -393 -424 -387 -422
rect -247 -413 -238 -411
rect -236 -406 -228 -404
rect -236 -408 -233 -406
rect -231 -408 -228 -406
rect -236 -413 -228 -408
rect -226 -408 -218 -404
rect -226 -410 -223 -408
rect -221 -410 -218 -408
rect -226 -413 -218 -410
rect -223 -416 -218 -413
rect -216 -416 -211 -404
rect -209 -416 -201 -404
rect -207 -418 -201 -416
rect -207 -420 -205 -418
rect -203 -420 -201 -418
rect -207 -422 -201 -420
rect -787 -431 -781 -429
rect -787 -433 -785 -431
rect -783 -433 -781 -431
rect -787 -435 -781 -433
rect -787 -447 -779 -435
rect -777 -447 -772 -435
rect -770 -438 -765 -435
rect -680 -432 -674 -430
rect -680 -434 -678 -432
rect -676 -434 -674 -432
rect -770 -441 -762 -438
rect -770 -443 -767 -441
rect -765 -443 -762 -441
rect -770 -447 -762 -443
rect -760 -443 -752 -438
rect -760 -445 -757 -443
rect -755 -445 -752 -443
rect -760 -447 -752 -445
rect -750 -443 -741 -438
rect -680 -439 -674 -434
rect -691 -441 -684 -439
rect -691 -443 -689 -441
rect -687 -443 -684 -441
rect -750 -447 -736 -443
rect -741 -452 -736 -447
rect -734 -446 -729 -443
rect -717 -446 -712 -443
rect -734 -448 -727 -446
rect -734 -450 -731 -448
rect -729 -450 -727 -448
rect -734 -452 -727 -450
rect -719 -448 -712 -446
rect -719 -450 -717 -448
rect -715 -450 -712 -448
rect -719 -452 -712 -450
rect -710 -445 -699 -443
rect -691 -445 -684 -443
rect -710 -447 -703 -445
rect -701 -447 -699 -445
rect -710 -452 -699 -447
rect -689 -451 -684 -445
rect -682 -441 -674 -439
rect -548 -432 -542 -430
rect -548 -434 -546 -432
rect -544 -434 -542 -432
rect -548 -439 -542 -434
rect -682 -451 -672 -441
rect -680 -453 -672 -451
rect -670 -453 -665 -441
rect -663 -449 -655 -441
rect -663 -451 -660 -449
rect -658 -451 -655 -449
rect -663 -453 -655 -451
rect -653 -443 -645 -441
rect -653 -445 -650 -443
rect -648 -445 -645 -443
rect -653 -453 -645 -445
rect -643 -443 -635 -441
rect -643 -445 -640 -443
rect -638 -445 -635 -443
rect -559 -441 -552 -439
rect -559 -443 -557 -441
rect -555 -443 -552 -441
rect -643 -453 -635 -445
rect -585 -447 -580 -444
rect -587 -449 -580 -447
rect -587 -451 -585 -449
rect -583 -451 -580 -449
rect -587 -453 -580 -451
rect -578 -446 -567 -444
rect -559 -445 -552 -443
rect -578 -448 -571 -446
rect -569 -448 -567 -446
rect -578 -453 -567 -448
rect -557 -451 -552 -445
rect -550 -441 -542 -439
rect -419 -431 -413 -429
rect -419 -433 -417 -431
rect -415 -433 -413 -431
rect -419 -438 -413 -433
rect -550 -451 -540 -441
rect -548 -453 -540 -451
rect -538 -453 -533 -441
rect -531 -449 -523 -441
rect -531 -451 -528 -449
rect -526 -451 -523 -449
rect -531 -453 -523 -451
rect -521 -443 -513 -441
rect -521 -445 -518 -443
rect -516 -445 -513 -443
rect -521 -453 -513 -445
rect -511 -443 -503 -441
rect -430 -440 -423 -438
rect -430 -442 -428 -440
rect -426 -442 -423 -440
rect -511 -445 -508 -443
rect -506 -445 -503 -443
rect -511 -453 -503 -445
rect -453 -446 -448 -443
rect -455 -448 -448 -446
rect -455 -450 -453 -448
rect -451 -450 -448 -448
rect -455 -452 -448 -450
rect -446 -445 -435 -443
rect -430 -444 -423 -442
rect -446 -447 -439 -445
rect -437 -447 -435 -445
rect -446 -452 -435 -447
rect -428 -450 -423 -444
rect -421 -440 -413 -438
rect -250 -429 -243 -427
rect -250 -431 -248 -429
rect -246 -431 -243 -429
rect -250 -437 -243 -431
rect -250 -439 -241 -437
rect -421 -450 -411 -440
rect -419 -452 -411 -450
rect -409 -452 -404 -440
rect -402 -448 -394 -440
rect -402 -450 -399 -448
rect -397 -450 -394 -448
rect -402 -452 -394 -450
rect -392 -442 -384 -440
rect -392 -444 -389 -442
rect -387 -444 -384 -442
rect -392 -452 -384 -444
rect -382 -442 -374 -440
rect -382 -444 -379 -442
rect -377 -444 -374 -442
rect -382 -452 -374 -444
rect -261 -441 -254 -439
rect -261 -443 -259 -441
rect -257 -443 -254 -441
rect -261 -445 -254 -443
rect -259 -448 -254 -445
rect -252 -448 -241 -439
rect -239 -448 -234 -437
rect -232 -439 -225 -437
rect -232 -441 -229 -439
rect -227 -441 -225 -439
rect -232 -443 -225 -441
rect -232 -448 -227 -443
<< pdif >>
rect -252 109 -245 111
rect -252 107 -250 109
rect -248 107 -245 109
rect -288 94 -280 106
rect -288 92 -286 94
rect -284 92 -280 94
rect -278 103 -270 106
rect -278 101 -275 103
rect -273 101 -270 103
rect -278 96 -270 101
rect -278 94 -275 96
rect -273 94 -270 96
rect -278 92 -270 94
rect -268 103 -260 106
rect -268 101 -264 103
rect -262 101 -260 103
rect -268 96 -260 101
rect -252 102 -245 107
rect -252 100 -250 102
rect -248 100 -245 102
rect -252 98 -245 100
rect -268 94 -264 96
rect -262 94 -260 96
rect -268 92 -260 94
rect -250 93 -245 98
rect -243 94 -234 111
rect -224 108 -217 110
rect -224 106 -222 108
rect -220 106 -217 108
rect -224 101 -217 106
rect -224 99 -222 101
rect -220 99 -217 101
rect -224 97 -217 99
rect -243 93 -239 94
rect -288 90 -282 92
rect -241 92 -239 93
rect -237 92 -234 94
rect -222 92 -217 97
rect -215 103 -209 110
rect -129 108 -122 110
rect -129 106 -127 108
rect -125 106 -122 108
rect -215 96 -207 103
rect -215 94 -212 96
rect -210 94 -207 96
rect -215 92 -207 94
rect -241 90 -234 92
rect -213 90 -207 92
rect -205 101 -197 103
rect -205 99 -202 101
rect -200 99 -197 101
rect -205 94 -197 99
rect -205 92 -202 94
rect -200 92 -197 94
rect -205 90 -197 92
rect -195 94 -188 103
rect -129 101 -122 106
rect -129 99 -127 101
rect -125 99 -122 101
rect -129 97 -122 99
rect -195 92 -192 94
rect -190 92 -188 94
rect -127 92 -122 97
rect -120 103 -114 110
rect -85 107 -78 109
rect -85 105 -83 107
rect -81 105 -78 107
rect -120 96 -112 103
rect -120 94 -117 96
rect -115 94 -112 96
rect -120 92 -112 94
rect -195 90 -188 92
rect -118 90 -112 92
rect -110 101 -102 103
rect -110 99 -107 101
rect -105 99 -102 101
rect -110 94 -102 99
rect -110 92 -107 94
rect -105 92 -102 94
rect -110 90 -102 92
rect -100 94 -93 103
rect -85 100 -78 105
rect -85 98 -83 100
rect -81 98 -78 100
rect -85 96 -78 98
rect -100 92 -97 94
rect -95 92 -93 94
rect -100 90 -93 92
rect -83 91 -78 96
rect -76 102 -70 109
rect -41 108 -34 110
rect -41 106 -39 108
rect -37 106 -34 108
rect -76 95 -68 102
rect -76 93 -73 95
rect -71 93 -68 95
rect -76 91 -68 93
rect -74 89 -68 91
rect -66 100 -58 102
rect -66 98 -63 100
rect -61 98 -58 100
rect -66 93 -58 98
rect -66 91 -63 93
rect -61 91 -58 93
rect -66 89 -58 91
rect -56 93 -49 102
rect -41 101 -34 106
rect -41 99 -39 101
rect -37 99 -34 101
rect -41 97 -34 99
rect -56 91 -53 93
rect -51 91 -49 93
rect -39 92 -34 97
rect -32 103 -26 110
rect 12 108 19 110
rect 12 106 14 108
rect 16 106 19 108
rect -32 96 -24 103
rect -32 94 -29 96
rect -27 94 -24 96
rect -32 92 -24 94
rect -56 89 -49 91
rect -30 90 -24 92
rect -22 101 -14 103
rect -22 99 -19 101
rect -17 99 -14 101
rect -22 94 -14 99
rect -22 92 -19 94
rect -17 92 -14 94
rect -22 90 -14 92
rect -12 94 -5 103
rect 12 101 19 106
rect 12 99 14 101
rect 16 99 19 101
rect 12 97 19 99
rect -12 92 -9 94
rect -7 92 -5 94
rect 14 92 19 97
rect 21 103 27 110
rect 56 108 63 110
rect 56 106 58 108
rect 60 106 63 108
rect 21 96 29 103
rect 21 94 24 96
rect 26 94 29 96
rect 21 92 29 94
rect -12 90 -5 92
rect 23 90 29 92
rect 31 101 39 103
rect 31 99 34 101
rect 36 99 39 101
rect 31 94 39 99
rect 31 92 34 94
rect 36 92 39 94
rect 31 90 39 92
rect 41 94 48 103
rect 56 101 63 106
rect 56 99 58 101
rect 60 99 63 101
rect 56 97 63 99
rect 41 92 44 94
rect 46 92 48 94
rect 58 92 63 97
rect 65 103 71 110
rect 99 108 106 110
rect 99 106 101 108
rect 103 106 106 108
rect 65 96 73 103
rect 65 94 68 96
rect 70 94 73 96
rect 65 92 73 94
rect 41 90 48 92
rect 67 90 73 92
rect 75 101 83 103
rect 75 99 78 101
rect 80 99 83 101
rect 75 94 83 99
rect 75 92 78 94
rect 80 92 83 94
rect 75 90 83 92
rect 85 94 92 103
rect 99 101 106 106
rect 99 99 101 101
rect 103 99 106 101
rect 99 97 106 99
rect 85 92 88 94
rect 90 92 92 94
rect 101 92 106 97
rect 108 103 114 110
rect 108 96 116 103
rect 108 94 111 96
rect 113 94 116 96
rect 108 92 116 94
rect 85 90 92 92
rect 110 90 116 92
rect 118 101 126 103
rect 118 99 121 101
rect 123 99 126 101
rect 118 94 126 99
rect 118 92 121 94
rect 123 92 126 94
rect 118 90 126 92
rect 128 94 135 103
rect 128 92 131 94
rect 133 92 135 94
rect 128 90 135 92
rect -386 64 -381 71
rect -388 62 -381 64
rect -388 60 -386 62
rect -384 60 -381 62
rect -388 58 -381 60
rect -386 43 -381 58
rect -379 54 -371 71
rect -379 52 -376 54
rect -374 52 -371 54
rect -379 43 -371 52
rect -369 54 -361 71
rect -369 52 -366 54
rect -364 52 -361 54
rect -369 47 -361 52
rect -369 45 -366 47
rect -364 45 -361 47
rect -369 43 -361 45
rect -359 69 -351 71
rect -359 67 -356 69
rect -354 67 -351 69
rect -359 57 -351 67
rect -349 62 -341 71
rect -349 60 -346 62
rect -344 60 -341 62
rect -349 57 -341 60
rect -339 69 -332 71
rect -339 67 -336 69
rect -334 67 -332 69
rect -339 62 -332 67
rect -326 64 -321 71
rect -339 60 -336 62
rect -334 60 -332 62
rect -339 57 -332 60
rect -328 62 -321 64
rect -328 60 -326 62
rect -324 60 -321 62
rect -328 58 -321 60
rect -359 43 -353 57
rect -326 43 -321 58
rect -319 54 -311 71
rect -319 52 -316 54
rect -314 52 -311 54
rect -319 43 -311 52
rect -309 54 -301 71
rect -309 52 -306 54
rect -304 52 -301 54
rect -309 47 -301 52
rect -309 45 -306 47
rect -304 45 -301 47
rect -309 43 -301 45
rect -299 69 -292 71
rect -299 67 -296 69
rect -294 67 -292 69
rect -299 64 -292 67
rect -255 64 -250 71
rect -299 50 -290 64
rect -288 54 -280 64
rect -288 52 -285 54
rect -283 52 -280 54
rect -288 50 -280 52
rect -278 62 -270 64
rect -278 60 -275 62
rect -273 60 -270 62
rect -278 50 -270 60
rect -257 62 -250 64
rect -257 60 -255 62
rect -253 60 -250 62
rect -257 58 -250 60
rect -299 43 -292 50
rect -255 43 -250 58
rect -248 54 -240 71
rect -248 52 -245 54
rect -243 52 -240 54
rect -248 43 -240 52
rect -238 54 -230 71
rect -238 52 -235 54
rect -233 52 -230 54
rect -238 47 -230 52
rect -238 45 -235 47
rect -233 45 -230 47
rect -238 43 -230 45
rect -228 69 -220 71
rect -228 67 -225 69
rect -223 67 -220 69
rect -228 57 -220 67
rect -218 62 -210 71
rect -218 60 -215 62
rect -213 60 -210 62
rect -218 57 -210 60
rect -208 69 -201 71
rect -208 67 -205 69
rect -203 67 -201 69
rect -208 62 -201 67
rect -195 64 -190 71
rect -208 60 -205 62
rect -203 60 -201 62
rect -208 57 -201 60
rect -197 62 -190 64
rect -197 60 -195 62
rect -193 60 -190 62
rect -197 58 -190 60
rect -228 43 -222 57
rect -195 43 -190 58
rect -188 54 -180 71
rect -188 52 -185 54
rect -183 52 -180 54
rect -188 43 -180 52
rect -178 54 -170 71
rect -178 52 -175 54
rect -173 52 -170 54
rect -178 47 -170 52
rect -178 45 -175 47
rect -173 45 -170 47
rect -178 43 -170 45
rect -168 69 -161 71
rect -168 67 -165 69
rect -163 67 -161 69
rect -168 64 -161 67
rect -123 64 -118 71
rect -168 50 -159 64
rect -157 54 -149 64
rect -157 52 -154 54
rect -152 52 -149 54
rect -157 50 -149 52
rect -147 62 -139 64
rect -147 60 -144 62
rect -142 60 -139 62
rect -147 50 -139 60
rect -125 62 -118 64
rect -125 60 -123 62
rect -121 60 -118 62
rect -125 58 -118 60
rect -168 43 -161 50
rect -123 43 -118 58
rect -116 54 -108 71
rect -116 52 -113 54
rect -111 52 -108 54
rect -116 43 -108 52
rect -106 54 -98 71
rect -106 52 -103 54
rect -101 52 -98 54
rect -106 47 -98 52
rect -106 45 -103 47
rect -101 45 -98 47
rect -106 43 -98 45
rect -96 69 -88 71
rect -96 67 -93 69
rect -91 67 -88 69
rect -96 57 -88 67
rect -86 62 -78 71
rect -86 60 -83 62
rect -81 60 -78 62
rect -86 57 -78 60
rect -76 69 -69 71
rect -76 67 -73 69
rect -71 67 -69 69
rect -76 62 -69 67
rect -63 64 -58 71
rect -76 60 -73 62
rect -71 60 -69 62
rect -76 57 -69 60
rect -65 62 -58 64
rect -65 60 -63 62
rect -61 60 -58 62
rect -65 58 -58 60
rect -96 43 -90 57
rect -63 43 -58 58
rect -56 54 -48 71
rect -56 52 -53 54
rect -51 52 -48 54
rect -56 43 -48 52
rect -46 54 -38 71
rect -46 52 -43 54
rect -41 52 -38 54
rect -46 47 -38 52
rect -46 45 -43 47
rect -41 45 -38 47
rect -46 43 -38 45
rect -36 69 -29 71
rect -36 67 -33 69
rect -31 67 -29 69
rect -36 64 -29 67
rect -36 50 -27 64
rect -25 54 -17 64
rect -25 52 -22 54
rect -20 52 -17 54
rect -25 50 -17 52
rect -15 62 -7 64
rect -15 60 -12 62
rect -10 60 -7 62
rect -15 50 -7 60
rect 17 50 22 71
rect -36 43 -29 50
rect 15 48 22 50
rect 15 46 17 48
rect 19 46 22 48
rect 15 44 22 46
rect 24 69 36 71
rect 24 67 27 69
rect 29 67 36 69
rect 24 62 36 67
rect 53 62 58 71
rect 24 60 27 62
rect 29 60 38 62
rect 24 44 38 60
rect 40 55 48 62
rect 40 53 43 55
rect 45 53 48 55
rect 40 48 48 53
rect 40 46 43 48
rect 45 46 48 48
rect 40 44 48 46
rect 50 55 58 62
rect 50 53 53 55
rect 55 53 58 55
rect 50 44 58 53
rect 60 65 65 71
rect 60 63 67 65
rect 60 61 63 63
rect 65 61 67 63
rect 60 59 67 61
rect 60 44 65 59
rect -378 -34 -371 -32
rect -378 -36 -376 -34
rect -374 -36 -371 -34
rect -378 -41 -371 -36
rect -378 -43 -376 -41
rect -374 -43 -371 -41
rect -378 -45 -371 -43
rect -376 -50 -371 -45
rect -369 -49 -360 -32
rect -347 -40 -342 -32
rect -369 -50 -365 -49
rect -367 -51 -365 -50
rect -363 -51 -360 -49
rect -367 -53 -360 -51
rect -349 -42 -342 -40
rect -349 -44 -347 -42
rect -345 -44 -342 -42
rect -349 -49 -342 -44
rect -349 -51 -347 -49
rect -345 -51 -342 -49
rect -349 -53 -342 -51
rect -347 -59 -342 -53
rect -340 -48 -332 -32
rect -340 -50 -337 -48
rect -335 -50 -332 -48
rect -340 -55 -332 -50
rect -340 -57 -337 -55
rect -335 -57 -332 -55
rect -340 -59 -332 -57
rect -330 -59 -325 -32
rect -323 -34 -315 -32
rect -323 -36 -320 -34
rect -318 -36 -315 -34
rect -323 -41 -315 -36
rect -323 -43 -320 -41
rect -318 -43 -315 -41
rect -323 -59 -315 -43
rect -313 -50 -305 -32
rect -313 -52 -310 -50
rect -308 -52 -305 -50
rect -313 -59 -305 -52
rect -303 -47 -296 -32
rect -284 -34 -277 -32
rect -284 -36 -282 -34
rect -280 -36 -277 -34
rect -284 -41 -277 -36
rect -284 -43 -282 -41
rect -280 -43 -277 -41
rect -284 -45 -277 -43
rect -303 -49 -300 -47
rect -298 -49 -296 -47
rect -303 -55 -296 -49
rect -282 -50 -277 -45
rect -275 -49 -266 -32
rect -251 -40 -246 -32
rect -275 -50 -271 -49
rect -273 -51 -271 -50
rect -269 -51 -266 -49
rect -273 -53 -266 -51
rect -253 -42 -246 -40
rect -253 -44 -251 -42
rect -249 -44 -246 -42
rect -253 -49 -246 -44
rect -253 -51 -251 -49
rect -249 -51 -246 -49
rect -253 -53 -246 -51
rect -303 -57 -300 -55
rect -298 -57 -296 -55
rect -303 -59 -296 -57
rect -251 -59 -246 -53
rect -244 -48 -236 -32
rect -244 -50 -241 -48
rect -239 -50 -236 -48
rect -244 -55 -236 -50
rect -244 -57 -241 -55
rect -239 -57 -236 -55
rect -244 -59 -236 -57
rect -234 -59 -229 -32
rect -227 -34 -219 -32
rect -227 -36 -224 -34
rect -222 -36 -219 -34
rect -227 -41 -219 -36
rect -227 -43 -224 -41
rect -222 -43 -219 -41
rect -227 -59 -219 -43
rect -217 -50 -209 -32
rect -217 -52 -214 -50
rect -212 -52 -209 -50
rect -217 -59 -209 -52
rect -207 -47 -200 -32
rect -151 -35 -144 -33
rect -151 -37 -149 -35
rect -147 -37 -144 -35
rect -151 -42 -144 -37
rect -151 -44 -149 -42
rect -147 -44 -144 -42
rect -151 -46 -144 -44
rect -207 -49 -204 -47
rect -202 -49 -200 -47
rect -207 -55 -200 -49
rect -149 -51 -144 -46
rect -142 -50 -133 -33
rect -119 -41 -114 -33
rect -142 -51 -138 -50
rect -207 -57 -204 -55
rect -202 -57 -200 -55
rect -140 -52 -138 -51
rect -136 -52 -133 -50
rect -140 -54 -133 -52
rect -121 -43 -114 -41
rect -121 -45 -119 -43
rect -117 -45 -114 -43
rect -121 -50 -114 -45
rect -121 -52 -119 -50
rect -117 -52 -114 -50
rect -121 -54 -114 -52
rect -207 -59 -200 -57
rect -119 -60 -114 -54
rect -112 -49 -104 -33
rect -112 -51 -109 -49
rect -107 -51 -104 -49
rect -112 -56 -104 -51
rect -112 -58 -109 -56
rect -107 -58 -104 -56
rect -112 -60 -104 -58
rect -102 -60 -97 -33
rect -95 -35 -87 -33
rect -95 -37 -92 -35
rect -90 -37 -87 -35
rect -95 -42 -87 -37
rect -95 -44 -92 -42
rect -90 -44 -87 -42
rect -95 -60 -87 -44
rect -85 -51 -77 -33
rect -85 -53 -82 -51
rect -80 -53 -77 -51
rect -85 -60 -77 -53
rect -75 -48 -68 -33
rect 9 -36 16 -34
rect 9 -38 11 -36
rect 13 -38 16 -36
rect 9 -43 16 -38
rect 9 -45 11 -43
rect 13 -45 16 -43
rect 9 -47 16 -45
rect -75 -50 -72 -48
rect -70 -50 -68 -48
rect -75 -56 -68 -50
rect 11 -52 16 -47
rect 18 -41 24 -34
rect 18 -48 26 -41
rect 18 -50 21 -48
rect 23 -50 26 -48
rect 18 -52 26 -50
rect 20 -54 26 -52
rect 28 -43 36 -41
rect 28 -45 31 -43
rect 33 -45 36 -43
rect 28 -50 36 -45
rect 28 -52 31 -50
rect 33 -52 36 -50
rect 28 -54 36 -52
rect 38 -50 45 -41
rect 38 -52 41 -50
rect 43 -52 45 -50
rect 38 -54 45 -52
rect -75 -58 -72 -56
rect -70 -58 -68 -56
rect -75 -60 -68 -58
rect -439 -83 -432 -81
rect -411 -82 -405 -80
rect -439 -84 -437 -83
rect -448 -89 -443 -84
rect -450 -91 -443 -89
rect -450 -93 -448 -91
rect -446 -93 -443 -91
rect -450 -98 -443 -93
rect -450 -100 -448 -98
rect -446 -100 -443 -98
rect -450 -102 -443 -100
rect -441 -85 -437 -84
rect -435 -85 -432 -83
rect -441 -102 -432 -85
rect -420 -87 -415 -82
rect -422 -89 -415 -87
rect -422 -91 -420 -89
rect -418 -91 -415 -89
rect -422 -96 -415 -91
rect -422 -98 -420 -96
rect -418 -98 -415 -96
rect -422 -100 -415 -98
rect -413 -84 -405 -82
rect -413 -86 -410 -84
rect -408 -86 -405 -84
rect -413 -93 -405 -86
rect -403 -82 -395 -80
rect -403 -84 -400 -82
rect -398 -84 -395 -82
rect -403 -89 -395 -84
rect -403 -91 -400 -89
rect -398 -91 -395 -89
rect -403 -93 -395 -91
rect -393 -82 -386 -80
rect -299 -81 -293 -79
rect -393 -84 -390 -82
rect -388 -84 -386 -82
rect -393 -93 -386 -84
rect -308 -86 -303 -81
rect -310 -88 -303 -86
rect -310 -90 -308 -88
rect -306 -90 -303 -88
rect -413 -100 -407 -93
rect -310 -95 -303 -90
rect -310 -97 -308 -95
rect -306 -97 -303 -95
rect -310 -99 -303 -97
rect -301 -83 -293 -81
rect -301 -85 -298 -83
rect -296 -85 -293 -83
rect -301 -92 -293 -85
rect -291 -81 -283 -79
rect -291 -83 -288 -81
rect -286 -83 -283 -81
rect -291 -88 -283 -83
rect -291 -90 -288 -88
rect -286 -90 -283 -88
rect -291 -92 -283 -90
rect -281 -81 -274 -79
rect -281 -83 -278 -81
rect -276 -83 -274 -81
rect -148 -82 -142 -80
rect -281 -92 -274 -83
rect -157 -87 -152 -82
rect -159 -89 -152 -87
rect -159 -91 -157 -89
rect -155 -91 -152 -89
rect -301 -99 -295 -92
rect -159 -96 -152 -91
rect -159 -98 -157 -96
rect -155 -98 -152 -96
rect -159 -100 -152 -98
rect -150 -84 -142 -82
rect -150 -86 -147 -84
rect -145 -86 -142 -84
rect -150 -93 -142 -86
rect -140 -82 -132 -80
rect -140 -84 -137 -82
rect -135 -84 -132 -82
rect -140 -89 -132 -84
rect -140 -91 -137 -89
rect -135 -91 -132 -89
rect -140 -93 -132 -91
rect -130 -82 -123 -80
rect -104 -82 -98 -80
rect -130 -84 -127 -82
rect -125 -84 -123 -82
rect -130 -93 -123 -84
rect -113 -87 -108 -82
rect -115 -89 -108 -87
rect -115 -91 -113 -89
rect -111 -91 -108 -89
rect -150 -100 -144 -93
rect -115 -96 -108 -91
rect -115 -98 -113 -96
rect -111 -98 -108 -96
rect -115 -100 -108 -98
rect -106 -84 -98 -82
rect -106 -86 -103 -84
rect -101 -86 -98 -84
rect -106 -93 -98 -86
rect -96 -82 -88 -80
rect -96 -84 -93 -82
rect -91 -84 -88 -82
rect -96 -89 -88 -84
rect -96 -91 -93 -89
rect -91 -91 -88 -89
rect -96 -93 -88 -91
rect -86 -82 -79 -80
rect -86 -84 -83 -82
rect -81 -84 -79 -82
rect -86 -93 -79 -84
rect -106 -100 -100 -93
rect -539 -193 -534 -178
rect -541 -195 -534 -193
rect -541 -197 -539 -195
rect -537 -197 -534 -195
rect -541 -199 -534 -197
rect -539 -206 -534 -199
rect -532 -187 -524 -178
rect -532 -189 -529 -187
rect -527 -189 -524 -187
rect -532 -206 -524 -189
rect -522 -180 -514 -178
rect -522 -182 -519 -180
rect -517 -182 -514 -180
rect -522 -187 -514 -182
rect -522 -189 -519 -187
rect -517 -189 -514 -187
rect -522 -206 -514 -189
rect -512 -192 -506 -178
rect -512 -202 -504 -192
rect -512 -204 -509 -202
rect -507 -204 -504 -202
rect -512 -206 -504 -204
rect -502 -195 -494 -192
rect -502 -197 -499 -195
rect -497 -197 -494 -195
rect -502 -206 -494 -197
rect -492 -195 -485 -192
rect -479 -193 -474 -178
rect -492 -197 -489 -195
rect -487 -197 -485 -195
rect -492 -202 -485 -197
rect -481 -195 -474 -193
rect -481 -197 -479 -195
rect -477 -197 -474 -195
rect -481 -199 -474 -197
rect -492 -204 -489 -202
rect -487 -204 -485 -202
rect -492 -206 -485 -204
rect -479 -206 -474 -199
rect -472 -187 -464 -178
rect -472 -189 -469 -187
rect -467 -189 -464 -187
rect -472 -206 -464 -189
rect -462 -180 -454 -178
rect -462 -182 -459 -180
rect -457 -182 -454 -180
rect -462 -187 -454 -182
rect -462 -189 -459 -187
rect -457 -189 -454 -187
rect -462 -206 -454 -189
rect -452 -185 -445 -178
rect -452 -199 -443 -185
rect -441 -187 -433 -185
rect -441 -189 -438 -187
rect -436 -189 -433 -187
rect -441 -199 -433 -189
rect -431 -195 -423 -185
rect -407 -193 -402 -178
rect -431 -197 -428 -195
rect -426 -197 -423 -195
rect -431 -199 -423 -197
rect -409 -195 -402 -193
rect -409 -197 -407 -195
rect -405 -197 -402 -195
rect -409 -199 -402 -197
rect -452 -202 -445 -199
rect -452 -204 -449 -202
rect -447 -204 -445 -202
rect -452 -206 -445 -204
rect -407 -206 -402 -199
rect -400 -187 -392 -178
rect -400 -189 -397 -187
rect -395 -189 -392 -187
rect -400 -206 -392 -189
rect -390 -180 -382 -178
rect -390 -182 -387 -180
rect -385 -182 -382 -180
rect -390 -187 -382 -182
rect -390 -189 -387 -187
rect -385 -189 -382 -187
rect -390 -206 -382 -189
rect -380 -192 -374 -178
rect -380 -202 -372 -192
rect -380 -204 -377 -202
rect -375 -204 -372 -202
rect -380 -206 -372 -204
rect -370 -195 -362 -192
rect -370 -197 -367 -195
rect -365 -197 -362 -195
rect -370 -206 -362 -197
rect -360 -195 -353 -192
rect -347 -193 -342 -178
rect -360 -197 -357 -195
rect -355 -197 -353 -195
rect -360 -202 -353 -197
rect -349 -195 -342 -193
rect -349 -197 -347 -195
rect -345 -197 -342 -195
rect -349 -199 -342 -197
rect -360 -204 -357 -202
rect -355 -204 -353 -202
rect -360 -206 -353 -204
rect -347 -206 -342 -199
rect -340 -187 -332 -178
rect -340 -189 -337 -187
rect -335 -189 -332 -187
rect -340 -206 -332 -189
rect -330 -180 -322 -178
rect -330 -182 -327 -180
rect -325 -182 -322 -180
rect -330 -187 -322 -182
rect -330 -189 -327 -187
rect -325 -189 -322 -187
rect -330 -206 -322 -189
rect -320 -185 -313 -178
rect -320 -199 -311 -185
rect -309 -187 -301 -185
rect -309 -189 -306 -187
rect -304 -189 -301 -187
rect -309 -199 -301 -189
rect -299 -195 -291 -185
rect -270 -192 -265 -177
rect -299 -197 -296 -195
rect -294 -197 -291 -195
rect -299 -199 -291 -197
rect -272 -194 -265 -192
rect -272 -196 -270 -194
rect -268 -196 -265 -194
rect -272 -198 -265 -196
rect -320 -202 -313 -199
rect -320 -204 -317 -202
rect -315 -204 -313 -202
rect -320 -206 -313 -204
rect -270 -205 -265 -198
rect -263 -186 -255 -177
rect -263 -188 -260 -186
rect -258 -188 -255 -186
rect -263 -205 -255 -188
rect -253 -179 -245 -177
rect -253 -181 -250 -179
rect -248 -181 -245 -179
rect -253 -186 -245 -181
rect -253 -188 -250 -186
rect -248 -188 -245 -186
rect -253 -205 -245 -188
rect -243 -191 -237 -177
rect -243 -201 -235 -191
rect -243 -203 -240 -201
rect -238 -203 -235 -201
rect -243 -205 -235 -203
rect -233 -194 -225 -191
rect -233 -196 -230 -194
rect -228 -196 -225 -194
rect -233 -205 -225 -196
rect -223 -194 -216 -191
rect -210 -192 -205 -177
rect -223 -196 -220 -194
rect -218 -196 -216 -194
rect -223 -201 -216 -196
rect -212 -194 -205 -192
rect -212 -196 -210 -194
rect -208 -196 -205 -194
rect -212 -198 -205 -196
rect -223 -203 -220 -201
rect -218 -203 -216 -201
rect -223 -205 -216 -203
rect -210 -205 -205 -198
rect -203 -186 -195 -177
rect -203 -188 -200 -186
rect -198 -188 -195 -186
rect -203 -205 -195 -188
rect -193 -179 -185 -177
rect -193 -181 -190 -179
rect -188 -181 -185 -179
rect -193 -186 -185 -181
rect -193 -188 -190 -186
rect -188 -188 -185 -186
rect -193 -205 -185 -188
rect -183 -184 -176 -177
rect -183 -198 -174 -184
rect -172 -186 -164 -184
rect -172 -188 -169 -186
rect -167 -188 -164 -186
rect -172 -198 -164 -188
rect -162 -194 -154 -184
rect -139 -193 -134 -178
rect -162 -196 -159 -194
rect -157 -196 -154 -194
rect -162 -198 -154 -196
rect -141 -195 -134 -193
rect -141 -197 -139 -195
rect -137 -197 -134 -195
rect -183 -201 -176 -198
rect -183 -203 -180 -201
rect -178 -203 -176 -201
rect -141 -199 -134 -197
rect -183 -205 -176 -203
rect -139 -205 -134 -199
rect -132 -187 -124 -178
rect -132 -189 -129 -187
rect -127 -189 -124 -187
rect -132 -196 -124 -189
rect -122 -180 -114 -178
rect -122 -182 -119 -180
rect -117 -182 -114 -180
rect -122 -187 -114 -182
rect -122 -189 -119 -187
rect -117 -189 -114 -187
rect -122 -196 -114 -189
rect -112 -194 -98 -178
rect -112 -196 -103 -194
rect -101 -196 -98 -194
rect -132 -205 -127 -196
rect -110 -201 -98 -196
rect -110 -203 -103 -201
rect -101 -203 -98 -201
rect -110 -205 -98 -203
rect -96 -180 -89 -178
rect -96 -182 -93 -180
rect -91 -182 -89 -180
rect -96 -184 -89 -182
rect -96 -205 -91 -184
rect -471 -225 -466 -219
rect -491 -227 -484 -225
rect -491 -228 -489 -227
rect -500 -233 -495 -228
rect -502 -235 -495 -233
rect -502 -237 -500 -235
rect -498 -237 -495 -235
rect -502 -242 -495 -237
rect -502 -244 -500 -242
rect -498 -244 -495 -242
rect -502 -246 -495 -244
rect -493 -229 -489 -228
rect -487 -229 -484 -227
rect -493 -246 -484 -229
rect -473 -227 -466 -225
rect -473 -229 -471 -227
rect -469 -229 -466 -227
rect -473 -234 -466 -229
rect -473 -236 -471 -234
rect -469 -236 -466 -234
rect -473 -238 -466 -236
rect -471 -246 -466 -238
rect -464 -221 -456 -219
rect -464 -223 -461 -221
rect -459 -223 -456 -221
rect -464 -228 -456 -223
rect -464 -230 -461 -228
rect -459 -230 -456 -228
rect -464 -246 -456 -230
rect -454 -246 -449 -219
rect -447 -235 -439 -219
rect -447 -237 -444 -235
rect -442 -237 -439 -235
rect -447 -242 -439 -237
rect -447 -244 -444 -242
rect -442 -244 -439 -242
rect -447 -246 -439 -244
rect -437 -226 -429 -219
rect -437 -228 -434 -226
rect -432 -228 -429 -226
rect -437 -246 -429 -228
rect -427 -221 -420 -219
rect -427 -223 -424 -221
rect -422 -223 -420 -221
rect -427 -229 -420 -223
rect -377 -225 -372 -219
rect -398 -227 -391 -225
rect -398 -228 -396 -227
rect -427 -231 -424 -229
rect -422 -231 -420 -229
rect -427 -246 -420 -231
rect -407 -233 -402 -228
rect -409 -235 -402 -233
rect -409 -237 -407 -235
rect -405 -237 -402 -235
rect -409 -242 -402 -237
rect -409 -244 -407 -242
rect -405 -244 -402 -242
rect -409 -246 -402 -244
rect -400 -229 -396 -228
rect -394 -229 -391 -227
rect -400 -246 -391 -229
rect -379 -227 -372 -225
rect -379 -229 -377 -227
rect -375 -229 -372 -227
rect -379 -234 -372 -229
rect -379 -236 -377 -234
rect -375 -236 -372 -234
rect -379 -238 -372 -236
rect -377 -246 -372 -238
rect -370 -221 -362 -219
rect -370 -223 -367 -221
rect -365 -223 -362 -221
rect -370 -228 -362 -223
rect -370 -230 -367 -228
rect -365 -230 -362 -228
rect -370 -246 -362 -230
rect -360 -246 -355 -219
rect -353 -235 -345 -219
rect -353 -237 -350 -235
rect -348 -237 -345 -235
rect -353 -242 -345 -237
rect -353 -244 -350 -242
rect -348 -244 -345 -242
rect -353 -246 -345 -244
rect -343 -226 -335 -219
rect -343 -228 -340 -226
rect -338 -228 -335 -226
rect -343 -246 -335 -228
rect -333 -221 -326 -219
rect -333 -223 -330 -221
rect -328 -223 -326 -221
rect -333 -229 -326 -223
rect -203 -224 -198 -218
rect -225 -226 -218 -224
rect -225 -227 -223 -226
rect -333 -231 -330 -229
rect -328 -231 -326 -229
rect -333 -246 -326 -231
rect -234 -232 -229 -227
rect -236 -234 -229 -232
rect -236 -236 -234 -234
rect -232 -236 -229 -234
rect -236 -241 -229 -236
rect -236 -243 -234 -241
rect -232 -243 -229 -241
rect -236 -245 -229 -243
rect -227 -228 -223 -227
rect -221 -228 -218 -226
rect -227 -245 -218 -228
rect -205 -226 -198 -224
rect -205 -228 -203 -226
rect -201 -228 -198 -226
rect -205 -233 -198 -228
rect -205 -235 -203 -233
rect -201 -235 -198 -233
rect -205 -237 -198 -235
rect -203 -245 -198 -237
rect -196 -220 -188 -218
rect -196 -222 -193 -220
rect -191 -222 -188 -220
rect -196 -227 -188 -222
rect -196 -229 -193 -227
rect -191 -229 -188 -227
rect -196 -245 -188 -229
rect -186 -245 -181 -218
rect -179 -234 -171 -218
rect -179 -236 -176 -234
rect -174 -236 -171 -234
rect -179 -241 -171 -236
rect -179 -243 -176 -241
rect -174 -243 -171 -241
rect -179 -245 -171 -243
rect -169 -225 -161 -218
rect -169 -227 -166 -225
rect -164 -227 -161 -225
rect -169 -245 -161 -227
rect -159 -220 -152 -218
rect -159 -222 -156 -220
rect -154 -222 -152 -220
rect -159 -228 -152 -222
rect -130 -226 -124 -224
rect -159 -230 -156 -228
rect -154 -230 -152 -228
rect -159 -245 -152 -230
rect -139 -231 -134 -226
rect -141 -233 -134 -231
rect -141 -235 -139 -233
rect -137 -235 -134 -233
rect -141 -240 -134 -235
rect -141 -242 -139 -240
rect -137 -242 -134 -240
rect -141 -244 -134 -242
rect -132 -228 -124 -226
rect -132 -230 -129 -228
rect -127 -230 -124 -228
rect -132 -237 -124 -230
rect -122 -226 -114 -224
rect -122 -228 -119 -226
rect -117 -228 -114 -226
rect -122 -233 -114 -228
rect -122 -235 -119 -233
rect -117 -235 -114 -233
rect -122 -237 -114 -235
rect -112 -226 -105 -224
rect -112 -228 -109 -226
rect -107 -228 -105 -226
rect -112 -237 -105 -228
rect -132 -244 -126 -237
rect -578 -325 -571 -323
rect -578 -327 -576 -325
rect -574 -327 -571 -325
rect -578 -332 -571 -327
rect -578 -334 -576 -332
rect -574 -334 -571 -332
rect -578 -336 -571 -334
rect -576 -341 -571 -336
rect -569 -330 -563 -323
rect -569 -337 -561 -330
rect -569 -339 -566 -337
rect -564 -339 -561 -337
rect -569 -341 -561 -339
rect -567 -343 -561 -341
rect -559 -332 -551 -330
rect -559 -334 -556 -332
rect -554 -334 -551 -332
rect -559 -339 -551 -334
rect -559 -341 -556 -339
rect -554 -341 -551 -339
rect -559 -343 -551 -341
rect -549 -339 -542 -330
rect -549 -341 -546 -339
rect -544 -341 -542 -339
rect -549 -343 -542 -341
rect -505 -339 -497 -327
rect -505 -341 -503 -339
rect -501 -341 -497 -339
rect -495 -330 -487 -327
rect -495 -332 -492 -330
rect -490 -332 -487 -330
rect -495 -337 -487 -332
rect -495 -339 -492 -337
rect -490 -339 -487 -337
rect -495 -341 -487 -339
rect -485 -330 -477 -327
rect -485 -332 -481 -330
rect -479 -332 -477 -330
rect -485 -337 -477 -332
rect -485 -339 -481 -337
rect -479 -339 -477 -337
rect -485 -341 -477 -339
rect -381 -339 -373 -327
rect -381 -341 -379 -339
rect -377 -341 -373 -339
rect -371 -330 -363 -327
rect -371 -332 -368 -330
rect -366 -332 -363 -330
rect -371 -337 -363 -332
rect -371 -339 -368 -337
rect -366 -339 -363 -337
rect -371 -341 -363 -339
rect -361 -330 -353 -327
rect -361 -332 -357 -330
rect -355 -332 -353 -330
rect -361 -337 -353 -332
rect -361 -339 -357 -337
rect -355 -339 -353 -337
rect -361 -341 -353 -339
rect -235 -338 -227 -326
rect -235 -340 -233 -338
rect -231 -340 -227 -338
rect -225 -329 -217 -326
rect -225 -331 -222 -329
rect -220 -331 -217 -329
rect -225 -336 -217 -331
rect -225 -338 -222 -336
rect -220 -338 -217 -336
rect -225 -340 -217 -338
rect -215 -329 -207 -326
rect -215 -331 -211 -329
rect -209 -331 -207 -329
rect -215 -336 -207 -331
rect -215 -338 -211 -336
rect -209 -338 -207 -336
rect -215 -340 -207 -338
rect -505 -343 -499 -341
rect -381 -343 -375 -341
rect -235 -342 -229 -340
rect -717 -368 -712 -361
rect -719 -370 -712 -368
rect -719 -372 -717 -370
rect -715 -372 -712 -370
rect -719 -374 -712 -372
rect -717 -389 -712 -374
rect -710 -378 -702 -361
rect -710 -380 -707 -378
rect -705 -380 -702 -378
rect -710 -389 -702 -380
rect -700 -378 -692 -361
rect -700 -380 -697 -378
rect -695 -380 -692 -378
rect -700 -385 -692 -380
rect -700 -387 -697 -385
rect -695 -387 -692 -385
rect -700 -389 -692 -387
rect -690 -363 -682 -361
rect -690 -365 -687 -363
rect -685 -365 -682 -363
rect -690 -375 -682 -365
rect -680 -370 -672 -361
rect -680 -372 -677 -370
rect -675 -372 -672 -370
rect -680 -375 -672 -372
rect -670 -363 -663 -361
rect -670 -365 -667 -363
rect -665 -365 -663 -363
rect -670 -370 -663 -365
rect -657 -368 -652 -361
rect -670 -372 -667 -370
rect -665 -372 -663 -370
rect -670 -375 -663 -372
rect -659 -370 -652 -368
rect -659 -372 -657 -370
rect -655 -372 -652 -370
rect -659 -374 -652 -372
rect -690 -389 -684 -375
rect -657 -389 -652 -374
rect -650 -378 -642 -361
rect -650 -380 -647 -378
rect -645 -380 -642 -378
rect -650 -389 -642 -380
rect -640 -378 -632 -361
rect -640 -380 -637 -378
rect -635 -380 -632 -378
rect -640 -385 -632 -380
rect -640 -387 -637 -385
rect -635 -387 -632 -385
rect -640 -389 -632 -387
rect -630 -363 -623 -361
rect -630 -365 -627 -363
rect -625 -365 -623 -363
rect -630 -368 -623 -365
rect -585 -368 -580 -361
rect -630 -382 -621 -368
rect -619 -378 -611 -368
rect -619 -380 -616 -378
rect -614 -380 -611 -378
rect -619 -382 -611 -380
rect -609 -370 -601 -368
rect -609 -372 -606 -370
rect -604 -372 -601 -370
rect -609 -382 -601 -372
rect -587 -370 -580 -368
rect -587 -372 -585 -370
rect -583 -372 -580 -370
rect -587 -374 -580 -372
rect -630 -389 -623 -382
rect -585 -389 -580 -374
rect -578 -378 -570 -361
rect -578 -380 -575 -378
rect -573 -380 -570 -378
rect -578 -389 -570 -380
rect -568 -378 -560 -361
rect -568 -380 -565 -378
rect -563 -380 -560 -378
rect -568 -385 -560 -380
rect -568 -387 -565 -385
rect -563 -387 -560 -385
rect -568 -389 -560 -387
rect -558 -363 -550 -361
rect -558 -365 -555 -363
rect -553 -365 -550 -363
rect -558 -375 -550 -365
rect -548 -370 -540 -361
rect -548 -372 -545 -370
rect -543 -372 -540 -370
rect -548 -375 -540 -372
rect -538 -363 -531 -361
rect -538 -365 -535 -363
rect -533 -365 -531 -363
rect -538 -370 -531 -365
rect -525 -368 -520 -361
rect -538 -372 -535 -370
rect -533 -372 -531 -370
rect -538 -375 -531 -372
rect -527 -370 -520 -368
rect -527 -372 -525 -370
rect -523 -372 -520 -370
rect -527 -374 -520 -372
rect -558 -389 -552 -375
rect -525 -389 -520 -374
rect -518 -378 -510 -361
rect -518 -380 -515 -378
rect -513 -380 -510 -378
rect -518 -389 -510 -380
rect -508 -378 -500 -361
rect -508 -380 -505 -378
rect -503 -380 -500 -378
rect -508 -385 -500 -380
rect -508 -387 -505 -385
rect -503 -387 -500 -385
rect -508 -389 -500 -387
rect -498 -363 -491 -361
rect -498 -365 -495 -363
rect -493 -365 -491 -363
rect -498 -368 -491 -365
rect -453 -368 -448 -361
rect -498 -382 -489 -368
rect -487 -378 -479 -368
rect -487 -380 -484 -378
rect -482 -380 -479 -378
rect -487 -382 -479 -380
rect -477 -370 -469 -368
rect -477 -372 -474 -370
rect -472 -372 -469 -370
rect -477 -382 -469 -372
rect -455 -370 -448 -368
rect -455 -372 -453 -370
rect -451 -372 -448 -370
rect -455 -374 -448 -372
rect -498 -389 -491 -382
rect -453 -389 -448 -374
rect -446 -378 -438 -361
rect -446 -380 -443 -378
rect -441 -380 -438 -378
rect -446 -389 -438 -380
rect -436 -378 -428 -361
rect -436 -380 -433 -378
rect -431 -380 -428 -378
rect -436 -385 -428 -380
rect -436 -387 -433 -385
rect -431 -387 -428 -385
rect -436 -389 -428 -387
rect -426 -363 -418 -361
rect -426 -365 -423 -363
rect -421 -365 -418 -363
rect -426 -375 -418 -365
rect -416 -370 -408 -361
rect -416 -372 -413 -370
rect -411 -372 -408 -370
rect -416 -375 -408 -372
rect -406 -363 -399 -361
rect -406 -365 -403 -363
rect -401 -365 -399 -363
rect -406 -370 -399 -365
rect -393 -368 -388 -361
rect -406 -372 -403 -370
rect -401 -372 -399 -370
rect -406 -375 -399 -372
rect -395 -370 -388 -368
rect -395 -372 -393 -370
rect -391 -372 -388 -370
rect -395 -374 -388 -372
rect -426 -389 -420 -375
rect -393 -389 -388 -374
rect -386 -378 -378 -361
rect -386 -380 -383 -378
rect -381 -380 -378 -378
rect -386 -389 -378 -380
rect -376 -378 -368 -361
rect -376 -380 -373 -378
rect -371 -380 -368 -378
rect -376 -385 -368 -380
rect -376 -387 -373 -385
rect -371 -387 -368 -385
rect -376 -389 -368 -387
rect -366 -363 -359 -361
rect -366 -365 -363 -363
rect -361 -365 -359 -363
rect -366 -368 -359 -365
rect -366 -382 -357 -368
rect -355 -378 -347 -368
rect -355 -380 -352 -378
rect -350 -380 -347 -378
rect -355 -382 -347 -380
rect -345 -370 -337 -368
rect -345 -372 -342 -370
rect -340 -372 -337 -370
rect -345 -382 -337 -372
rect -251 -380 -246 -359
rect -253 -382 -246 -380
rect -366 -389 -359 -382
rect -253 -384 -251 -382
rect -249 -384 -246 -382
rect -253 -386 -246 -384
rect -244 -361 -232 -359
rect -244 -363 -241 -361
rect -239 -363 -232 -361
rect -244 -368 -232 -363
rect -215 -368 -210 -359
rect -244 -370 -241 -368
rect -239 -370 -230 -368
rect -244 -386 -230 -370
rect -228 -375 -220 -368
rect -228 -377 -225 -375
rect -223 -377 -220 -375
rect -228 -382 -220 -377
rect -228 -384 -225 -382
rect -223 -384 -220 -382
rect -228 -386 -220 -384
rect -218 -375 -210 -368
rect -218 -377 -215 -375
rect -213 -377 -210 -375
rect -218 -386 -210 -377
rect -208 -365 -203 -359
rect -208 -367 -201 -365
rect -208 -369 -205 -367
rect -203 -369 -201 -367
rect -208 -371 -201 -369
rect -208 -386 -203 -371
rect -785 -480 -780 -465
rect -787 -482 -780 -480
rect -787 -484 -785 -482
rect -783 -484 -780 -482
rect -787 -486 -780 -484
rect -785 -492 -780 -486
rect -778 -474 -770 -465
rect -778 -476 -775 -474
rect -773 -476 -770 -474
rect -778 -483 -770 -476
rect -768 -467 -760 -465
rect -768 -469 -765 -467
rect -763 -469 -760 -467
rect -768 -474 -760 -469
rect -768 -476 -765 -474
rect -763 -476 -760 -474
rect -768 -483 -760 -476
rect -758 -481 -744 -465
rect -758 -483 -749 -481
rect -747 -483 -744 -481
rect -778 -492 -773 -483
rect -756 -488 -744 -483
rect -756 -490 -749 -488
rect -747 -490 -744 -488
rect -756 -492 -744 -490
rect -742 -467 -735 -465
rect -742 -469 -739 -467
rect -737 -469 -735 -467
rect -719 -466 -712 -464
rect -719 -468 -717 -466
rect -715 -468 -712 -466
rect -742 -471 -735 -469
rect -742 -492 -737 -471
rect -719 -473 -712 -468
rect -719 -475 -717 -473
rect -715 -475 -712 -473
rect -719 -477 -712 -475
rect -717 -482 -712 -477
rect -710 -481 -701 -464
rect -686 -473 -681 -465
rect -710 -482 -706 -481
rect -708 -483 -706 -482
rect -704 -483 -701 -481
rect -708 -485 -701 -483
rect -688 -475 -681 -473
rect -688 -477 -686 -475
rect -684 -477 -681 -475
rect -688 -482 -681 -477
rect -688 -484 -686 -482
rect -684 -484 -681 -482
rect -688 -486 -681 -484
rect -686 -492 -681 -486
rect -679 -481 -671 -465
rect -679 -483 -676 -481
rect -674 -483 -671 -481
rect -679 -488 -671 -483
rect -679 -490 -676 -488
rect -674 -490 -671 -488
rect -679 -492 -671 -490
rect -669 -492 -664 -465
rect -662 -467 -654 -465
rect -662 -469 -659 -467
rect -657 -469 -654 -467
rect -662 -474 -654 -469
rect -662 -476 -659 -474
rect -657 -476 -654 -474
rect -662 -492 -654 -476
rect -652 -483 -644 -465
rect -652 -485 -649 -483
rect -647 -485 -644 -483
rect -652 -492 -644 -485
rect -642 -480 -635 -465
rect -587 -467 -580 -465
rect -587 -469 -585 -467
rect -583 -469 -580 -467
rect -587 -474 -580 -469
rect -587 -476 -585 -474
rect -583 -476 -580 -474
rect -587 -478 -580 -476
rect -642 -482 -639 -480
rect -637 -482 -635 -480
rect -642 -488 -635 -482
rect -585 -483 -580 -478
rect -578 -482 -569 -465
rect -554 -473 -549 -465
rect -578 -483 -574 -482
rect -576 -484 -574 -483
rect -572 -484 -569 -482
rect -576 -486 -569 -484
rect -556 -475 -549 -473
rect -556 -477 -554 -475
rect -552 -477 -549 -475
rect -556 -482 -549 -477
rect -556 -484 -554 -482
rect -552 -484 -549 -482
rect -556 -486 -549 -484
rect -642 -490 -639 -488
rect -637 -490 -635 -488
rect -642 -492 -635 -490
rect -554 -492 -549 -486
rect -547 -481 -539 -465
rect -547 -483 -544 -481
rect -542 -483 -539 -481
rect -547 -488 -539 -483
rect -547 -490 -544 -488
rect -542 -490 -539 -488
rect -547 -492 -539 -490
rect -537 -492 -532 -465
rect -530 -467 -522 -465
rect -530 -469 -527 -467
rect -525 -469 -522 -467
rect -530 -474 -522 -469
rect -530 -476 -527 -474
rect -525 -476 -522 -474
rect -530 -492 -522 -476
rect -520 -483 -512 -465
rect -520 -485 -517 -483
rect -515 -485 -512 -483
rect -520 -492 -512 -485
rect -510 -480 -503 -465
rect -455 -466 -448 -464
rect -455 -468 -453 -466
rect -451 -468 -448 -466
rect -455 -473 -448 -468
rect -455 -475 -453 -473
rect -451 -475 -448 -473
rect -455 -477 -448 -475
rect -510 -482 -507 -480
rect -505 -482 -503 -480
rect -453 -482 -448 -477
rect -446 -481 -437 -464
rect -425 -472 -420 -464
rect -446 -482 -442 -481
rect -510 -488 -503 -482
rect -444 -483 -442 -482
rect -440 -483 -437 -481
rect -444 -485 -437 -483
rect -427 -474 -420 -472
rect -427 -476 -425 -474
rect -423 -476 -420 -474
rect -427 -481 -420 -476
rect -427 -483 -425 -481
rect -423 -483 -420 -481
rect -427 -485 -420 -483
rect -510 -490 -507 -488
rect -505 -490 -503 -488
rect -510 -492 -503 -490
rect -425 -491 -420 -485
rect -418 -480 -410 -464
rect -418 -482 -415 -480
rect -413 -482 -410 -480
rect -418 -487 -410 -482
rect -418 -489 -415 -487
rect -413 -489 -410 -487
rect -418 -491 -410 -489
rect -408 -491 -403 -464
rect -401 -466 -393 -464
rect -401 -468 -398 -466
rect -396 -468 -393 -466
rect -401 -473 -393 -468
rect -401 -475 -398 -473
rect -396 -475 -393 -473
rect -401 -491 -393 -475
rect -391 -482 -383 -464
rect -391 -484 -388 -482
rect -386 -484 -383 -482
rect -391 -491 -383 -484
rect -381 -479 -374 -464
rect -261 -465 -254 -463
rect -261 -467 -259 -465
rect -257 -467 -254 -465
rect -261 -472 -254 -467
rect -261 -474 -259 -472
rect -257 -474 -254 -472
rect -261 -476 -254 -474
rect -381 -481 -378 -479
rect -376 -481 -374 -479
rect -259 -481 -254 -476
rect -252 -470 -246 -463
rect -252 -477 -244 -470
rect -252 -479 -249 -477
rect -247 -479 -244 -477
rect -252 -481 -244 -479
rect -381 -487 -374 -481
rect -250 -483 -244 -481
rect -242 -472 -234 -470
rect -242 -474 -239 -472
rect -237 -474 -234 -472
rect -242 -479 -234 -474
rect -242 -481 -239 -479
rect -237 -481 -234 -479
rect -242 -483 -234 -481
rect -232 -479 -225 -470
rect -232 -481 -229 -479
rect -227 -481 -225 -479
rect -232 -483 -225 -481
rect -381 -489 -378 -487
rect -376 -489 -374 -487
rect -381 -491 -374 -489
<< alu1 >>
rect -292 148 -89 149
rect -45 148 172 149
rect -292 145 172 148
rect -292 144 168 145
rect -292 142 -249 144
rect -247 142 -237 144
rect -235 142 -221 144
rect -219 142 -211 144
rect -209 142 -126 144
rect -124 142 -116 144
rect -114 143 -38 144
rect -114 142 -82 143
rect -292 141 -82 142
rect -80 141 -72 143
rect -70 142 -38 143
rect -36 142 -28 144
rect -26 142 15 144
rect 17 142 25 144
rect 27 142 59 144
rect 61 142 69 144
rect 71 142 102 144
rect 104 142 112 144
rect 114 143 168 144
rect 170 143 172 145
rect 114 142 172 143
rect -70 141 172 142
rect -288 134 -283 136
rect -288 132 -286 134
rect -284 132 -283 134
rect -288 130 -283 132
rect -288 103 -284 130
rect -272 128 -268 136
rect -272 126 -260 128
rect -272 125 -265 126
rect -272 123 -268 125
rect -266 124 -265 125
rect -263 124 -260 126
rect -266 123 -260 124
rect -272 122 -260 123
rect -252 127 -248 136
rect -89 140 -45 141
rect -252 125 -250 127
rect -280 118 -276 120
rect -280 116 -279 118
rect -277 116 -276 118
rect -280 115 -276 116
rect -280 111 -267 115
rect -273 110 -267 111
rect -273 108 -272 110
rect -270 108 -267 110
rect -273 107 -267 108
rect -252 109 -248 125
rect -244 120 -240 128
rect -224 132 -212 136
rect -224 130 -222 132
rect -220 130 -212 132
rect -129 132 -117 136
rect -224 120 -220 130
rect -129 130 -127 132
rect -125 130 -117 132
rect -85 131 -73 135
rect -244 118 -220 120
rect -244 116 -243 118
rect -241 116 -220 118
rect -244 114 -220 116
rect -252 107 -250 109
rect -252 104 -248 107
rect -224 110 -220 114
rect -200 126 -195 128
rect -200 124 -199 126
rect -197 124 -195 126
rect -200 119 -195 124
rect -129 120 -125 130
rect -85 129 -83 131
rect -81 129 -73 131
rect -41 132 -29 135
rect -41 130 -39 132
rect -37 130 -29 132
rect 12 132 24 136
rect -224 108 -219 110
rect -224 106 -222 108
rect -220 106 -219 108
rect -288 102 -275 103
rect -288 100 -283 102
rect -281 100 -275 102
rect -288 99 -275 100
rect -252 103 -240 104
rect -252 102 -243 103
rect -252 100 -250 102
rect -248 101 -243 102
rect -241 101 -240 103
rect -248 100 -240 101
rect -252 98 -240 100
rect -224 101 -219 106
rect -224 99 -222 101
rect -220 99 -219 101
rect -209 118 -195 119
rect -209 116 -205 118
rect -203 116 -195 118
rect -209 115 -195 116
rect -164 118 -125 120
rect -164 116 -155 118
rect -153 116 -125 118
rect -164 114 -125 116
rect -201 110 -188 111
rect -201 108 -195 110
rect -193 108 -188 110
rect -201 107 -188 108
rect -224 97 -219 99
rect -192 101 -188 107
rect -192 99 -191 101
rect -189 99 -188 101
rect -192 98 -188 99
rect -129 110 -125 114
rect -105 126 -100 128
rect -105 124 -103 126
rect -101 124 -100 126
rect -105 119 -100 124
rect -129 108 -124 110
rect -129 106 -127 108
rect -125 106 -124 108
rect -129 101 -124 106
rect -129 99 -127 101
rect -125 99 -124 101
rect -114 118 -100 119
rect -114 116 -110 118
rect -108 116 -100 118
rect -114 115 -100 116
rect -106 110 -93 111
rect -106 108 -100 110
rect -98 108 -96 110
rect -94 108 -93 110
rect -106 107 -93 108
rect -129 97 -124 99
rect -97 98 -93 107
rect -85 109 -81 129
rect -61 126 -56 127
rect -61 124 -59 126
rect -57 124 -56 126
rect -61 118 -56 124
rect -85 107 -80 109
rect -85 105 -83 107
rect -81 105 -80 107
rect -85 103 -80 105
rect -85 101 -84 103
rect -82 101 -80 103
rect -85 100 -80 101
rect -85 98 -83 100
rect -81 98 -80 100
rect -70 117 -56 118
rect -70 115 -66 117
rect -64 115 -56 117
rect -70 114 -56 115
rect -41 112 -37 130
rect 12 130 14 132
rect 16 130 24 132
rect 56 132 68 136
rect -41 110 -40 112
rect -38 110 -37 112
rect -17 127 -12 128
rect -17 125 -16 127
rect -14 125 -12 127
rect -17 119 -12 125
rect -62 109 -49 110
rect -62 107 -56 109
rect -54 107 -49 109
rect -62 106 -49 107
rect -85 96 -80 98
rect -292 84 -89 85
rect -53 100 -49 106
rect -53 98 -52 100
rect -50 98 -49 100
rect -53 97 -49 98
rect -41 108 -36 110
rect -41 106 -39 108
rect -37 106 -36 108
rect -41 101 -36 106
rect -41 99 -39 101
rect -37 99 -36 101
rect -26 118 -12 119
rect -26 116 -22 118
rect -20 116 -12 118
rect -26 115 -12 116
rect 12 114 16 130
rect 56 130 58 132
rect 60 130 68 132
rect 99 132 111 136
rect 12 112 13 114
rect 15 112 16 114
rect -18 110 -5 111
rect -18 108 -12 110
rect -10 108 -8 110
rect -6 108 -5 110
rect -18 107 -5 108
rect -41 97 -36 99
rect -9 98 -5 107
rect 12 110 16 112
rect 36 127 41 128
rect 36 125 37 127
rect 39 125 41 127
rect 36 119 41 125
rect 12 108 17 110
rect 12 106 14 108
rect 16 106 17 108
rect 12 101 17 106
rect 12 99 14 101
rect 16 99 17 101
rect 27 118 41 119
rect 27 116 31 118
rect 33 116 41 118
rect 27 115 41 116
rect 56 112 60 130
rect 99 130 101 132
rect 103 130 111 132
rect 35 110 48 111
rect 35 108 41 110
rect 43 108 48 110
rect 35 107 48 108
rect 12 97 17 99
rect 44 101 48 107
rect 44 99 45 101
rect 47 99 48 101
rect 44 98 48 99
rect 56 110 57 112
rect 59 110 60 112
rect 80 127 85 128
rect 80 125 82 127
rect 84 125 85 127
rect 80 119 85 125
rect 56 108 61 110
rect 56 106 58 108
rect 60 106 61 108
rect 56 101 61 106
rect 56 99 58 101
rect 60 99 61 101
rect 71 118 85 119
rect 71 116 75 118
rect 77 116 85 118
rect 71 115 85 116
rect 79 110 92 111
rect 79 108 80 110
rect 82 108 85 110
rect 87 108 92 110
rect 79 107 92 108
rect 56 97 61 99
rect 88 98 92 107
rect 99 110 103 130
rect 123 127 128 128
rect 123 125 125 127
rect 127 125 128 127
rect 123 119 128 125
rect 99 108 104 110
rect 99 106 101 108
rect 103 106 104 108
rect 99 101 104 106
rect 99 99 101 101
rect 103 99 104 101
rect 114 118 128 119
rect 114 116 118 118
rect 120 116 128 118
rect 114 115 128 116
rect 122 110 135 111
rect 122 108 128 110
rect 130 108 135 110
rect 122 107 135 108
rect 99 97 104 99
rect 131 101 135 107
rect 131 99 132 101
rect 134 99 135 101
rect 131 98 135 99
rect -49 84 139 85
rect -292 82 -273 84
rect -271 82 -265 84
rect -263 82 -249 84
rect -247 82 -237 84
rect -235 82 -221 84
rect -219 82 -126 84
rect -124 83 -38 84
rect -124 82 -82 83
rect -292 81 -82 82
rect -80 82 -38 83
rect -36 82 15 84
rect 17 82 59 84
rect 61 82 102 84
rect 104 82 139 84
rect -80 81 139 82
rect -292 77 139 81
rect -392 75 71 77
rect -392 73 -347 75
rect -345 73 71 75
rect -392 71 -377 73
rect -375 72 71 73
rect -375 71 -269 72
rect -392 70 -269 71
rect -267 70 -138 72
rect -136 70 -6 72
rect -4 70 43 72
rect 45 70 71 72
rect -392 69 71 70
rect 7 63 19 64
rect 7 61 13 63
rect 15 61 19 63
rect -388 54 -372 55
rect -388 52 -376 54
rect -374 52 -372 54
rect -388 51 -372 52
rect -388 23 -384 51
rect -349 52 -336 55
rect -349 50 -347 52
rect -345 50 -343 52
rect -341 50 -336 52
rect -349 49 -336 50
rect -388 21 -387 23
rect -385 22 -364 23
rect -385 21 -368 22
rect -388 20 -368 21
rect -366 20 -364 22
rect -388 19 -364 20
rect -340 32 -336 49
rect -340 30 -339 32
rect -337 30 -336 32
rect -340 28 -336 30
rect -277 51 -264 56
rect -268 47 -264 51
rect -292 38 -279 40
rect -292 37 -283 38
rect -292 35 -291 37
rect -289 36 -283 37
rect -281 36 -279 38
rect -289 35 -279 36
rect -292 34 -279 35
rect -285 27 -279 34
rect -269 45 -264 47
rect -269 43 -268 45
rect -266 43 -264 45
rect -269 41 -264 43
rect -268 37 -264 41
rect -268 35 -267 37
rect -265 35 -264 37
rect -268 34 -264 35
rect -257 54 -241 55
rect -257 52 -245 54
rect -243 52 -241 54
rect -257 51 -241 52
rect -257 23 -253 51
rect -218 52 -205 55
rect -218 50 -216 52
rect -214 50 -212 52
rect -210 50 -205 52
rect -218 49 -205 50
rect -257 22 -233 23
rect -257 20 -245 22
rect -243 20 -237 22
rect -235 20 -233 22
rect -257 19 -233 20
rect -209 32 -205 49
rect -209 30 -208 32
rect -206 30 -205 32
rect -209 28 -205 30
rect -146 51 -133 56
rect -137 47 -133 51
rect -161 39 -148 40
rect -161 37 -153 39
rect -151 37 -148 39
rect -161 35 -160 37
rect -158 35 -148 37
rect -161 34 -148 35
rect -154 27 -148 34
rect -138 45 -133 47
rect -138 43 -137 45
rect -135 43 -133 45
rect -138 41 -133 43
rect -137 38 -133 41
rect -137 36 -136 38
rect -134 36 -133 38
rect -137 34 -133 36
rect -125 54 -109 55
rect -125 52 -113 54
rect -111 52 -109 54
rect -125 51 -109 52
rect -125 23 -121 51
rect 7 58 19 61
rect -86 52 -73 55
rect -86 50 -83 52
rect -81 50 -80 52
rect -78 50 -73 52
rect -86 49 -73 50
rect -125 22 -101 23
rect -125 20 -110 22
rect -108 20 -105 22
rect -103 20 -101 22
rect -125 19 -101 20
rect -77 32 -73 49
rect -77 30 -76 32
rect -74 30 -73 32
rect -77 28 -73 30
rect -14 51 -1 56
rect -5 47 -1 51
rect -29 39 -16 40
rect -29 37 -25 39
rect -23 37 -16 39
rect -29 35 -28 37
rect -26 35 -16 37
rect -29 34 -16 35
rect -22 27 -16 34
rect -6 45 -1 47
rect -6 43 -5 45
rect -3 43 -1 45
rect -6 41 -1 43
rect 7 46 12 58
rect 7 44 9 46
rect 11 44 12 46
rect 7 42 12 44
rect -5 37 -1 41
rect -5 35 -4 37
rect -2 35 -1 37
rect -5 34 -1 35
rect 23 39 28 40
rect 23 37 25 39
rect 27 37 28 39
rect 23 33 28 37
rect 51 55 67 56
rect 51 53 53 55
rect 55 53 67 55
rect 51 51 67 53
rect 23 32 25 33
rect 15 31 25 32
rect 27 31 28 33
rect 15 26 28 31
rect 63 23 67 51
rect 43 22 67 23
rect 43 20 45 22
rect 47 20 67 22
rect 43 19 67 20
rect -392 12 71 13
rect -392 10 -386 12
rect -384 10 -324 12
rect -322 10 -269 12
rect -267 10 -255 12
rect -253 10 -193 12
rect -191 10 -138 12
rect -136 10 -123 12
rect -121 10 -61 12
rect -59 10 -6 12
rect -4 10 10 12
rect 12 10 63 12
rect 65 10 71 12
rect -392 8 71 10
rect -392 6 63 8
rect 65 6 71 8
rect -392 5 71 6
rect -382 1 49 5
rect -382 -1 -375 1
rect -373 -1 -363 1
rect -361 -1 -339 1
rect -337 -1 -281 1
rect -279 -1 -269 1
rect -267 -1 -243 1
rect -241 0 49 1
rect -241 -1 -148 0
rect -382 -2 -148 -1
rect -146 -2 -136 0
rect -134 -2 -111 0
rect -109 -2 12 0
rect 14 -2 22 0
rect 24 -2 49 0
rect -378 -16 -374 -7
rect -284 -8 -280 -7
rect -284 -10 -283 -8
rect -281 -10 -280 -8
rect -378 -18 -376 -16
rect -378 -34 -374 -18
rect -370 -23 -366 -15
rect -336 -16 -317 -15
rect -284 -16 -280 -10
rect -155 -3 49 -2
rect -336 -18 -321 -16
rect -319 -18 -317 -16
rect -336 -20 -317 -18
rect -313 -20 -299 -16
rect -284 -18 -282 -16
rect -370 -24 -358 -23
rect -370 -25 -364 -24
rect -370 -27 -369 -25
rect -367 -26 -364 -25
rect -362 -26 -358 -24
rect -367 -27 -358 -26
rect -370 -29 -358 -27
rect -352 -25 -340 -23
rect -352 -27 -343 -25
rect -341 -27 -340 -25
rect -352 -29 -340 -27
rect -336 -25 -332 -20
rect -313 -24 -309 -20
rect -284 -24 -280 -18
rect -336 -27 -335 -25
rect -333 -27 -332 -25
rect -378 -36 -376 -34
rect -378 -39 -374 -36
rect -352 -34 -348 -29
rect -352 -36 -351 -34
rect -349 -36 -348 -34
rect -336 -32 -332 -27
rect -321 -25 -309 -24
rect -321 -27 -320 -25
rect -318 -27 -317 -25
rect -315 -27 -309 -25
rect -321 -28 -309 -27
rect -305 -25 -280 -24
rect -305 -27 -303 -25
rect -301 -27 -280 -25
rect -305 -29 -280 -27
rect -276 -23 -272 -15
rect -240 -16 -221 -15
rect -240 -18 -239 -16
rect -237 -18 -225 -16
rect -223 -18 -221 -16
rect -240 -20 -221 -18
rect -217 -17 -184 -16
rect -217 -19 -189 -17
rect -187 -19 -184 -17
rect -217 -20 -184 -19
rect -151 -17 -147 -8
rect 9 -12 21 -8
rect -51 -14 11 -12
rect 13 -14 21 -12
rect -151 -19 -149 -17
rect -276 -24 -264 -23
rect -276 -25 -267 -24
rect -276 -27 -275 -25
rect -273 -26 -267 -25
rect -265 -26 -264 -24
rect -273 -27 -264 -26
rect -276 -29 -264 -27
rect -256 -25 -244 -23
rect -256 -27 -255 -25
rect -253 -27 -247 -25
rect -245 -27 -244 -25
rect -256 -29 -244 -27
rect -305 -32 -299 -29
rect -336 -34 -316 -32
rect -336 -36 -320 -34
rect -318 -36 -316 -34
rect -352 -37 -348 -36
rect -405 -41 -366 -39
rect -405 -43 -404 -41
rect -402 -43 -376 -41
rect -374 -43 -366 -41
rect -405 -45 -366 -43
rect -321 -41 -316 -36
rect -321 -43 -320 -41
rect -318 -43 -316 -41
rect -321 -45 -316 -43
rect -312 -37 -299 -32
rect -284 -34 -280 -29
rect -284 -36 -282 -34
rect -312 -45 -308 -37
rect -284 -39 -280 -36
rect -256 -37 -252 -29
rect -240 -32 -236 -20
rect -217 -24 -213 -20
rect -225 -25 -213 -24
rect -225 -27 -221 -25
rect -219 -27 -213 -25
rect -225 -28 -213 -27
rect -209 -25 -203 -24
rect -209 -27 -207 -25
rect -205 -27 -196 -25
rect -209 -29 -200 -27
rect -198 -29 -196 -27
rect -209 -31 -196 -29
rect -151 -27 -147 -19
rect -51 -16 0 -14
rect 2 -16 13 -14
rect -151 -29 -150 -27
rect -148 -29 -147 -27
rect -209 -32 -203 -31
rect -240 -34 -220 -32
rect -240 -36 -224 -34
rect -222 -36 -220 -34
rect -284 -41 -272 -39
rect -284 -43 -282 -41
rect -280 -43 -272 -41
rect -284 -45 -272 -43
rect -225 -41 -220 -36
rect -225 -43 -224 -41
rect -222 -43 -220 -41
rect -225 -45 -220 -43
rect -216 -37 -203 -32
rect -151 -35 -147 -29
rect -143 -24 -139 -16
rect -124 -17 -89 -16
rect -51 -17 13 -16
rect -124 -19 -122 -17
rect -120 -19 -93 -17
rect -91 -19 -89 -17
rect -124 -20 -89 -19
rect -108 -21 -89 -20
rect -85 -18 13 -17
rect -85 -21 -46 -18
rect -143 -25 -131 -24
rect -143 -26 -135 -25
rect -143 -28 -142 -26
rect -140 -27 -135 -26
rect -133 -27 -131 -25
rect -140 -28 -131 -27
rect -143 -30 -131 -28
rect -124 -26 -112 -24
rect -124 -28 -122 -26
rect -120 -28 -115 -26
rect -113 -28 -112 -26
rect -124 -30 -112 -28
rect -151 -37 -149 -35
rect -216 -45 -212 -37
rect -151 -40 -147 -37
rect -124 -38 -120 -30
rect -108 -33 -104 -21
rect -85 -25 -81 -21
rect -93 -26 -81 -25
rect -93 -28 -89 -26
rect -87 -28 -81 -26
rect -93 -29 -81 -28
rect -77 -26 -52 -25
rect -77 -28 -75 -26
rect -73 -27 -52 -26
rect -73 -28 -59 -27
rect -77 -29 -59 -28
rect -57 -29 -52 -27
rect -77 -32 -52 -29
rect -77 -33 -71 -32
rect -108 -35 -88 -33
rect -108 -37 -92 -35
rect -90 -37 -88 -35
rect -151 -42 -139 -40
rect -151 -44 -149 -42
rect -147 -44 -139 -42
rect -151 -46 -139 -44
rect -384 -59 -192 -58
rect -93 -42 -88 -37
rect -93 -44 -92 -42
rect -90 -44 -88 -42
rect -93 -46 -88 -44
rect -84 -38 -71 -33
rect 9 -34 13 -18
rect 33 -25 38 -16
rect 9 -36 14 -34
rect 9 -38 11 -36
rect 13 -38 14 -36
rect -84 -46 -80 -38
rect 9 -43 14 -38
rect 9 -45 11 -43
rect 13 -45 14 -43
rect 24 -26 38 -25
rect 24 -28 25 -26
rect 27 -28 28 -26
rect 30 -28 38 -26
rect 24 -29 38 -28
rect 32 -34 45 -33
rect 32 -36 38 -34
rect 40 -36 42 -34
rect 44 -36 45 -34
rect 32 -37 45 -36
rect 9 -47 14 -45
rect 41 -46 45 -37
rect -384 -61 -375 -59
rect -373 -61 -363 -59
rect -361 -61 -320 -59
rect -318 -61 -281 -59
rect -279 -61 -269 -59
rect -267 -60 49 -59
rect -267 -61 -148 -60
rect -384 -62 -148 -61
rect -146 -62 -136 -60
rect -134 -62 12 -60
rect 14 -62 49 -60
rect -384 -66 49 -62
rect -426 -67 49 -66
rect -426 -68 -75 -67
rect -454 -69 -75 -68
rect -454 -71 -442 -69
rect -440 -71 -75 -69
rect -454 -72 -307 -71
rect -454 -73 -419 -72
rect -454 -75 -447 -73
rect -445 -75 -435 -73
rect -433 -74 -419 -73
rect -417 -73 -307 -72
rect -305 -72 -75 -71
rect -305 -73 -156 -72
rect -417 -74 -156 -73
rect -154 -74 -112 -72
rect -110 -74 -75 -72
rect -433 -75 -314 -74
rect -454 -76 -426 -75
rect -422 -89 -417 -87
rect -450 -91 -438 -89
rect -450 -93 -448 -91
rect -446 -93 -438 -91
rect -450 -95 -438 -93
rect -422 -91 -420 -89
rect -418 -91 -417 -89
rect -310 -88 -305 -86
rect -450 -98 -446 -95
rect -450 -100 -448 -98
rect -510 -106 -467 -105
rect -510 -108 -508 -106
rect -506 -108 -472 -106
rect -470 -108 -467 -106
rect -510 -109 -467 -108
rect -450 -116 -446 -100
rect -422 -96 -417 -91
rect -422 -98 -420 -96
rect -418 -98 -417 -96
rect -422 -100 -417 -98
rect -422 -105 -418 -100
rect -442 -107 -418 -105
rect -442 -109 -441 -107
rect -439 -109 -418 -107
rect -442 -111 -418 -109
rect -450 -118 -448 -116
rect -450 -124 -446 -118
rect -442 -119 -438 -111
rect -450 -126 -449 -124
rect -447 -126 -446 -124
rect -450 -127 -446 -126
rect -422 -120 -418 -111
rect -390 -97 -386 -88
rect -310 -90 -308 -88
rect -306 -90 -305 -88
rect -163 -75 -75 -74
rect -310 -95 -305 -90
rect -310 -97 -308 -95
rect -306 -97 -305 -95
rect -399 -98 -367 -97
rect -399 -100 -393 -98
rect -391 -100 -371 -98
rect -369 -100 -367 -98
rect -399 -101 -367 -100
rect -310 -99 -305 -97
rect -278 -90 -274 -87
rect -278 -92 -277 -90
rect -275 -92 -274 -90
rect -407 -106 -393 -105
rect -407 -108 -403 -106
rect -401 -108 -397 -106
rect -395 -108 -393 -106
rect -407 -109 -393 -108
rect -422 -122 -420 -120
rect -418 -122 -410 -120
rect -422 -126 -410 -122
rect -398 -118 -393 -109
rect -310 -119 -306 -99
rect -278 -96 -274 -92
rect -259 -90 -223 -88
rect -259 -92 -258 -90
rect -256 -92 -229 -90
rect -227 -92 -223 -90
rect -259 -93 -223 -92
rect -159 -89 -154 -87
rect -159 -91 -157 -89
rect -155 -91 -154 -89
rect -287 -97 -274 -96
rect -287 -99 -286 -97
rect -284 -99 -281 -97
rect -279 -99 -274 -97
rect -287 -100 -274 -99
rect -159 -96 -154 -91
rect -159 -98 -157 -96
rect -155 -98 -154 -96
rect -159 -100 -154 -98
rect -127 -90 -123 -88
rect -127 -92 -126 -90
rect -124 -92 -123 -90
rect -295 -105 -281 -104
rect -295 -107 -291 -105
rect -289 -107 -281 -105
rect -295 -108 -281 -107
rect -310 -121 -308 -119
rect -306 -121 -298 -119
rect -310 -123 -305 -121
rect -303 -123 -298 -121
rect -310 -125 -298 -123
rect -286 -113 -281 -108
rect -286 -115 -285 -113
rect -283 -115 -281 -113
rect -286 -117 -281 -115
rect -159 -109 -155 -100
rect -159 -111 -158 -109
rect -156 -111 -155 -109
rect -159 -120 -155 -111
rect -127 -97 -123 -92
rect -136 -98 -123 -97
rect -136 -100 -130 -98
rect -128 -100 -123 -98
rect -136 -101 -123 -100
rect -115 -89 -110 -87
rect -115 -91 -113 -89
rect -111 -91 -110 -89
rect -115 -96 -110 -91
rect -115 -98 -113 -96
rect -111 -98 -110 -96
rect -115 -100 -110 -98
rect -83 -90 -79 -88
rect -83 -92 -82 -90
rect -80 -92 -79 -90
rect -144 -106 -130 -105
rect -144 -108 -140 -106
rect -138 -108 -133 -106
rect -131 -108 -130 -106
rect -144 -109 -130 -108
rect -159 -122 -157 -120
rect -155 -122 -147 -120
rect -159 -126 -147 -122
rect -135 -118 -130 -109
rect -115 -117 -111 -100
rect -83 -97 -79 -92
rect -92 -98 -79 -97
rect -92 -100 -86 -98
rect -84 -100 -79 -98
rect -92 -101 -79 -100
rect -100 -106 -86 -105
rect -100 -108 -96 -106
rect -94 -108 -86 -106
rect -100 -109 -86 -108
rect 129 -106 154 -105
rect 129 -108 130 -106
rect 132 -108 151 -106
rect 153 -108 154 -106
rect 129 -109 154 -108
rect -115 -119 -114 -117
rect -112 -119 -111 -117
rect -115 -120 -111 -119
rect -115 -122 -113 -120
rect -111 -122 -103 -120
rect -115 -126 -103 -122
rect -91 -115 -86 -109
rect -91 -117 -90 -115
rect -88 -117 -86 -115
rect -91 -118 -86 -117
rect -382 -131 -270 -130
rect -426 -132 -307 -131
rect -454 -133 -419 -132
rect -454 -135 -447 -133
rect -445 -135 -435 -133
rect -433 -134 -419 -133
rect -417 -134 -409 -132
rect -407 -133 -307 -132
rect -305 -133 -297 -131
rect -295 -132 -75 -131
rect -295 -133 -156 -132
rect -407 -134 -156 -133
rect -154 -134 -146 -132
rect -144 -134 -112 -132
rect -110 -134 -102 -132
rect -100 -134 -75 -132
rect -433 -135 -75 -134
rect -454 -137 -75 -135
rect -454 -139 -82 -137
rect -80 -139 -75 -137
rect 150 -135 154 -109
rect 150 -137 151 -135
rect 153 -137 154 -135
rect 150 -139 154 -137
rect -454 -140 -77 -139
rect -545 -144 -77 -140
rect -545 -145 -270 -144
rect -545 -147 -539 -145
rect -537 -147 -477 -145
rect -475 -147 -422 -145
rect -420 -147 -407 -145
rect -405 -147 -345 -145
rect -343 -147 -290 -145
rect -288 -146 -270 -145
rect -268 -146 -208 -144
rect -206 -146 -153 -144
rect -151 -146 -139 -144
rect -137 -146 -86 -144
rect -84 -146 -77 -144
rect -288 -147 -77 -146
rect -545 -148 -276 -147
rect -541 -155 -517 -154
rect -541 -157 -521 -155
rect -519 -157 -517 -155
rect -541 -158 -517 -157
rect -541 -185 -537 -158
rect -409 -155 -385 -154
rect -409 -157 -389 -155
rect -387 -157 -385 -155
rect -409 -158 -385 -157
rect -493 -165 -489 -163
rect -493 -167 -492 -165
rect -490 -167 -489 -165
rect -493 -168 -489 -167
rect -493 -170 -492 -168
rect -490 -170 -489 -168
rect -541 -187 -540 -185
rect -538 -186 -537 -185
rect -538 -187 -525 -186
rect -541 -189 -529 -187
rect -527 -189 -525 -187
rect -541 -190 -525 -189
rect -493 -184 -489 -170
rect -502 -185 -489 -184
rect -502 -187 -496 -185
rect -494 -187 -489 -185
rect -502 -190 -489 -187
rect -438 -169 -432 -162
rect -445 -170 -432 -169
rect -445 -172 -444 -170
rect -442 -171 -432 -170
rect -442 -172 -438 -171
rect -445 -173 -438 -172
rect -436 -173 -432 -171
rect -445 -175 -432 -173
rect -421 -176 -417 -169
rect -422 -178 -417 -176
rect -422 -180 -421 -178
rect -419 -180 -417 -178
rect -422 -182 -417 -180
rect -421 -186 -417 -182
rect -430 -187 -417 -186
rect -430 -189 -420 -187
rect -418 -189 -417 -187
rect -430 -191 -417 -189
rect -409 -186 -405 -158
rect -272 -154 -248 -153
rect -272 -156 -252 -154
rect -250 -156 -248 -154
rect -272 -157 -248 -156
rect -361 -165 -357 -163
rect -361 -167 -360 -165
rect -358 -167 -357 -165
rect -361 -170 -357 -167
rect -361 -172 -360 -170
rect -358 -172 -357 -170
rect -409 -187 -393 -186
rect -409 -189 -408 -187
rect -406 -189 -397 -187
rect -395 -189 -393 -187
rect -409 -190 -393 -189
rect -361 -184 -357 -172
rect -370 -185 -357 -184
rect -370 -187 -364 -185
rect -362 -187 -357 -185
rect -370 -190 -357 -187
rect -306 -165 -300 -162
rect -306 -167 -305 -165
rect -303 -167 -300 -165
rect -306 -169 -300 -167
rect -313 -170 -300 -169
rect -313 -172 -312 -170
rect -310 -172 -300 -170
rect -313 -175 -300 -172
rect -289 -176 -285 -169
rect -290 -178 -285 -176
rect -290 -180 -289 -178
rect -287 -180 -285 -178
rect -290 -182 -285 -180
rect -289 -186 -285 -182
rect -298 -188 -285 -186
rect -298 -190 -288 -188
rect -286 -190 -285 -188
rect -272 -185 -268 -157
rect -141 -154 -117 -153
rect -141 -156 -121 -154
rect -119 -156 -117 -154
rect -141 -157 -117 -156
rect -224 -164 -220 -162
rect -224 -166 -223 -164
rect -221 -166 -220 -164
rect -224 -169 -220 -166
rect -224 -171 -223 -169
rect -221 -171 -220 -169
rect -272 -186 -256 -185
rect -272 -188 -271 -186
rect -269 -188 -260 -186
rect -258 -188 -256 -186
rect -272 -189 -256 -188
rect -298 -191 -285 -190
rect -224 -183 -220 -171
rect -233 -184 -220 -183
rect -233 -186 -227 -184
rect -225 -186 -220 -184
rect -233 -189 -220 -186
rect -169 -163 -163 -161
rect -169 -165 -167 -163
rect -165 -165 -163 -163
rect -169 -168 -163 -165
rect -176 -169 -163 -168
rect -176 -171 -175 -169
rect -173 -171 -163 -169
rect -176 -174 -163 -171
rect -152 -175 -148 -168
rect -153 -177 -148 -175
rect -153 -179 -152 -177
rect -150 -179 -148 -177
rect -153 -181 -148 -179
rect -152 -185 -148 -181
rect -161 -186 -148 -185
rect -161 -188 -151 -186
rect -149 -188 -148 -186
rect -161 -190 -148 -188
rect -141 -185 -137 -157
rect -102 -161 -89 -160
rect -102 -163 -100 -161
rect -98 -163 -89 -161
rect -102 -165 -89 -163
rect -102 -167 -101 -165
rect -99 -166 -89 -165
rect -99 -167 -97 -166
rect -141 -187 -125 -185
rect -141 -189 -129 -187
rect -127 -189 -125 -187
rect -141 -190 -125 -189
rect -102 -174 -97 -167
rect -86 -178 -81 -176
rect -86 -180 -85 -178
rect -83 -180 -81 -178
rect -86 -181 -81 -180
rect -86 -183 -84 -181
rect -82 -183 -81 -181
rect -86 -192 -81 -183
rect -93 -198 -81 -192
rect -276 -204 -77 -203
rect -545 -205 -153 -204
rect -545 -207 -422 -205
rect -420 -207 -290 -205
rect -288 -206 -153 -205
rect -151 -206 -119 -204
rect -117 -206 -77 -204
rect -288 -207 -77 -206
rect -545 -208 -77 -207
rect -545 -210 -517 -208
rect -515 -210 -77 -208
rect -545 -211 -77 -210
rect -545 -212 -101 -211
rect -506 -216 -101 -212
rect -506 -217 -233 -216
rect -506 -219 -499 -217
rect -497 -219 -487 -217
rect -485 -219 -406 -217
rect -404 -219 -394 -217
rect -392 -218 -233 -217
rect -231 -218 -221 -216
rect -219 -218 -138 -216
rect -136 -218 -101 -216
rect -392 -219 -318 -218
rect -240 -219 -101 -218
rect -506 -220 -318 -219
rect -502 -235 -490 -233
rect -502 -237 -500 -235
rect -498 -237 -490 -235
rect -502 -239 -490 -237
rect -445 -235 -440 -233
rect -445 -237 -444 -235
rect -442 -237 -440 -235
rect -502 -242 -498 -239
rect -502 -244 -500 -242
rect -502 -250 -498 -244
rect -476 -242 -472 -241
rect -445 -242 -440 -237
rect -476 -244 -475 -242
rect -473 -244 -472 -242
rect -476 -249 -472 -244
rect -460 -244 -444 -242
rect -442 -244 -440 -242
rect -460 -246 -440 -244
rect -436 -236 -432 -233
rect -436 -238 -435 -236
rect -433 -238 -432 -236
rect -436 -241 -432 -238
rect -409 -235 -397 -233
rect -409 -237 -407 -235
rect -405 -237 -404 -235
rect -402 -237 -397 -235
rect -409 -239 -397 -237
rect -272 -229 -268 -226
rect -272 -231 -271 -229
rect -269 -231 -268 -229
rect -351 -235 -346 -233
rect -351 -237 -350 -235
rect -348 -237 -346 -235
rect -436 -246 -423 -241
rect -572 -253 -498 -250
rect -572 -255 -568 -253
rect -566 -255 -498 -253
rect -572 -256 -498 -255
rect -502 -260 -498 -256
rect -494 -251 -482 -249
rect -494 -253 -493 -251
rect -491 -252 -482 -251
rect -491 -253 -485 -252
rect -494 -254 -485 -253
rect -483 -254 -482 -252
rect -494 -255 -482 -254
rect -476 -251 -464 -249
rect -476 -253 -467 -251
rect -465 -253 -464 -251
rect -476 -255 -464 -253
rect -460 -251 -456 -246
rect -460 -253 -459 -251
rect -457 -253 -456 -251
rect -502 -262 -500 -260
rect -502 -271 -498 -262
rect -494 -263 -490 -255
rect -460 -258 -456 -253
rect -445 -251 -433 -250
rect -445 -253 -444 -251
rect -442 -253 -441 -251
rect -439 -253 -433 -251
rect -445 -254 -433 -253
rect -429 -251 -423 -246
rect -429 -253 -427 -251
rect -425 -253 -423 -251
rect -429 -254 -423 -253
rect -409 -242 -405 -239
rect -409 -244 -407 -242
rect -437 -258 -433 -254
rect -460 -260 -441 -258
rect -460 -262 -445 -260
rect -443 -262 -441 -260
rect -437 -262 -423 -258
rect -409 -260 -405 -244
rect -382 -243 -378 -241
rect -351 -242 -346 -237
rect -382 -245 -381 -243
rect -379 -245 -378 -243
rect -382 -249 -378 -245
rect -366 -244 -350 -242
rect -348 -244 -346 -242
rect -366 -246 -346 -244
rect -342 -241 -338 -233
rect -342 -243 -329 -241
rect -342 -245 -333 -243
rect -331 -245 -329 -243
rect -342 -246 -329 -245
rect -401 -251 -389 -249
rect -401 -253 -400 -251
rect -398 -253 -389 -251
rect -401 -255 -389 -253
rect -382 -251 -370 -249
rect -382 -253 -373 -251
rect -371 -253 -370 -251
rect -382 -255 -370 -253
rect -409 -262 -407 -260
rect -460 -263 -441 -262
rect -409 -271 -405 -262
rect -401 -260 -397 -255
rect -401 -262 -400 -260
rect -398 -262 -397 -260
rect -366 -258 -362 -246
rect -351 -251 -339 -250
rect -351 -253 -347 -251
rect -345 -253 -342 -251
rect -340 -253 -339 -251
rect -351 -254 -339 -253
rect -335 -251 -329 -246
rect -335 -253 -333 -251
rect -331 -253 -329 -251
rect -335 -254 -329 -253
rect -343 -258 -339 -254
rect -272 -255 -268 -231
rect -272 -257 -271 -255
rect -269 -257 -268 -255
rect -272 -258 -268 -257
rect -236 -234 -224 -232
rect -236 -236 -234 -234
rect -232 -236 -224 -234
rect -236 -238 -224 -236
rect -177 -234 -172 -232
rect -177 -236 -176 -234
rect -174 -236 -172 -234
rect -236 -241 -232 -238
rect -236 -243 -234 -241
rect -236 -244 -232 -243
rect -236 -246 -235 -244
rect -233 -246 -232 -244
rect -208 -242 -204 -240
rect -177 -241 -172 -236
rect -208 -244 -207 -242
rect -205 -244 -204 -242
rect -366 -260 -347 -258
rect -401 -263 -397 -262
rect -366 -262 -364 -260
rect -362 -262 -351 -260
rect -349 -262 -347 -260
rect -343 -262 -329 -258
rect -236 -259 -232 -246
rect -208 -248 -204 -244
rect -192 -243 -176 -241
rect -174 -243 -172 -241
rect -192 -245 -172 -243
rect -168 -240 -164 -232
rect -141 -233 -136 -231
rect -141 -235 -139 -233
rect -137 -235 -136 -233
rect -141 -236 -136 -235
rect -141 -238 -140 -236
rect -138 -238 -136 -236
rect -141 -240 -136 -238
rect -168 -242 -155 -240
rect -168 -244 -158 -242
rect -156 -244 -155 -242
rect -168 -245 -155 -244
rect -228 -250 -216 -248
rect -228 -252 -227 -250
rect -225 -252 -216 -250
rect -228 -254 -216 -252
rect -208 -250 -196 -248
rect -208 -252 -199 -250
rect -197 -252 -196 -250
rect -208 -254 -196 -252
rect -236 -261 -234 -259
rect -366 -263 -347 -262
rect -236 -270 -232 -261
rect -228 -259 -224 -254
rect -228 -261 -227 -259
rect -225 -261 -224 -259
rect -192 -257 -188 -245
rect -177 -250 -165 -249
rect -177 -252 -173 -250
rect -171 -252 -168 -250
rect -166 -252 -165 -250
rect -177 -253 -165 -252
rect -161 -250 -155 -245
rect -161 -252 -159 -250
rect -157 -252 -155 -250
rect -161 -253 -155 -252
rect -141 -242 -139 -240
rect -137 -242 -136 -240
rect -141 -244 -136 -242
rect -109 -235 -105 -232
rect -109 -237 -108 -235
rect -106 -237 -105 -235
rect -169 -257 -165 -253
rect -192 -259 -173 -257
rect -228 -262 -224 -261
rect -192 -261 -190 -259
rect -188 -261 -177 -259
rect -175 -261 -173 -259
rect -169 -261 -155 -257
rect -192 -262 -173 -261
rect -141 -264 -137 -244
rect -109 -241 -105 -237
rect -118 -242 -105 -241
rect -118 -244 -112 -242
rect -110 -244 -105 -242
rect -118 -245 -105 -244
rect -126 -250 -112 -249
rect -126 -252 -125 -250
rect -123 -252 -122 -250
rect -120 -252 -112 -250
rect -126 -253 -112 -252
rect -322 -274 -240 -273
rect -322 -275 -236 -274
rect -141 -266 -139 -264
rect -137 -266 -129 -264
rect -141 -270 -129 -266
rect -117 -262 -112 -253
rect -322 -276 -101 -275
rect -506 -277 -233 -276
rect -506 -279 -499 -277
rect -497 -279 -487 -277
rect -485 -279 -463 -277
rect -461 -279 -406 -277
rect -404 -279 -394 -277
rect -392 -279 -369 -277
rect -367 -278 -233 -277
rect -231 -278 -221 -276
rect -219 -278 -195 -276
rect -193 -278 -138 -276
rect -136 -278 -128 -276
rect -126 -278 -113 -276
rect -111 -278 -101 -276
rect -367 -279 -318 -278
rect -506 -284 -318 -279
rect -240 -283 -101 -278
rect -582 -289 -349 -284
rect -285 -285 -255 -284
rect -285 -287 -284 -285
rect -282 -287 -259 -285
rect -257 -287 -255 -285
rect -285 -288 -255 -287
rect -582 -291 -575 -289
rect -573 -291 -565 -289
rect -563 -291 -349 -289
rect -239 -291 -203 -283
rect 132 -285 162 -284
rect 132 -287 133 -285
rect 135 -287 159 -285
rect 161 -287 162 -285
rect 132 -288 162 -287
rect -582 -292 -349 -291
rect -288 -297 -254 -296
rect -578 -301 -566 -297
rect -578 -303 -576 -301
rect -574 -303 -566 -301
rect -505 -299 -500 -297
rect -505 -301 -503 -299
rect -501 -301 -500 -299
rect -578 -319 -574 -303
rect -505 -303 -500 -301
rect -578 -321 -577 -319
rect -575 -321 -574 -319
rect -578 -323 -574 -321
rect -554 -307 -549 -305
rect -554 -309 -552 -307
rect -550 -309 -549 -307
rect -554 -314 -549 -309
rect -578 -325 -573 -323
rect -578 -327 -576 -325
rect -574 -327 -573 -325
rect -578 -332 -573 -327
rect -578 -334 -576 -332
rect -574 -334 -573 -332
rect -563 -315 -549 -314
rect -563 -317 -559 -315
rect -557 -317 -549 -315
rect -563 -318 -549 -317
rect -532 -322 -528 -321
rect -555 -323 -531 -322
rect -555 -325 -549 -323
rect -547 -324 -531 -323
rect -529 -324 -528 -322
rect -547 -325 -528 -324
rect -555 -326 -528 -325
rect -578 -336 -573 -334
rect -546 -335 -542 -326
rect -505 -330 -501 -303
rect -489 -305 -485 -297
rect -381 -299 -376 -297
rect -381 -301 -379 -299
rect -377 -301 -376 -299
rect -381 -303 -376 -301
rect -365 -301 -361 -297
rect -288 -299 -286 -297
rect -284 -299 -258 -297
rect -256 -299 -254 -297
rect -288 -300 -254 -299
rect -235 -298 -230 -296
rect -235 -300 -233 -298
rect -231 -300 -230 -298
rect -365 -303 -364 -301
rect -362 -303 -361 -301
rect -489 -306 -477 -305
rect -489 -308 -480 -306
rect -478 -308 -477 -306
rect -489 -310 -485 -308
rect -483 -310 -477 -308
rect -489 -311 -477 -310
rect -497 -315 -493 -313
rect -497 -317 -496 -315
rect -494 -317 -493 -315
rect -497 -318 -493 -317
rect -497 -321 -484 -318
rect -497 -322 -488 -321
rect -490 -323 -488 -322
rect -486 -323 -484 -321
rect -490 -326 -484 -323
rect -505 -331 -492 -330
rect -505 -333 -503 -331
rect -501 -333 -492 -331
rect -505 -334 -492 -333
rect -381 -330 -377 -303
rect -365 -305 -361 -303
rect -235 -302 -230 -300
rect -365 -308 -353 -305
rect -365 -310 -361 -308
rect -359 -310 -353 -308
rect -365 -311 -353 -310
rect -373 -315 -369 -313
rect -373 -317 -372 -315
rect -370 -317 -369 -315
rect -373 -318 -369 -317
rect -287 -318 -245 -317
rect -373 -321 -360 -318
rect -287 -320 -286 -318
rect -284 -320 -248 -318
rect -246 -320 -245 -318
rect -287 -321 -245 -320
rect -373 -322 -363 -321
rect -366 -323 -363 -322
rect -361 -323 -360 -321
rect -366 -326 -360 -323
rect -235 -329 -231 -302
rect -219 -304 -215 -296
rect 133 -297 154 -296
rect 133 -299 134 -297
rect 136 -299 151 -297
rect 153 -299 154 -297
rect 133 -300 154 -299
rect -219 -305 -207 -304
rect -219 -307 -210 -305
rect -208 -307 -207 -305
rect -219 -309 -215 -307
rect -213 -309 -207 -307
rect -219 -310 -207 -309
rect -227 -314 -223 -312
rect -227 -316 -226 -314
rect -224 -316 -223 -314
rect -227 -317 -223 -316
rect -227 -318 -214 -317
rect -227 -320 -225 -318
rect -223 -320 -214 -318
rect -227 -321 -214 -320
rect -220 -325 -214 -321
rect -381 -331 -368 -330
rect -381 -333 -371 -331
rect -369 -333 -368 -331
rect -381 -334 -368 -333
rect -235 -330 -222 -329
rect -235 -332 -234 -330
rect -232 -332 -222 -330
rect -235 -333 -222 -332
rect -239 -348 -203 -347
rect -582 -349 -220 -348
rect -582 -351 -575 -349
rect -573 -351 -490 -349
rect -488 -351 -482 -349
rect -480 -351 -366 -349
rect -364 -351 -358 -349
rect -356 -350 -220 -349
rect -218 -350 -212 -348
rect -210 -350 -203 -348
rect -356 -351 -203 -350
rect -582 -353 -203 -351
rect -582 -355 -197 -353
rect -723 -357 -197 -355
rect -723 -359 -709 -357
rect -707 -358 -197 -357
rect -707 -359 -225 -358
rect -723 -360 -225 -359
rect -223 -360 -197 -358
rect -723 -362 -600 -360
rect -598 -362 -468 -360
rect -466 -362 -336 -360
rect -334 -361 -197 -360
rect -334 -362 -327 -361
rect -723 -363 -327 -362
rect -261 -368 -249 -366
rect -261 -370 -260 -368
rect -258 -370 -249 -368
rect -261 -372 -249 -370
rect -719 -378 -703 -377
rect -719 -380 -707 -378
rect -705 -380 -703 -378
rect -719 -381 -703 -380
rect -719 -409 -715 -381
rect -680 -379 -667 -377
rect -680 -380 -670 -379
rect -680 -382 -674 -380
rect -672 -381 -670 -380
rect -668 -381 -667 -379
rect -672 -382 -667 -381
rect -680 -383 -667 -382
rect -719 -410 -695 -409
rect -719 -412 -699 -410
rect -697 -412 -695 -410
rect -719 -413 -695 -412
rect -671 -400 -667 -383
rect -671 -402 -670 -400
rect -668 -402 -667 -400
rect -671 -404 -667 -402
rect -608 -381 -595 -376
rect -599 -385 -595 -381
rect -623 -394 -610 -392
rect -623 -395 -615 -394
rect -623 -397 -622 -395
rect -620 -396 -615 -395
rect -613 -396 -610 -394
rect -620 -397 -610 -396
rect -623 -398 -610 -397
rect -616 -405 -610 -398
rect -600 -387 -595 -385
rect -600 -389 -599 -387
rect -597 -389 -595 -387
rect -600 -391 -595 -389
rect -599 -395 -595 -391
rect -599 -397 -598 -395
rect -596 -397 -595 -395
rect -599 -398 -595 -397
rect -587 -378 -571 -377
rect -587 -380 -575 -378
rect -573 -380 -571 -378
rect -587 -381 -571 -380
rect -587 -409 -583 -381
rect -548 -380 -535 -377
rect -548 -382 -542 -380
rect -540 -382 -538 -380
rect -536 -382 -535 -380
rect -548 -383 -535 -382
rect -587 -410 -563 -409
rect -587 -412 -567 -410
rect -565 -412 -563 -410
rect -587 -413 -563 -412
rect -539 -400 -535 -383
rect -539 -402 -538 -400
rect -536 -402 -535 -400
rect -539 -404 -535 -402
rect -476 -381 -463 -376
rect -467 -385 -463 -381
rect -491 -394 -478 -392
rect -491 -395 -484 -394
rect -491 -397 -490 -395
rect -488 -396 -484 -395
rect -482 -396 -478 -394
rect -488 -397 -478 -396
rect -491 -398 -478 -397
rect -484 -405 -478 -398
rect -468 -387 -463 -385
rect -468 -389 -467 -387
rect -465 -389 -463 -387
rect -468 -391 -463 -389
rect -467 -394 -463 -391
rect -467 -396 -466 -394
rect -464 -396 -463 -394
rect -467 -398 -463 -396
rect -455 -378 -439 -377
rect -455 -380 -443 -378
rect -441 -380 -439 -378
rect -455 -381 -439 -380
rect -455 -409 -451 -381
rect -416 -378 -403 -377
rect -416 -380 -406 -378
rect -404 -380 -403 -378
rect -416 -382 -410 -380
rect -408 -382 -403 -380
rect -416 -383 -403 -382
rect -455 -410 -431 -409
rect -455 -412 -435 -410
rect -433 -412 -431 -410
rect -455 -413 -431 -412
rect -407 -400 -403 -383
rect -407 -402 -406 -400
rect -404 -402 -403 -400
rect -407 -404 -403 -402
rect -344 -381 -331 -376
rect -335 -385 -331 -381
rect -359 -395 -346 -392
rect -359 -397 -358 -395
rect -356 -397 -355 -395
rect -353 -397 -346 -395
rect -359 -398 -346 -397
rect -352 -405 -346 -398
rect -336 -387 -331 -385
rect -336 -389 -335 -387
rect -333 -389 -331 -387
rect -261 -384 -256 -372
rect -261 -386 -259 -384
rect -257 -386 -256 -384
rect -261 -388 -256 -386
rect -336 -391 -331 -389
rect -335 -395 -331 -391
rect -335 -397 -334 -395
rect -332 -397 -331 -395
rect -335 -398 -331 -397
rect -245 -391 -240 -390
rect -245 -393 -244 -391
rect -242 -393 -240 -391
rect -245 -397 -240 -393
rect -217 -375 -201 -374
rect -217 -377 -215 -375
rect -213 -377 -201 -375
rect -217 -379 -201 -377
rect -245 -398 -243 -397
rect -253 -399 -243 -398
rect -241 -399 -240 -397
rect -253 -404 -240 -399
rect -205 -407 -201 -379
rect -225 -408 -201 -407
rect -225 -410 -223 -408
rect -221 -410 -201 -408
rect -225 -411 -201 -410
rect -265 -418 -197 -417
rect -327 -419 -258 -418
rect -723 -420 -258 -419
rect -256 -420 -205 -418
rect -203 -420 -197 -418
rect -723 -422 -717 -420
rect -715 -422 -655 -420
rect -653 -422 -600 -420
rect -598 -422 -585 -420
rect -583 -422 -523 -420
rect -521 -422 -468 -420
rect -466 -422 -453 -420
rect -451 -422 -391 -420
rect -389 -422 -336 -420
rect -334 -421 -197 -420
rect -334 -422 -208 -421
rect -723 -423 -208 -422
rect -206 -423 -197 -421
rect -723 -425 -197 -423
rect -723 -426 -221 -425
rect -791 -429 -221 -426
rect -791 -431 -258 -429
rect -256 -431 -248 -429
rect -246 -431 -221 -429
rect -791 -433 -785 -431
rect -783 -433 -732 -431
rect -730 -433 -716 -431
rect -714 -433 -704 -431
rect -702 -432 -452 -431
rect -702 -433 -678 -432
rect -791 -434 -678 -433
rect -676 -434 -584 -432
rect -582 -434 -572 -432
rect -570 -434 -546 -432
rect -544 -433 -452 -432
rect -450 -433 -440 -431
rect -438 -433 -417 -431
rect -415 -433 -366 -431
rect -265 -432 -221 -431
rect -544 -434 -366 -433
rect -787 -441 -763 -440
rect -787 -443 -767 -441
rect -765 -443 -763 -441
rect -787 -444 -763 -443
rect -787 -472 -783 -444
rect -749 -452 -735 -447
rect -749 -454 -747 -452
rect -745 -453 -735 -452
rect -745 -454 -743 -453
rect -787 -474 -771 -472
rect -787 -476 -775 -474
rect -773 -476 -771 -474
rect -787 -477 -771 -476
rect -749 -458 -743 -454
rect -749 -460 -747 -458
rect -745 -460 -743 -458
rect -749 -461 -743 -460
rect -719 -448 -715 -439
rect -695 -435 -495 -434
rect -719 -450 -717 -448
rect -749 -470 -745 -466
rect -732 -465 -727 -463
rect -732 -467 -731 -465
rect -729 -467 -727 -465
rect -732 -471 -727 -467
rect -719 -466 -715 -450
rect -587 -442 -583 -440
rect -587 -444 -586 -442
rect -584 -444 -583 -442
rect -711 -455 -707 -447
rect -675 -449 -656 -448
rect -587 -449 -583 -444
rect -675 -451 -660 -449
rect -658 -451 -656 -449
rect -675 -453 -656 -451
rect -652 -450 -638 -449
rect -652 -452 -642 -450
rect -640 -452 -638 -450
rect -652 -453 -638 -452
rect -587 -451 -585 -449
rect -711 -456 -699 -455
rect -711 -457 -702 -456
rect -711 -459 -710 -457
rect -708 -458 -702 -457
rect -700 -458 -699 -456
rect -708 -459 -699 -458
rect -711 -461 -699 -459
rect -691 -458 -679 -456
rect -691 -460 -686 -458
rect -684 -460 -682 -458
rect -680 -460 -679 -458
rect -691 -462 -679 -460
rect -719 -468 -717 -466
rect -719 -471 -715 -468
rect -691 -470 -687 -462
rect -675 -465 -671 -453
rect -652 -457 -648 -453
rect -660 -458 -648 -457
rect -660 -460 -656 -458
rect -654 -460 -648 -458
rect -660 -461 -648 -460
rect -644 -458 -638 -457
rect -644 -460 -642 -458
rect -640 -460 -638 -458
rect -644 -465 -638 -460
rect -675 -467 -655 -465
rect -675 -469 -659 -467
rect -657 -469 -655 -467
rect -660 -471 -655 -469
rect -732 -473 -707 -471
rect -660 -473 -659 -471
rect -657 -473 -655 -471
rect -732 -475 -717 -473
rect -715 -475 -707 -473
rect -732 -477 -707 -475
rect -732 -479 -727 -477
rect -749 -481 -745 -479
rect -747 -483 -745 -481
rect -749 -488 -745 -483
rect -739 -485 -727 -479
rect -747 -490 -745 -488
rect -660 -474 -655 -473
rect -660 -476 -659 -474
rect -657 -476 -655 -474
rect -660 -478 -655 -476
rect -651 -467 -638 -465
rect -651 -469 -642 -467
rect -640 -469 -638 -467
rect -651 -470 -638 -469
rect -587 -467 -583 -451
rect -455 -448 -451 -439
rect -261 -438 -249 -437
rect -261 -440 -259 -438
rect -257 -440 -249 -438
rect -261 -441 -249 -440
rect -261 -443 -259 -441
rect -257 -443 -249 -441
rect -579 -456 -575 -448
rect -543 -449 -524 -448
rect -543 -451 -528 -449
rect -526 -451 -524 -449
rect -543 -453 -524 -451
rect -520 -450 -506 -449
rect -520 -452 -514 -450
rect -512 -452 -506 -450
rect -520 -453 -506 -452
rect -455 -450 -453 -448
rect -579 -458 -567 -456
rect -579 -460 -578 -458
rect -576 -460 -572 -458
rect -570 -460 -567 -458
rect -579 -462 -567 -460
rect -559 -458 -547 -456
rect -559 -460 -554 -458
rect -552 -460 -550 -458
rect -548 -460 -547 -458
rect -559 -462 -547 -460
rect -587 -469 -585 -467
rect -651 -478 -647 -470
rect -587 -472 -583 -469
rect -559 -470 -555 -462
rect -543 -465 -539 -453
rect -520 -457 -516 -453
rect -528 -458 -516 -457
rect -528 -460 -524 -458
rect -522 -460 -516 -458
rect -528 -461 -516 -460
rect -512 -458 -506 -457
rect -512 -460 -510 -458
rect -508 -460 -506 -458
rect -512 -465 -506 -460
rect -543 -466 -523 -465
rect -543 -468 -542 -466
rect -540 -467 -523 -466
rect -540 -468 -527 -467
rect -543 -469 -527 -468
rect -525 -469 -523 -467
rect -587 -474 -575 -472
rect -587 -476 -585 -474
rect -583 -476 -575 -474
rect -587 -478 -575 -476
rect -791 -491 -695 -490
rect -528 -474 -523 -469
rect -528 -476 -527 -474
rect -525 -476 -523 -474
rect -528 -478 -523 -476
rect -519 -470 -506 -465
rect -455 -466 -451 -450
rect -447 -455 -443 -447
rect -414 -448 -395 -447
rect -414 -450 -399 -448
rect -397 -450 -395 -448
rect -414 -452 -395 -450
rect -391 -449 -377 -448
rect -391 -451 -380 -449
rect -378 -451 -377 -449
rect -391 -452 -377 -451
rect -447 -456 -435 -455
rect -447 -457 -439 -456
rect -447 -459 -446 -457
rect -444 -458 -439 -457
rect -437 -458 -435 -456
rect -444 -459 -435 -458
rect -447 -461 -435 -459
rect -430 -457 -418 -455
rect -430 -459 -428 -457
rect -426 -459 -421 -457
rect -419 -459 -418 -457
rect -430 -461 -418 -459
rect -455 -468 -453 -466
rect -519 -473 -515 -470
rect -519 -475 -518 -473
rect -516 -475 -515 -473
rect -519 -478 -515 -475
rect -455 -471 -451 -468
rect -430 -469 -426 -461
rect -414 -464 -410 -452
rect -391 -456 -387 -452
rect -399 -457 -387 -456
rect -399 -459 -395 -457
rect -393 -459 -387 -457
rect -399 -460 -387 -459
rect -383 -457 -377 -456
rect -383 -459 -381 -457
rect -379 -459 -377 -457
rect -383 -464 -377 -459
rect -414 -466 -394 -464
rect -414 -468 -398 -466
rect -396 -468 -394 -466
rect -399 -469 -394 -468
rect -399 -471 -397 -469
rect -395 -471 -394 -469
rect -455 -473 -443 -471
rect -455 -475 -453 -473
rect -451 -475 -450 -473
rect -448 -475 -443 -473
rect -455 -477 -443 -475
rect -399 -473 -394 -471
rect -399 -475 -398 -473
rect -396 -475 -394 -473
rect -399 -477 -394 -475
rect -390 -466 -377 -464
rect -390 -468 -381 -466
rect -379 -468 -377 -466
rect -390 -469 -377 -468
rect -261 -463 -257 -443
rect -237 -448 -232 -445
rect -237 -450 -236 -448
rect -234 -450 -232 -448
rect -237 -454 -232 -450
rect -261 -465 -256 -463
rect -261 -467 -259 -465
rect -257 -467 -256 -465
rect -390 -477 -386 -469
rect -261 -472 -256 -467
rect -261 -474 -259 -472
rect -257 -474 -256 -472
rect -246 -455 -232 -454
rect -246 -457 -242 -455
rect -240 -457 -232 -455
rect -246 -458 -232 -457
rect -238 -463 -225 -462
rect -238 -465 -232 -463
rect -230 -465 -228 -463
rect -226 -465 -225 -463
rect -238 -466 -225 -465
rect -261 -476 -256 -474
rect -229 -475 -225 -466
rect -265 -489 -221 -488
rect -366 -490 -258 -489
rect -459 -491 -258 -490
rect -256 -491 -221 -489
rect -791 -493 -765 -491
rect -763 -493 -716 -491
rect -714 -493 -704 -491
rect -702 -492 -452 -491
rect -702 -493 -584 -492
rect -791 -494 -584 -493
rect -582 -494 -572 -492
rect -570 -493 -452 -492
rect -450 -493 -440 -491
rect -438 -493 -221 -491
rect -570 -494 -221 -493
rect -791 -496 -776 -494
rect -774 -496 -748 -494
rect -746 -496 -221 -494
rect -791 -498 -265 -496
rect -695 -499 -459 -498
<< alu2 >>
rect -61 149 162 153
rect -61 128 -56 149
rect 36 135 154 139
rect 36 128 41 135
rect -305 126 -195 128
rect -305 124 -265 126
rect -263 124 -199 126
rect -197 124 -195 126
rect -305 122 -195 124
rect -105 126 -56 128
rect -105 124 -103 126
rect -101 124 -59 126
rect -57 124 -56 126
rect -17 127 41 128
rect -17 125 -16 127
rect -14 125 37 127
rect 39 125 41 127
rect -17 124 41 125
rect 80 127 146 128
rect 80 125 82 127
rect 84 125 125 127
rect 127 125 146 127
rect -105 123 -56 124
rect 80 123 146 125
rect -392 73 -372 77
rect -392 71 -389 73
rect -387 71 -377 73
rect -375 71 -372 73
rect -392 69 -372 71
rect -349 75 -344 77
rect -349 73 -347 75
rect -345 73 -344 75
rect -349 52 -344 73
rect -349 50 -347 52
rect -345 50 -344 52
rect -349 49 -344 50
rect -305 40 -299 122
rect -160 118 -147 120
rect -160 116 -155 118
rect -153 116 -147 118
rect -273 110 -256 111
rect -273 108 -272 110
rect -270 108 -260 110
rect -258 108 -256 110
rect -273 107 -256 108
rect -285 102 -279 104
rect -285 100 -283 102
rect -281 100 -279 102
rect -285 40 -279 100
rect -244 103 -240 104
rect -244 101 -243 103
rect -241 101 -240 103
rect -244 69 -240 101
rect -192 101 -176 103
rect -192 99 -191 101
rect -189 99 -180 101
rect -178 99 -176 101
rect -192 97 -176 99
rect -244 65 -212 69
rect -351 38 -279 40
rect -218 52 -212 65
rect -218 50 -216 52
rect -214 50 -212 52
rect -351 36 -350 38
rect -348 36 -283 38
rect -281 36 -279 38
rect -351 35 -279 36
rect -388 23 -384 27
rect -388 21 -387 23
rect -385 21 -384 23
rect -493 -41 -399 -39
rect -493 -43 -404 -41
rect -402 -43 -399 -41
rect -493 -45 -399 -43
rect -554 -106 -504 -105
rect -554 -108 -508 -106
rect -506 -108 -504 -106
rect -554 -109 -504 -108
rect -671 -253 -564 -250
rect -671 -255 -568 -253
rect -566 -255 -564 -253
rect -671 -256 -564 -255
rect -723 -357 -704 -355
rect -723 -358 -709 -357
rect -723 -360 -720 -358
rect -718 -359 -709 -358
rect -707 -359 -704 -357
rect -718 -360 -704 -359
rect -723 -363 -704 -360
rect -671 -377 -667 -256
rect -554 -307 -549 -109
rect -493 -168 -489 -45
rect -454 -69 -438 -68
rect -454 -71 -442 -69
rect -440 -71 -438 -69
rect -454 -73 -451 -71
rect -449 -73 -438 -71
rect -454 -75 -438 -73
rect -398 -73 -393 -71
rect -398 -75 -397 -73
rect -395 -75 -393 -73
rect -398 -105 -393 -75
rect -474 -106 -393 -105
rect -474 -108 -472 -106
rect -470 -108 -397 -106
rect -395 -108 -393 -106
rect -474 -109 -393 -108
rect -388 -108 -384 21
rect -365 -24 -332 -23
rect -365 -26 -364 -24
rect -362 -25 -332 -24
rect -362 -26 -335 -25
rect -365 -27 -335 -26
rect -333 -27 -332 -25
rect -365 -29 -332 -27
rect -321 -25 -317 -24
rect -321 -27 -320 -25
rect -318 -27 -317 -25
rect -352 -34 -346 -33
rect -352 -36 -351 -34
rect -349 -36 -346 -34
rect -352 -42 -346 -36
rect -352 -44 -351 -42
rect -349 -44 -346 -42
rect -352 -45 -346 -44
rect -321 -59 -317 -27
rect -321 -61 -320 -59
rect -318 -61 -317 -59
rect -321 -62 -317 -61
rect -305 -71 -299 35
rect -285 34 -279 35
rect -268 37 -264 39
rect -268 35 -267 37
rect -265 35 -264 37
rect -268 -7 -264 35
rect -246 22 -242 23
rect -246 20 -245 22
rect -243 20 -242 22
rect -246 12 -242 20
rect -246 10 -245 12
rect -243 10 -242 12
rect -246 9 -242 10
rect -284 -8 -264 -7
rect -284 -10 -283 -8
rect -281 -10 -264 -8
rect -284 -11 -264 -10
rect -269 -16 -233 -15
rect -269 -18 -239 -16
rect -237 -18 -233 -16
rect -269 -19 -233 -18
rect -269 -24 -261 -19
rect -218 -23 -212 50
rect -160 39 -147 116
rect -25 114 -21 116
rect -41 112 -37 114
rect -97 110 -89 111
rect -97 108 -96 110
rect -94 108 -92 110
rect -90 108 -89 110
rect -97 107 -89 108
rect -41 110 -40 112
rect -38 110 -37 112
rect -41 104 -37 110
rect -25 112 -24 114
rect -22 112 -21 114
rect 12 114 17 116
rect -25 111 -21 112
rect -4 111 3 113
rect -25 110 -3 111
rect -25 108 -8 110
rect -6 109 -3 110
rect -1 109 3 111
rect -6 108 3 109
rect -25 107 3 108
rect 12 112 13 114
rect 15 112 17 114
rect -85 103 -80 104
rect -85 101 -84 103
rect -82 101 -80 103
rect -85 52 -80 101
rect -53 101 -37 104
rect -53 100 -47 101
rect -53 98 -52 100
rect -50 99 -47 100
rect -45 99 -37 101
rect -50 98 -37 99
rect -53 97 -37 98
rect -85 50 -83 52
rect -81 50 -80 52
rect -160 37 -153 39
rect -151 37 -147 39
rect -160 34 -147 37
rect -137 38 -133 41
rect -137 36 -136 38
rect -134 36 -133 38
rect -155 -15 -148 34
rect -137 1 -133 36
rect -111 22 -101 23
rect -111 20 -110 22
rect -108 20 -101 22
rect -111 19 -101 20
rect -106 14 -101 19
rect -106 12 -105 14
rect -103 12 -101 14
rect -106 11 -101 12
rect -137 -1 -136 1
rect -134 -1 -133 1
rect -137 -13 -133 -1
rect -192 -17 -148 -15
rect -192 -19 -189 -17
rect -187 -19 -148 -17
rect -192 -20 -148 -19
rect -129 -17 -117 -16
rect -129 -19 -128 -17
rect -126 -19 -122 -17
rect -120 -19 -117 -17
rect -129 -20 -117 -19
rect -269 -26 -267 -24
rect -265 -26 -261 -24
rect -269 -29 -261 -26
rect -256 -25 -212 -23
rect -85 -24 -80 50
rect -41 40 -37 97
rect 12 64 17 112
rect 23 112 61 113
rect 23 110 57 112
rect 59 110 61 112
rect 23 107 61 110
rect 73 111 83 113
rect 73 109 74 111
rect 76 110 83 111
rect 76 109 80 110
rect 73 108 80 109
rect 82 108 83 110
rect 73 107 83 108
rect 12 63 19 64
rect 12 61 13 63
rect 15 61 19 63
rect 12 60 19 61
rect -41 39 -22 40
rect -41 37 -25 39
rect -23 37 -22 39
rect -41 34 -22 37
rect -5 37 4 38
rect -5 35 -4 37
rect -2 35 4 37
rect -5 34 4 35
rect -41 33 -37 34
rect -137 -25 -128 -24
rect -256 -27 -255 -25
rect -253 -27 -212 -25
rect -256 -29 -212 -27
rect -218 -30 -212 -29
rect -201 -27 -147 -25
rect -201 -29 -200 -27
rect -198 -29 -166 -27
rect -164 -29 -150 -27
rect -148 -29 -147 -27
rect -201 -31 -147 -29
rect -137 -27 -135 -25
rect -133 -27 -131 -25
rect -129 -27 -128 -25
rect -137 -30 -128 -27
rect -124 -26 -80 -24
rect -30 -25 -24 34
rect -1 -14 4 34
rect -1 -16 0 -14
rect 2 -16 4 -14
rect -1 -18 4 -16
rect -124 -28 -122 -26
rect -120 -28 -80 -26
rect -124 -29 -80 -28
rect -65 -27 -24 -25
rect -65 -29 -59 -27
rect -57 -29 -24 -27
rect 15 -25 19 60
rect 23 39 28 107
rect 44 101 135 103
rect 44 99 45 101
rect 47 99 49 101
rect 51 99 132 101
rect 134 99 135 101
rect 44 98 135 99
rect 23 37 25 39
rect 27 37 28 39
rect 23 10 28 37
rect 61 10 71 13
rect 23 5 46 10
rect 61 8 67 10
rect 69 8 71 10
rect 61 6 63 8
rect 65 6 71 8
rect 61 5 71 6
rect 15 -26 28 -25
rect 15 -28 25 -26
rect 27 -28 28 -26
rect 15 -29 28 -28
rect -65 -32 -24 -29
rect 40 -34 46 5
rect 40 -36 42 -34
rect 44 -36 46 -34
rect 40 -37 46 -36
rect -367 -74 -299 -71
rect -367 -76 -365 -74
rect -363 -76 -299 -74
rect -367 -77 -299 -76
rect -246 -69 -242 -64
rect -246 -71 -245 -69
rect -243 -71 -242 -69
rect -278 -90 -253 -88
rect -278 -92 -277 -90
rect -275 -92 -258 -90
rect -256 -92 -253 -90
rect -278 -93 -253 -92
rect -373 -97 -283 -96
rect -373 -98 -286 -97
rect -373 -100 -371 -98
rect -369 -99 -286 -98
rect -284 -99 -283 -97
rect -369 -100 -283 -99
rect -373 -101 -283 -100
rect -388 -112 -357 -108
rect -493 -170 -492 -168
rect -490 -170 -489 -168
rect -554 -309 -552 -307
rect -550 -309 -549 -307
rect -554 -310 -549 -309
rect -541 -185 -537 -176
rect -541 -187 -540 -185
rect -538 -187 -537 -185
rect -687 -379 -667 -377
rect -687 -381 -670 -379
rect -668 -381 -667 -379
rect -687 -383 -667 -381
rect -616 -319 -574 -315
rect -616 -321 -577 -319
rect -575 -321 -574 -319
rect -616 -323 -574 -321
rect -703 -456 -699 -455
rect -749 -458 -744 -456
rect -749 -460 -747 -458
rect -745 -460 -744 -458
rect -791 -494 -769 -490
rect -791 -496 -787 -494
rect -785 -496 -776 -494
rect -774 -496 -769 -494
rect -791 -498 -769 -496
rect -749 -494 -744 -460
rect -703 -458 -702 -456
rect -700 -458 -699 -456
rect -703 -470 -699 -458
rect -687 -458 -683 -383
rect -616 -392 -609 -323
rect -541 -377 -537 -187
rect -527 -208 -511 -204
rect -527 -210 -525 -208
rect -523 -210 -517 -208
rect -515 -210 -511 -208
rect -527 -212 -511 -210
rect -493 -241 -489 -170
rect -450 -124 -446 -123
rect -450 -126 -449 -124
rect -447 -126 -446 -124
rect -450 -169 -446 -126
rect -361 -169 -357 -112
rect -286 -113 -255 -112
rect -286 -115 -285 -113
rect -283 -114 -255 -113
rect -283 -115 -258 -114
rect -286 -116 -258 -115
rect -256 -116 -255 -114
rect -286 -117 -255 -116
rect -306 -121 -302 -119
rect -306 -123 -305 -121
rect -303 -123 -302 -121
rect -306 -164 -302 -123
rect -352 -165 -302 -164
rect -352 -167 -305 -165
rect -303 -167 -302 -165
rect -352 -168 -302 -167
rect -450 -171 -433 -169
rect -450 -173 -438 -171
rect -436 -173 -433 -171
rect -385 -170 -357 -169
rect -385 -172 -360 -170
rect -358 -172 -357 -170
rect -385 -173 -357 -172
rect -450 -175 -433 -173
rect -493 -242 -472 -241
rect -493 -244 -475 -242
rect -473 -244 -472 -242
rect -493 -245 -472 -244
rect -487 -251 -456 -249
rect -487 -252 -459 -251
rect -487 -254 -485 -252
rect -483 -253 -459 -252
rect -457 -253 -456 -251
rect -483 -254 -456 -253
rect -445 -251 -440 -175
rect -421 -187 -417 -184
rect -421 -189 -420 -187
rect -418 -189 -417 -187
rect -421 -233 -417 -189
rect -409 -187 -388 -186
rect -409 -189 -408 -187
rect -406 -189 -388 -187
rect -409 -190 -388 -189
rect -436 -235 -401 -233
rect -436 -236 -404 -235
rect -436 -238 -435 -236
rect -433 -237 -404 -236
rect -402 -237 -401 -235
rect -433 -238 -401 -237
rect -436 -239 -401 -238
rect -445 -253 -444 -251
rect -442 -253 -440 -251
rect -445 -254 -440 -253
rect -487 -255 -456 -254
rect -392 -259 -388 -190
rect -382 -243 -378 -173
rect -382 -245 -381 -243
rect -379 -245 -378 -243
rect -382 -246 -378 -245
rect -343 -251 -339 -168
rect -306 -169 -302 -168
rect -246 -168 -242 -71
rect -232 -90 -79 -88
rect -232 -92 -229 -90
rect -227 -92 -126 -90
rect -124 -92 -82 -90
rect -80 -92 -79 -90
rect -232 -93 -79 -92
rect -135 -106 133 -105
rect -169 -109 -155 -107
rect -135 -108 -133 -106
rect -131 -108 130 -106
rect 132 -108 133 -106
rect -135 -109 133 -108
rect -169 -111 -158 -109
rect -156 -111 -155 -109
rect -169 -114 -155 -111
rect 142 -113 146 123
rect 150 -106 154 135
rect 150 -108 151 -106
rect 153 -108 154 -106
rect 150 -109 154 -108
rect -91 -114 146 -113
rect -169 -163 -163 -114
rect -91 -115 143 -114
rect -169 -165 -167 -163
rect -165 -165 -163 -163
rect -246 -169 -220 -168
rect -246 -171 -223 -169
rect -221 -171 -220 -169
rect -246 -173 -220 -171
rect -289 -188 -285 -185
rect -289 -190 -288 -188
rect -286 -190 -285 -188
rect -289 -240 -285 -190
rect -272 -186 -268 -185
rect -272 -188 -271 -186
rect -269 -188 -268 -186
rect -272 -229 -268 -188
rect -272 -231 -271 -229
rect -269 -231 -268 -229
rect -272 -233 -268 -231
rect -289 -241 -232 -240
rect -335 -243 -232 -241
rect -335 -245 -333 -243
rect -331 -244 -232 -243
rect -331 -245 -235 -244
rect -335 -246 -235 -245
rect -233 -246 -232 -244
rect -224 -241 -220 -173
rect -224 -242 -204 -241
rect -224 -244 -207 -242
rect -205 -244 -204 -242
rect -224 -245 -204 -244
rect -335 -247 -232 -246
rect -343 -253 -342 -251
rect -340 -253 -339 -251
rect -169 -250 -163 -165
rect -125 -117 -111 -116
rect -125 -119 -114 -117
rect -112 -119 -111 -117
rect -91 -117 -90 -115
rect -88 -116 143 -115
rect 145 -116 146 -114
rect -88 -117 146 -116
rect -91 -118 146 -117
rect -125 -120 -111 -119
rect -125 -176 -121 -120
rect 158 -122 162 149
rect 167 146 186 149
rect 167 145 181 146
rect 167 143 168 145
rect 170 144 181 145
rect 183 144 186 146
rect 170 143 186 144
rect 167 141 186 143
rect -21 -123 162 -122
rect -21 -125 -19 -123
rect -17 -125 162 -123
rect -21 -126 162 -125
rect -106 -132 -101 -127
rect -106 -134 -105 -132
rect -103 -134 -101 -132
rect -106 -160 -101 -134
rect -84 -137 -79 -134
rect -84 -139 -82 -137
rect -80 -139 -79 -137
rect -84 -143 -79 -139
rect -84 -145 -82 -143
rect -80 -145 -79 -143
rect -84 -147 -79 -145
rect 142 -137 146 -134
rect 142 -139 143 -137
rect 145 -139 146 -137
rect -106 -161 -62 -160
rect -106 -163 -100 -161
rect -98 -163 -62 -161
rect -106 -164 -62 -163
rect -102 -166 -62 -164
rect -125 -181 -81 -176
rect -125 -183 -84 -181
rect -82 -183 -81 -181
rect -125 -184 -81 -183
rect -152 -186 -148 -184
rect -152 -188 -151 -186
rect -149 -188 -148 -186
rect -152 -234 -148 -188
rect -120 -213 -116 -184
rect -126 -217 -116 -213
rect -152 -236 -136 -234
rect -152 -238 -140 -236
rect -138 -238 -136 -236
rect -152 -239 -136 -238
rect -152 -241 -148 -239
rect -159 -242 -148 -241
rect -159 -244 -158 -242
rect -156 -244 -148 -242
rect -159 -245 -148 -244
rect -169 -252 -168 -250
rect -166 -252 -163 -250
rect -169 -253 -163 -252
rect -126 -250 -121 -217
rect -68 -232 -62 -166
rect -109 -235 -62 -232
rect -109 -237 -108 -235
rect -106 -237 -62 -235
rect -109 -238 -62 -237
rect -126 -252 -125 -250
rect -123 -252 -121 -250
rect -126 -253 -121 -252
rect -343 -254 -339 -253
rect -272 -255 -268 -254
rect -272 -257 -271 -255
rect -269 -257 -268 -255
rect -401 -260 -360 -259
rect -401 -262 -400 -260
rect -398 -262 -364 -260
rect -362 -262 -360 -260
rect -401 -263 -360 -262
rect -481 -285 -400 -284
rect -481 -287 -404 -285
rect -402 -287 -400 -285
rect -481 -288 -400 -287
rect -481 -306 -477 -288
rect -481 -308 -480 -306
rect -478 -308 -477 -306
rect -481 -311 -477 -308
rect -490 -321 -401 -320
rect -532 -322 -488 -321
rect -532 -324 -531 -322
rect -529 -323 -488 -322
rect -486 -323 -405 -321
rect -403 -323 -401 -321
rect -529 -324 -401 -323
rect -532 -325 -401 -324
rect -505 -331 -486 -329
rect -505 -333 -503 -331
rect -501 -333 -486 -331
rect -505 -334 -486 -333
rect -556 -380 -535 -377
rect -556 -382 -538 -380
rect -536 -382 -535 -380
rect -556 -383 -535 -382
rect -644 -394 -609 -392
rect -644 -396 -615 -394
rect -613 -396 -609 -394
rect -644 -398 -609 -396
rect -599 -395 -595 -392
rect -599 -397 -598 -395
rect -596 -397 -595 -395
rect -644 -450 -638 -398
rect -644 -452 -642 -450
rect -640 -452 -638 -450
rect -644 -453 -638 -452
rect -599 -440 -595 -397
rect -599 -442 -583 -440
rect -599 -444 -586 -442
rect -584 -444 -583 -442
rect -599 -445 -583 -444
rect -687 -460 -686 -458
rect -684 -460 -683 -458
rect -687 -462 -683 -460
rect -599 -465 -595 -445
rect -644 -467 -595 -465
rect -644 -469 -642 -467
rect -640 -469 -595 -467
rect -644 -470 -595 -469
rect -573 -458 -569 -456
rect -573 -460 -572 -458
rect -570 -460 -569 -458
rect -703 -471 -655 -470
rect -703 -473 -659 -471
rect -657 -473 -655 -471
rect -703 -474 -655 -473
rect -573 -471 -569 -460
rect -555 -458 -550 -383
rect -491 -392 -486 -334
rect -392 -377 -388 -263
rect -362 -285 -280 -284
rect -362 -287 -360 -285
rect -358 -287 -284 -285
rect -282 -287 -280 -285
rect -362 -288 -280 -287
rect -365 -297 -282 -296
rect -365 -299 -286 -297
rect -284 -299 -282 -297
rect -365 -300 -282 -299
rect -365 -301 -361 -300
rect -365 -303 -364 -301
rect -362 -303 -361 -301
rect -365 -304 -361 -303
rect -365 -318 -282 -317
rect -365 -320 -286 -318
rect -284 -320 -282 -318
rect -381 -321 -282 -320
rect -381 -323 -379 -321
rect -377 -323 -363 -321
rect -361 -323 -360 -321
rect -381 -325 -360 -323
rect -407 -378 -388 -377
rect -407 -380 -406 -378
rect -404 -380 -388 -378
rect -407 -381 -388 -380
rect -515 -394 -479 -392
rect -515 -396 -484 -394
rect -482 -396 -479 -394
rect -515 -398 -479 -396
rect -467 -394 -463 -392
rect -467 -396 -466 -394
rect -464 -396 -463 -394
rect -515 -450 -510 -398
rect -515 -452 -514 -450
rect -512 -452 -510 -450
rect -515 -453 -510 -452
rect -555 -460 -554 -458
rect -552 -460 -550 -458
rect -555 -462 -550 -460
rect -543 -466 -537 -465
rect -543 -468 -542 -466
rect -540 -468 -537 -466
rect -543 -471 -537 -468
rect -467 -471 -463 -396
rect -407 -400 -403 -381
rect -392 -382 -388 -381
rect -372 -331 -368 -330
rect -372 -333 -371 -331
rect -369 -333 -368 -331
rect -372 -392 -368 -333
rect -272 -366 -268 -257
rect -228 -259 -186 -258
rect -228 -261 -227 -259
rect -225 -261 -190 -259
rect -188 -261 -186 -259
rect -228 -262 -186 -261
rect -115 -276 -102 -275
rect -115 -278 -113 -276
rect -111 -278 -106 -276
rect -104 -278 -102 -276
rect -115 -279 -102 -278
rect -260 -285 136 -284
rect -260 -287 -259 -285
rect -257 -287 133 -285
rect 135 -287 136 -285
rect -260 -288 136 -287
rect -261 -297 137 -296
rect -261 -299 -258 -297
rect -256 -299 134 -297
rect 136 -299 137 -297
rect -261 -300 137 -299
rect 142 -304 146 -139
rect 150 -135 154 -132
rect 150 -137 151 -135
rect 153 -137 154 -135
rect 150 -297 154 -137
rect 158 -285 162 -126
rect 158 -287 159 -285
rect 161 -287 162 -285
rect 158 -288 162 -287
rect 150 -299 151 -297
rect 153 -299 154 -297
rect 150 -300 154 -299
rect -212 -305 146 -304
rect -212 -307 -210 -305
rect -208 -307 146 -305
rect -212 -310 146 -307
rect -250 -318 -221 -317
rect -250 -320 -248 -318
rect -246 -320 -225 -318
rect -223 -320 -221 -318
rect -250 -321 -221 -320
rect -245 -330 -231 -329
rect -245 -332 -234 -330
rect -232 -332 -231 -330
rect -245 -333 -231 -332
rect -272 -368 -256 -366
rect -272 -370 -260 -368
rect -258 -370 -256 -368
rect -272 -372 -256 -370
rect -425 -404 -403 -400
rect -381 -395 -352 -392
rect -381 -397 -355 -395
rect -353 -397 -352 -395
rect -381 -398 -352 -397
rect -335 -395 -290 -394
rect -335 -397 -334 -395
rect -332 -397 -290 -395
rect -335 -398 -290 -397
rect -423 -455 -419 -404
rect -381 -449 -377 -398
rect -381 -451 -380 -449
rect -378 -451 -377 -449
rect -381 -452 -377 -451
rect -295 -437 -290 -398
rect -261 -401 -256 -372
rect -245 -390 -240 -333
rect -245 -391 -223 -390
rect -245 -393 -244 -391
rect -242 -393 -223 -391
rect -245 -394 -223 -393
rect -261 -406 -233 -401
rect -295 -438 -255 -437
rect -295 -440 -259 -438
rect -257 -440 -255 -438
rect -295 -442 -255 -440
rect -440 -456 -435 -455
rect -440 -458 -439 -456
rect -437 -458 -435 -456
rect -440 -470 -435 -458
rect -430 -457 -419 -455
rect -430 -459 -428 -457
rect -426 -459 -419 -457
rect -430 -461 -419 -459
rect -295 -461 -290 -442
rect -237 -448 -233 -406
rect -237 -450 -236 -448
rect -234 -450 -233 -448
rect -237 -457 -233 -450
rect -399 -469 -394 -464
rect -383 -466 -290 -461
rect -229 -463 -225 -394
rect -211 -421 -197 -419
rect -211 -423 -208 -421
rect -206 -423 -201 -421
rect -199 -423 -197 -421
rect -211 -425 -197 -423
rect -229 -465 -228 -463
rect -226 -465 -225 -463
rect -229 -466 -225 -465
rect -383 -468 -381 -466
rect -379 -468 -290 -466
rect -383 -469 -290 -468
rect -399 -470 -397 -469
rect -440 -471 -397 -470
rect -395 -471 -394 -469
rect -573 -475 -537 -471
rect -519 -473 -445 -471
rect -519 -475 -518 -473
rect -516 -475 -450 -473
rect -448 -475 -445 -473
rect -440 -475 -394 -471
rect -519 -477 -445 -475
rect -399 -477 -394 -475
rect -749 -496 -748 -494
rect -746 -496 -744 -494
rect -749 -497 -744 -496
<< alu3 >>
rect 179 146 186 149
rect 179 144 181 146
rect 183 144 186 146
rect -93 114 -21 116
rect -93 112 -24 114
rect -22 112 -21 114
rect -93 111 -21 112
rect -4 111 77 113
rect -262 110 -89 111
rect -262 108 -260 110
rect -258 108 -92 110
rect -90 108 -89 110
rect -4 109 -3 111
rect -1 109 74 111
rect 76 109 77 111
rect -4 108 77 109
rect -262 107 -89 108
rect -48 103 52 104
rect -182 101 52 103
rect -182 99 -180 101
rect -178 99 -47 101
rect -45 99 49 101
rect 51 99 52 101
rect -182 97 52 99
rect -454 73 -381 77
rect -454 71 -389 73
rect -387 71 -381 73
rect -454 69 -381 71
rect -454 -67 -445 69
rect -352 38 -346 39
rect -352 36 -350 38
rect -348 36 -346 38
rect -352 -42 -346 36
rect -106 14 -101 16
rect -352 -44 -351 -42
rect -349 -44 -346 -42
rect -352 -45 -346 -44
rect -246 12 -242 13
rect -246 10 -245 12
rect -243 10 -242 12
rect -568 -71 -445 -67
rect -246 -69 -242 10
rect -106 12 -105 14
rect -103 12 -101 14
rect 179 13 186 144
rect -167 1 -133 2
rect -167 -1 -136 1
rect -134 -1 -133 1
rect -167 -2 -133 -1
rect -167 -27 -163 -2
rect -167 -29 -166 -27
rect -164 -29 -163 -27
rect -167 -31 -163 -29
rect -132 -17 -125 -16
rect -132 -19 -128 -17
rect -126 -19 -125 -17
rect -132 -20 -125 -19
rect -132 -25 -128 -20
rect -132 -27 -131 -25
rect -129 -27 -128 -25
rect -132 -30 -128 -27
rect -246 -71 -245 -69
rect -243 -71 -242 -69
rect -568 -73 -451 -71
rect -449 -73 -445 -71
rect -568 -75 -445 -73
rect -399 -73 -361 -71
rect -246 -73 -242 -71
rect -399 -75 -397 -73
rect -395 -74 -361 -73
rect -395 -75 -365 -74
rect -568 -204 -560 -75
rect -399 -76 -365 -75
rect -363 -76 -361 -74
rect -399 -77 -361 -76
rect -259 -114 -255 -112
rect -259 -116 -258 -114
rect -256 -116 -255 -114
rect -259 -122 -255 -116
rect -259 -123 -177 -122
rect -259 -125 -181 -123
rect -179 -125 -177 -123
rect -259 -126 -177 -125
rect -106 -132 -101 12
rect 66 10 186 13
rect 66 8 67 10
rect 69 8 186 10
rect 66 5 186 8
rect 142 -114 146 -112
rect 142 -116 143 -114
rect 145 -116 146 -114
rect -59 -123 -15 -122
rect -59 -125 -57 -123
rect -55 -125 -19 -123
rect -17 -125 -15 -123
rect -59 -126 -15 -125
rect -106 -134 -105 -132
rect -103 -134 -101 -132
rect -106 -135 -101 -134
rect 142 -137 146 -116
rect 142 -139 143 -137
rect 145 -139 146 -137
rect 142 -140 146 -139
rect -84 -143 123 -141
rect -84 -145 -82 -143
rect -80 -145 123 -143
rect -84 -147 123 -145
rect 118 -150 123 -147
rect 179 -150 186 5
rect 118 -156 186 -150
rect -723 -208 -520 -204
rect -723 -210 -525 -208
rect -523 -210 -520 -208
rect -723 -212 -520 -210
rect -723 -355 -714 -212
rect 179 -275 186 -156
rect -108 -276 186 -275
rect -108 -278 -106 -276
rect -104 -278 186 -276
rect -108 -279 186 -278
rect -406 -285 -356 -284
rect -406 -287 -404 -285
rect -402 -287 -360 -285
rect -358 -287 -356 -285
rect -406 -288 -356 -287
rect -406 -321 -375 -320
rect -406 -323 -405 -321
rect -403 -323 -379 -321
rect -377 -323 -375 -321
rect -406 -325 -375 -323
rect -828 -358 -714 -355
rect -828 -360 -720 -358
rect -718 -360 -714 -358
rect -828 -363 -714 -360
rect -828 -491 -819 -363
rect 179 -419 186 -279
rect -204 -421 186 -419
rect -204 -423 -201 -421
rect -199 -423 186 -421
rect -204 -425 186 -423
rect -828 -494 -780 -491
rect -828 -496 -787 -494
rect -785 -496 -780 -494
rect -828 -499 -780 -496
<< alu4 >>
rect -183 -123 -52 -122
rect -183 -125 -181 -123
rect -179 -125 -57 -123
rect -55 -125 -52 -123
rect -183 -126 -52 -125
<< ptie >>
rect -251 144 -233 146
rect -251 142 -249 144
rect -247 142 -237 144
rect -235 142 -233 144
rect -251 140 -233 142
rect -223 144 -217 146
rect -223 142 -221 144
rect -219 142 -217 144
rect -223 140 -217 142
rect -128 144 -122 146
rect -128 142 -126 144
rect -124 142 -122 144
rect -128 140 -122 142
rect -84 143 -78 145
rect -84 141 -82 143
rect -80 141 -78 143
rect -84 139 -78 141
rect -40 144 -34 146
rect -40 142 -38 144
rect -36 142 -34 144
rect -40 140 -34 142
rect 13 144 19 146
rect 13 142 15 144
rect 17 142 19 144
rect 13 140 19 142
rect 57 144 63 146
rect 57 142 59 144
rect 61 142 63 144
rect 57 140 63 142
rect 100 144 106 146
rect 100 142 102 144
rect 104 142 106 144
rect 100 140 106 142
rect -271 12 -265 14
rect -271 10 -269 12
rect -267 10 -265 12
rect -271 8 -265 10
rect -140 12 -134 14
rect -140 10 -138 12
rect -136 10 -134 12
rect -140 8 -134 10
rect -8 12 -2 14
rect -8 10 -6 12
rect -4 10 -2 12
rect -8 8 -2 10
rect 8 12 14 14
rect 8 10 10 12
rect 12 10 14 12
rect 8 8 14 10
rect -377 1 -359 3
rect -377 -1 -375 1
rect -373 -1 -363 1
rect -361 -1 -359 1
rect -377 -3 -359 -1
rect -283 1 -265 3
rect -283 -1 -281 1
rect -279 -1 -269 1
rect -267 -1 -265 1
rect -283 -3 -265 -1
rect -150 0 -132 2
rect -150 -2 -148 0
rect -146 -2 -136 0
rect -134 -2 -132 0
rect -150 -4 -132 -2
rect 10 0 16 2
rect 10 -2 12 0
rect 14 -2 16 0
rect 10 -4 16 -2
rect -449 -133 -431 -131
rect -449 -135 -447 -133
rect -445 -135 -435 -133
rect -433 -135 -431 -133
rect -449 -137 -431 -135
rect -421 -132 -415 -130
rect -421 -134 -419 -132
rect -417 -134 -415 -132
rect -421 -136 -415 -134
rect -309 -131 -303 -129
rect -309 -133 -307 -131
rect -305 -133 -303 -131
rect -309 -135 -303 -133
rect -158 -132 -152 -130
rect -158 -134 -156 -132
rect -154 -134 -152 -132
rect -158 -136 -152 -134
rect -114 -132 -108 -130
rect -114 -134 -112 -132
rect -110 -134 -108 -132
rect -114 -136 -108 -134
rect -424 -145 -418 -143
rect -424 -147 -422 -145
rect -420 -147 -418 -145
rect -424 -149 -418 -147
rect -292 -145 -286 -143
rect -292 -147 -290 -145
rect -288 -147 -286 -145
rect -292 -149 -286 -147
rect -155 -144 -149 -142
rect -155 -146 -153 -144
rect -151 -146 -149 -144
rect -155 -148 -149 -146
rect -88 -144 -82 -142
rect -88 -146 -86 -144
rect -84 -146 -82 -144
rect -88 -148 -82 -146
rect -501 -277 -483 -275
rect -501 -279 -499 -277
rect -497 -279 -487 -277
rect -485 -279 -483 -277
rect -501 -281 -483 -279
rect -408 -277 -390 -275
rect -408 -279 -406 -277
rect -404 -279 -394 -277
rect -392 -279 -390 -277
rect -408 -281 -390 -279
rect -235 -276 -217 -274
rect -235 -278 -233 -276
rect -231 -278 -221 -276
rect -219 -278 -217 -276
rect -235 -280 -217 -278
rect -140 -276 -134 -274
rect -140 -278 -138 -276
rect -136 -278 -134 -276
rect -140 -280 -134 -278
rect -577 -289 -571 -287
rect -577 -291 -575 -289
rect -573 -291 -571 -289
rect -577 -293 -571 -291
rect -602 -420 -596 -418
rect -602 -422 -600 -420
rect -598 -422 -596 -420
rect -602 -424 -596 -422
rect -470 -420 -464 -418
rect -470 -422 -468 -420
rect -466 -422 -464 -420
rect -470 -424 -464 -422
rect -260 -418 -254 -416
rect -338 -420 -332 -418
rect -338 -422 -336 -420
rect -334 -422 -332 -420
rect -260 -420 -258 -418
rect -256 -420 -254 -418
rect -260 -422 -254 -420
rect -338 -424 -332 -422
rect -260 -429 -254 -427
rect -734 -431 -728 -429
rect -734 -433 -732 -431
rect -730 -433 -728 -431
rect -734 -435 -728 -433
rect -718 -431 -700 -429
rect -718 -433 -716 -431
rect -714 -433 -704 -431
rect -702 -433 -700 -431
rect -718 -435 -700 -433
rect -586 -432 -568 -430
rect -586 -434 -584 -432
rect -582 -434 -572 -432
rect -570 -434 -568 -432
rect -586 -436 -568 -434
rect -454 -431 -436 -429
rect -454 -433 -452 -431
rect -450 -433 -440 -431
rect -438 -433 -436 -431
rect -454 -435 -436 -433
rect -260 -431 -258 -429
rect -256 -431 -254 -429
rect -260 -433 -254 -431
<< ntie >>
rect -275 84 -261 86
rect -275 82 -273 84
rect -271 82 -265 84
rect -263 82 -261 84
rect -275 80 -261 82
rect -251 84 -233 86
rect -251 82 -249 84
rect -247 82 -237 84
rect -235 82 -233 84
rect -251 80 -233 82
rect -223 84 -217 86
rect -223 82 -221 84
rect -219 82 -217 84
rect -223 80 -217 82
rect -128 84 -122 86
rect -128 82 -126 84
rect -124 82 -122 84
rect -128 80 -122 82
rect -84 83 -78 85
rect -40 84 -34 86
rect -84 81 -82 83
rect -80 81 -78 83
rect -84 79 -78 81
rect -40 82 -38 84
rect -36 82 -34 84
rect -40 80 -34 82
rect 13 84 19 86
rect 13 82 15 84
rect 17 82 19 84
rect 13 80 19 82
rect 57 84 63 86
rect 57 82 59 84
rect 61 82 63 84
rect 57 80 63 82
rect 100 84 106 86
rect 100 82 102 84
rect 104 82 106 84
rect 100 80 106 82
rect -271 72 -265 74
rect -271 70 -269 72
rect -267 70 -265 72
rect -140 72 -134 74
rect -271 68 -265 70
rect -140 70 -138 72
rect -136 70 -134 72
rect -8 72 -2 74
rect -140 68 -134 70
rect -8 70 -6 72
rect -4 70 -2 72
rect 41 72 47 74
rect -8 68 -2 70
rect 41 70 43 72
rect 45 70 47 72
rect 41 68 47 70
rect -377 -59 -359 -57
rect -283 -59 -265 -57
rect -377 -61 -375 -59
rect -373 -61 -363 -59
rect -361 -61 -359 -59
rect -377 -63 -359 -61
rect -283 -61 -281 -59
rect -279 -61 -269 -59
rect -267 -61 -265 -59
rect -283 -63 -265 -61
rect -150 -60 -132 -58
rect 10 -60 16 -58
rect -150 -62 -148 -60
rect -146 -62 -136 -60
rect -134 -62 -132 -60
rect -150 -64 -132 -62
rect 10 -62 12 -60
rect 14 -62 16 -60
rect 10 -64 16 -62
rect -449 -73 -431 -71
rect -449 -75 -447 -73
rect -445 -75 -435 -73
rect -433 -75 -431 -73
rect -449 -77 -431 -75
rect -421 -72 -415 -70
rect -421 -74 -419 -72
rect -417 -74 -415 -72
rect -421 -76 -415 -74
rect -309 -71 -303 -69
rect -309 -73 -307 -71
rect -305 -73 -303 -71
rect -309 -75 -303 -73
rect -158 -72 -152 -70
rect -158 -74 -156 -72
rect -154 -74 -152 -72
rect -158 -76 -152 -74
rect -114 -72 -108 -70
rect -114 -74 -112 -72
rect -110 -74 -108 -72
rect -114 -76 -108 -74
rect -424 -205 -418 -203
rect -424 -207 -422 -205
rect -420 -207 -418 -205
rect -292 -205 -286 -203
rect -155 -204 -149 -202
rect -424 -209 -418 -207
rect -292 -207 -290 -205
rect -288 -207 -286 -205
rect -292 -209 -286 -207
rect -155 -206 -153 -204
rect -151 -206 -149 -204
rect -121 -204 -115 -202
rect -155 -208 -149 -206
rect -121 -206 -119 -204
rect -117 -206 -115 -204
rect -121 -208 -115 -206
rect -501 -217 -483 -215
rect -501 -219 -499 -217
rect -497 -219 -487 -217
rect -485 -219 -483 -217
rect -408 -217 -390 -215
rect -408 -219 -406 -217
rect -404 -219 -394 -217
rect -392 -219 -390 -217
rect -235 -216 -217 -214
rect -235 -218 -233 -216
rect -231 -218 -221 -216
rect -219 -218 -217 -216
rect -140 -216 -134 -214
rect -140 -218 -138 -216
rect -136 -218 -134 -216
rect -501 -221 -483 -219
rect -408 -221 -390 -219
rect -235 -220 -217 -218
rect -140 -220 -134 -218
rect -577 -349 -571 -347
rect -577 -351 -575 -349
rect -573 -351 -571 -349
rect -577 -353 -571 -351
rect -492 -349 -478 -347
rect -492 -351 -490 -349
rect -488 -351 -482 -349
rect -480 -351 -478 -349
rect -492 -353 -478 -351
rect -368 -349 -354 -347
rect -368 -351 -366 -349
rect -364 -351 -358 -349
rect -356 -351 -354 -349
rect -368 -353 -354 -351
rect -222 -348 -208 -346
rect -222 -350 -220 -348
rect -218 -350 -212 -348
rect -210 -350 -208 -348
rect -222 -352 -208 -350
rect -602 -360 -596 -358
rect -602 -362 -600 -360
rect -598 -362 -596 -360
rect -470 -360 -464 -358
rect -602 -364 -596 -362
rect -470 -362 -468 -360
rect -466 -362 -464 -360
rect -338 -360 -332 -358
rect -227 -358 -221 -356
rect -470 -364 -464 -362
rect -338 -362 -336 -360
rect -334 -362 -332 -360
rect -338 -364 -332 -362
rect -227 -360 -225 -358
rect -223 -360 -221 -358
rect -227 -362 -221 -360
rect -767 -491 -761 -489
rect -767 -493 -765 -491
rect -763 -493 -761 -491
rect -718 -491 -700 -489
rect -767 -495 -761 -493
rect -718 -493 -716 -491
rect -714 -493 -704 -491
rect -702 -493 -700 -491
rect -586 -492 -568 -490
rect -454 -491 -436 -489
rect -260 -489 -254 -487
rect -260 -491 -258 -489
rect -256 -491 -254 -489
rect -718 -495 -700 -493
rect -586 -494 -584 -492
rect -582 -494 -572 -492
rect -570 -494 -568 -492
rect -586 -496 -568 -494
rect -454 -493 -452 -491
rect -450 -493 -440 -491
rect -438 -493 -436 -491
rect -454 -495 -436 -493
rect -260 -493 -254 -491
<< nmos >>
rect -281 130 -279 142
rect -274 130 -272 142
rect -245 123 -243 132
rect -217 125 -215 134
rect -204 125 -202 136
rect -197 125 -195 136
rect -122 125 -120 134
rect -109 125 -107 136
rect -102 125 -100 136
rect -78 124 -76 133
rect -65 124 -63 135
rect -58 124 -56 135
rect -34 125 -32 134
rect -21 125 -19 136
rect -14 125 -12 136
rect 19 125 21 134
rect 32 125 34 136
rect 39 125 41 136
rect 63 125 65 134
rect 76 125 78 136
rect 83 125 85 136
rect 106 125 108 134
rect 119 125 121 136
rect 126 125 128 136
rect -380 12 -378 25
rect -373 12 -371 25
rect -363 12 -361 25
rect -353 17 -351 30
rect -341 14 -339 25
rect -318 12 -316 25
rect -311 12 -309 25
rect -301 12 -299 25
rect -291 17 -289 30
rect -280 20 -278 31
rect -249 12 -247 25
rect -242 12 -240 25
rect -232 12 -230 25
rect -222 17 -220 30
rect -210 14 -208 25
rect -187 12 -185 25
rect -180 12 -178 25
rect -170 12 -168 25
rect -160 17 -158 30
rect -149 20 -147 31
rect -117 12 -115 25
rect -110 12 -108 25
rect -100 12 -98 25
rect -90 17 -88 30
rect -78 14 -76 25
rect -55 12 -53 25
rect -48 12 -46 25
rect -38 12 -36 25
rect -28 17 -26 30
rect -17 20 -15 31
rect 14 22 16 31
rect 30 17 32 26
rect 40 17 42 26
rect 50 14 52 26
rect 57 14 59 26
rect -371 -20 -369 -11
rect -345 -18 -343 -6
rect -333 -20 -331 -8
rect -326 -20 -324 -8
rect -316 -20 -314 -8
rect -306 -20 -304 -8
rect -277 -20 -275 -11
rect -249 -18 -247 -6
rect -237 -20 -235 -8
rect -230 -20 -228 -8
rect -220 -20 -218 -8
rect -210 -20 -208 -8
rect -144 -21 -142 -12
rect -117 -19 -115 -7
rect -105 -21 -103 -9
rect -98 -21 -96 -9
rect -88 -21 -86 -9
rect -78 -21 -76 -9
rect 16 -19 18 -10
rect 29 -19 31 -8
rect 36 -19 38 -8
rect -443 -123 -441 -114
rect -415 -124 -413 -115
rect -402 -126 -400 -115
rect -395 -126 -393 -115
rect -303 -123 -301 -114
rect -290 -125 -288 -114
rect -283 -125 -281 -114
rect -152 -124 -150 -115
rect -139 -126 -137 -115
rect -132 -126 -130 -115
rect -108 -124 -106 -115
rect -95 -126 -93 -115
rect -88 -126 -86 -115
rect -533 -160 -531 -147
rect -526 -160 -524 -147
rect -516 -160 -514 -147
rect -506 -165 -504 -152
rect -494 -160 -492 -149
rect -471 -160 -469 -147
rect -464 -160 -462 -147
rect -454 -160 -452 -147
rect -444 -165 -442 -152
rect -433 -166 -431 -155
rect -401 -160 -399 -147
rect -394 -160 -392 -147
rect -384 -160 -382 -147
rect -374 -165 -372 -152
rect -362 -160 -360 -149
rect -339 -160 -337 -147
rect -332 -160 -330 -147
rect -322 -160 -320 -147
rect -312 -165 -310 -152
rect -301 -166 -299 -155
rect -264 -159 -262 -146
rect -257 -159 -255 -146
rect -247 -159 -245 -146
rect -237 -164 -235 -151
rect -225 -159 -223 -148
rect -202 -159 -200 -146
rect -195 -159 -193 -146
rect -185 -159 -183 -146
rect -175 -164 -173 -151
rect -164 -165 -162 -154
rect -133 -160 -131 -148
rect -126 -160 -124 -148
rect -116 -160 -114 -151
rect -106 -160 -104 -151
rect -90 -165 -88 -156
rect -495 -267 -493 -258
rect -469 -272 -467 -260
rect -457 -270 -455 -258
rect -450 -270 -448 -258
rect -440 -270 -438 -258
rect -430 -270 -428 -258
rect -402 -267 -400 -258
rect -375 -272 -373 -260
rect -363 -270 -361 -258
rect -356 -270 -354 -258
rect -346 -270 -344 -258
rect -336 -270 -334 -258
rect -229 -266 -227 -257
rect -201 -271 -199 -259
rect -189 -269 -187 -257
rect -182 -269 -180 -257
rect -172 -269 -170 -257
rect -162 -269 -160 -257
rect -134 -268 -132 -259
rect -121 -270 -119 -259
rect -114 -270 -112 -259
rect -571 -308 -569 -299
rect -558 -308 -556 -297
rect -551 -308 -549 -297
rect -498 -303 -496 -291
rect -491 -303 -489 -291
rect -374 -303 -372 -291
rect -367 -303 -365 -291
rect -228 -302 -226 -290
rect -221 -302 -219 -290
rect -711 -420 -709 -407
rect -704 -420 -702 -407
rect -694 -420 -692 -407
rect -684 -415 -682 -402
rect -672 -418 -670 -407
rect -649 -420 -647 -407
rect -642 -420 -640 -407
rect -632 -420 -630 -407
rect -622 -415 -620 -402
rect -611 -412 -609 -401
rect -579 -420 -577 -407
rect -572 -420 -570 -407
rect -562 -420 -560 -407
rect -552 -415 -550 -402
rect -540 -418 -538 -407
rect -517 -420 -515 -407
rect -510 -420 -508 -407
rect -500 -420 -498 -407
rect -490 -415 -488 -402
rect -479 -412 -477 -401
rect -447 -420 -445 -407
rect -440 -420 -438 -407
rect -430 -420 -428 -407
rect -420 -415 -418 -402
rect -408 -418 -406 -407
rect -385 -420 -383 -407
rect -378 -420 -376 -407
rect -368 -420 -366 -407
rect -358 -415 -356 -402
rect -347 -412 -345 -401
rect -254 -408 -252 -399
rect -238 -413 -236 -404
rect -228 -413 -226 -404
rect -218 -416 -216 -404
rect -211 -416 -209 -404
rect -779 -447 -777 -435
rect -772 -447 -770 -435
rect -762 -447 -760 -438
rect -752 -447 -750 -438
rect -736 -452 -734 -443
rect -712 -452 -710 -443
rect -684 -451 -682 -439
rect -672 -453 -670 -441
rect -665 -453 -663 -441
rect -655 -453 -653 -441
rect -645 -453 -643 -441
rect -580 -453 -578 -444
rect -552 -451 -550 -439
rect -540 -453 -538 -441
rect -533 -453 -531 -441
rect -523 -453 -521 -441
rect -513 -453 -511 -441
rect -448 -452 -446 -443
rect -423 -450 -421 -438
rect -411 -452 -409 -440
rect -404 -452 -402 -440
rect -394 -452 -392 -440
rect -384 -452 -382 -440
rect -254 -448 -252 -439
rect -241 -448 -239 -437
rect -234 -448 -232 -437
<< pmos >>
rect -280 92 -278 106
rect -270 92 -268 106
rect -245 93 -243 111
rect -217 92 -215 110
rect -207 90 -205 103
rect -197 90 -195 103
rect -122 92 -120 110
rect -112 90 -110 103
rect -102 90 -100 103
rect -78 91 -76 109
rect -68 89 -66 102
rect -58 89 -56 102
rect -34 92 -32 110
rect -24 90 -22 103
rect -14 90 -12 103
rect 19 92 21 110
rect 29 90 31 103
rect 39 90 41 103
rect 63 92 65 110
rect 73 90 75 103
rect 83 90 85 103
rect 106 92 108 110
rect 116 90 118 103
rect 126 90 128 103
rect -381 43 -379 71
rect -371 43 -369 71
rect -361 43 -359 71
rect -351 57 -349 71
rect -341 57 -339 71
rect -321 43 -319 71
rect -311 43 -309 71
rect -301 43 -299 71
rect -290 50 -288 64
rect -280 50 -278 64
rect -250 43 -248 71
rect -240 43 -238 71
rect -230 43 -228 71
rect -220 57 -218 71
rect -210 57 -208 71
rect -190 43 -188 71
rect -180 43 -178 71
rect -170 43 -168 71
rect -159 50 -157 64
rect -149 50 -147 64
rect -118 43 -116 71
rect -108 43 -106 71
rect -98 43 -96 71
rect -88 57 -86 71
rect -78 57 -76 71
rect -58 43 -56 71
rect -48 43 -46 71
rect -38 43 -36 71
rect -27 50 -25 64
rect -17 50 -15 64
rect 22 44 24 71
rect 38 44 40 62
rect 48 44 50 62
rect 58 44 60 71
rect -371 -50 -369 -32
rect -342 -59 -340 -32
rect -332 -59 -330 -32
rect -325 -59 -323 -32
rect -315 -59 -313 -32
rect -305 -59 -303 -32
rect -277 -50 -275 -32
rect -246 -59 -244 -32
rect -236 -59 -234 -32
rect -229 -59 -227 -32
rect -219 -59 -217 -32
rect -209 -59 -207 -32
rect -144 -51 -142 -33
rect -114 -60 -112 -33
rect -104 -60 -102 -33
rect -97 -60 -95 -33
rect -87 -60 -85 -33
rect -77 -60 -75 -33
rect 16 -52 18 -34
rect 26 -54 28 -41
rect 36 -54 38 -41
rect -443 -102 -441 -84
rect -415 -100 -413 -82
rect -405 -93 -403 -80
rect -395 -93 -393 -80
rect -303 -99 -301 -81
rect -293 -92 -291 -79
rect -283 -92 -281 -79
rect -152 -100 -150 -82
rect -142 -93 -140 -80
rect -132 -93 -130 -80
rect -108 -100 -106 -82
rect -98 -93 -96 -80
rect -88 -93 -86 -80
rect -534 -206 -532 -178
rect -524 -206 -522 -178
rect -514 -206 -512 -178
rect -504 -206 -502 -192
rect -494 -206 -492 -192
rect -474 -206 -472 -178
rect -464 -206 -462 -178
rect -454 -206 -452 -178
rect -443 -199 -441 -185
rect -433 -199 -431 -185
rect -402 -206 -400 -178
rect -392 -206 -390 -178
rect -382 -206 -380 -178
rect -372 -206 -370 -192
rect -362 -206 -360 -192
rect -342 -206 -340 -178
rect -332 -206 -330 -178
rect -322 -206 -320 -178
rect -311 -199 -309 -185
rect -301 -199 -299 -185
rect -265 -205 -263 -177
rect -255 -205 -253 -177
rect -245 -205 -243 -177
rect -235 -205 -233 -191
rect -225 -205 -223 -191
rect -205 -205 -203 -177
rect -195 -205 -193 -177
rect -185 -205 -183 -177
rect -174 -198 -172 -184
rect -164 -198 -162 -184
rect -134 -205 -132 -178
rect -124 -196 -122 -178
rect -114 -196 -112 -178
rect -98 -205 -96 -178
rect -495 -246 -493 -228
rect -466 -246 -464 -219
rect -456 -246 -454 -219
rect -449 -246 -447 -219
rect -439 -246 -437 -219
rect -429 -246 -427 -219
rect -402 -246 -400 -228
rect -372 -246 -370 -219
rect -362 -246 -360 -219
rect -355 -246 -353 -219
rect -345 -246 -343 -219
rect -335 -246 -333 -219
rect -229 -245 -227 -227
rect -198 -245 -196 -218
rect -188 -245 -186 -218
rect -181 -245 -179 -218
rect -171 -245 -169 -218
rect -161 -245 -159 -218
rect -134 -244 -132 -226
rect -124 -237 -122 -224
rect -114 -237 -112 -224
rect -571 -341 -569 -323
rect -561 -343 -559 -330
rect -551 -343 -549 -330
rect -497 -341 -495 -327
rect -487 -341 -485 -327
rect -373 -341 -371 -327
rect -363 -341 -361 -327
rect -227 -340 -225 -326
rect -217 -340 -215 -326
rect -712 -389 -710 -361
rect -702 -389 -700 -361
rect -692 -389 -690 -361
rect -682 -375 -680 -361
rect -672 -375 -670 -361
rect -652 -389 -650 -361
rect -642 -389 -640 -361
rect -632 -389 -630 -361
rect -621 -382 -619 -368
rect -611 -382 -609 -368
rect -580 -389 -578 -361
rect -570 -389 -568 -361
rect -560 -389 -558 -361
rect -550 -375 -548 -361
rect -540 -375 -538 -361
rect -520 -389 -518 -361
rect -510 -389 -508 -361
rect -500 -389 -498 -361
rect -489 -382 -487 -368
rect -479 -382 -477 -368
rect -448 -389 -446 -361
rect -438 -389 -436 -361
rect -428 -389 -426 -361
rect -418 -375 -416 -361
rect -408 -375 -406 -361
rect -388 -389 -386 -361
rect -378 -389 -376 -361
rect -368 -389 -366 -361
rect -357 -382 -355 -368
rect -347 -382 -345 -368
rect -246 -386 -244 -359
rect -230 -386 -228 -368
rect -220 -386 -218 -368
rect -210 -386 -208 -359
rect -780 -492 -778 -465
rect -770 -483 -768 -465
rect -760 -483 -758 -465
rect -744 -492 -742 -465
rect -712 -482 -710 -464
rect -681 -492 -679 -465
rect -671 -492 -669 -465
rect -664 -492 -662 -465
rect -654 -492 -652 -465
rect -644 -492 -642 -465
rect -580 -483 -578 -465
rect -549 -492 -547 -465
rect -539 -492 -537 -465
rect -532 -492 -530 -465
rect -522 -492 -520 -465
rect -512 -492 -510 -465
rect -448 -482 -446 -464
rect -420 -491 -418 -464
rect -410 -491 -408 -464
rect -403 -491 -401 -464
rect -393 -491 -391 -464
rect -383 -491 -381 -464
rect -254 -481 -252 -463
rect -244 -483 -242 -470
rect -234 -483 -232 -470
<< polyct0 >>
rect -215 116 -213 118
rect -120 116 -118 118
rect -76 115 -74 117
rect -32 116 -30 118
rect 21 116 23 118
rect 65 116 67 118
rect 108 116 110 118
rect -379 36 -377 38
rect -369 36 -367 38
rect -329 36 -327 38
rect -319 36 -317 38
rect -309 36 -307 38
rect -248 36 -246 38
rect -238 36 -236 38
rect -198 36 -196 38
rect -188 36 -186 38
rect -178 36 -176 38
rect -116 36 -114 38
rect -106 36 -104 38
rect -66 36 -64 38
rect -56 36 -54 38
rect -46 36 -44 38
rect 46 36 48 38
rect 56 37 58 39
rect 18 -28 20 -26
rect -413 -108 -411 -106
rect -301 -107 -299 -105
rect -150 -108 -148 -106
rect -106 -108 -104 -106
rect -532 -173 -530 -171
rect -522 -173 -520 -171
rect -482 -173 -480 -171
rect -472 -173 -470 -171
rect -462 -173 -460 -171
rect -400 -173 -398 -171
rect -390 -173 -388 -171
rect -350 -173 -348 -171
rect -340 -173 -338 -171
rect -330 -173 -328 -171
rect -263 -172 -261 -170
rect -253 -172 -251 -170
rect -213 -172 -211 -170
rect -203 -172 -201 -170
rect -193 -172 -191 -170
rect -132 -173 -130 -171
rect -122 -172 -120 -170
rect -132 -252 -130 -250
rect -569 -317 -567 -315
rect -710 -396 -708 -394
rect -700 -396 -698 -394
rect -660 -396 -658 -394
rect -650 -396 -648 -394
rect -640 -396 -638 -394
rect -578 -396 -576 -394
rect -568 -396 -566 -394
rect -528 -396 -526 -394
rect -518 -396 -516 -394
rect -508 -396 -506 -394
rect -446 -396 -444 -394
rect -436 -396 -434 -394
rect -396 -396 -394 -394
rect -386 -396 -384 -394
rect -376 -396 -374 -394
rect -222 -394 -220 -392
rect -212 -393 -210 -391
rect -778 -460 -776 -458
rect -768 -459 -766 -457
rect -252 -457 -250 -455
<< polyct1 >>
rect -268 123 -266 125
rect -279 116 -277 118
rect -243 116 -241 118
rect -205 116 -203 118
rect -110 116 -108 118
rect -195 108 -193 110
rect -66 115 -64 117
rect -100 108 -98 110
rect -22 116 -20 118
rect -56 107 -54 109
rect 31 116 33 118
rect -12 108 -10 110
rect 75 116 77 118
rect 41 108 43 110
rect 118 116 120 118
rect 85 108 87 110
rect 128 108 130 110
rect -343 50 -341 52
rect -291 35 -289 37
rect -339 30 -337 32
rect -268 43 -266 45
rect -212 50 -210 52
rect -160 35 -158 37
rect -208 30 -206 32
rect -137 43 -135 45
rect -80 50 -78 52
rect -28 35 -26 37
rect -76 30 -74 32
rect -5 43 -3 45
rect 9 44 11 46
rect 25 31 27 33
rect -369 -27 -367 -25
rect -343 -27 -341 -25
rect -317 -27 -315 -25
rect -303 -27 -301 -25
rect -275 -27 -273 -25
rect -247 -27 -245 -25
rect -221 -27 -219 -25
rect -207 -27 -205 -25
rect -142 -28 -140 -26
rect -115 -28 -113 -26
rect -89 -28 -87 -26
rect -75 -28 -73 -26
rect 28 -28 30 -26
rect 38 -36 40 -34
rect -393 -100 -391 -98
rect -441 -109 -439 -107
rect -403 -108 -401 -106
rect -281 -99 -279 -97
rect -291 -107 -289 -105
rect -130 -100 -128 -98
rect -140 -108 -138 -106
rect -86 -100 -84 -98
rect -96 -108 -94 -106
rect -492 -167 -490 -165
rect -444 -172 -442 -170
rect -496 -187 -494 -185
rect -360 -167 -358 -165
rect -312 -172 -310 -170
rect -421 -180 -419 -178
rect -364 -187 -362 -185
rect -223 -166 -221 -164
rect -175 -171 -173 -169
rect -289 -180 -287 -178
rect -227 -186 -225 -184
rect -101 -167 -99 -165
rect -152 -179 -150 -177
rect -85 -180 -83 -178
rect -493 -253 -491 -251
rect -467 -253 -465 -251
rect -441 -253 -439 -251
rect -427 -253 -425 -251
rect -400 -253 -398 -251
rect -373 -253 -371 -251
rect -347 -253 -345 -251
rect -333 -253 -331 -251
rect -227 -252 -225 -250
rect -199 -252 -197 -250
rect -112 -244 -110 -242
rect -173 -252 -171 -250
rect -159 -252 -157 -250
rect -122 -252 -120 -250
rect -559 -317 -557 -315
rect -485 -310 -483 -308
rect -496 -317 -494 -315
rect -549 -325 -547 -323
rect -361 -310 -359 -308
rect -215 -309 -213 -307
rect -372 -317 -370 -315
rect -226 -316 -224 -314
rect -674 -382 -672 -380
rect -622 -397 -620 -395
rect -670 -402 -668 -400
rect -599 -389 -597 -387
rect -542 -382 -540 -380
rect -490 -397 -488 -395
rect -538 -402 -536 -400
rect -467 -389 -465 -387
rect -410 -382 -408 -380
rect -358 -397 -356 -395
rect -406 -402 -404 -400
rect -335 -389 -333 -387
rect -259 -386 -257 -384
rect -243 -399 -241 -397
rect -747 -454 -745 -452
rect -710 -459 -708 -457
rect -682 -460 -680 -458
rect -731 -467 -729 -465
rect -656 -460 -654 -458
rect -642 -460 -640 -458
rect -578 -460 -576 -458
rect -550 -460 -548 -458
rect -524 -460 -522 -458
rect -510 -460 -508 -458
rect -446 -459 -444 -457
rect -421 -459 -419 -457
rect -395 -459 -393 -457
rect -381 -459 -379 -457
rect -242 -457 -240 -455
rect -232 -465 -230 -463
<< ndifct0 >>
rect -264 138 -262 140
rect -236 128 -234 130
rect -192 132 -190 134
rect -97 132 -95 134
rect -53 131 -51 133
rect -9 132 -7 134
rect 44 132 46 134
rect 88 132 90 134
rect 131 132 133 134
rect -358 21 -356 23
rect -347 13 -345 15
rect -336 21 -334 23
rect -306 20 -304 22
rect -296 21 -294 23
rect -286 19 -284 21
rect -275 27 -273 29
rect -227 21 -225 23
rect -216 13 -214 15
rect -205 21 -203 23
rect -175 20 -173 22
rect -165 21 -163 23
rect -155 19 -153 21
rect -144 27 -142 29
rect -95 21 -93 23
rect -84 13 -82 15
rect -73 21 -71 23
rect -43 20 -41 22
rect -33 21 -31 23
rect -23 19 -21 21
rect -12 27 -10 29
rect 9 27 11 29
rect 23 19 25 21
rect 35 22 37 24
rect -350 -10 -348 -8
rect -362 -15 -360 -13
rect -311 -12 -309 -10
rect -301 -12 -299 -10
rect -254 -10 -252 -8
rect -268 -15 -266 -13
rect -215 -12 -213 -10
rect -205 -12 -203 -10
rect -122 -11 -120 -9
rect -135 -16 -133 -14
rect -83 -13 -81 -11
rect -73 -13 -71 -11
rect 41 -12 43 -10
rect -434 -121 -432 -119
rect -390 -124 -388 -122
rect -278 -123 -276 -121
rect -127 -124 -125 -122
rect -83 -124 -81 -122
rect -500 -150 -498 -148
rect -511 -158 -509 -156
rect -489 -158 -487 -156
rect -459 -157 -457 -155
rect -449 -158 -447 -156
rect -439 -156 -437 -154
rect -368 -150 -366 -148
rect -379 -158 -377 -156
rect -428 -164 -426 -162
rect -357 -158 -355 -156
rect -327 -157 -325 -155
rect -317 -158 -315 -156
rect -307 -156 -305 -154
rect -231 -149 -229 -147
rect -242 -157 -240 -155
rect -296 -164 -294 -162
rect -220 -157 -218 -155
rect -190 -156 -188 -154
rect -180 -157 -178 -155
rect -170 -155 -168 -153
rect -111 -158 -109 -156
rect -99 -155 -97 -153
rect -159 -163 -157 -161
rect -85 -163 -83 -161
rect -486 -265 -484 -263
rect -474 -270 -472 -268
rect -435 -268 -433 -266
rect -425 -268 -423 -266
rect -393 -265 -391 -263
rect -380 -270 -378 -268
rect -341 -268 -339 -266
rect -220 -264 -218 -262
rect -331 -268 -329 -266
rect -206 -269 -204 -267
rect -167 -267 -165 -265
rect -157 -267 -155 -265
rect -109 -268 -107 -266
rect -546 -301 -544 -299
rect -481 -295 -479 -293
rect -357 -295 -355 -293
rect -211 -294 -209 -292
rect -689 -411 -687 -409
rect -678 -419 -676 -417
rect -667 -411 -665 -409
rect -637 -412 -635 -410
rect -627 -411 -625 -409
rect -617 -413 -615 -411
rect -606 -405 -604 -403
rect -557 -411 -555 -409
rect -546 -419 -544 -417
rect -535 -411 -533 -409
rect -505 -412 -503 -410
rect -495 -411 -493 -409
rect -485 -413 -483 -411
rect -474 -405 -472 -403
rect -425 -411 -423 -409
rect -414 -419 -412 -417
rect -403 -411 -401 -409
rect -373 -412 -371 -410
rect -363 -411 -361 -409
rect -353 -413 -351 -411
rect -342 -405 -340 -403
rect -259 -403 -257 -401
rect -245 -411 -243 -409
rect -233 -408 -231 -406
rect -757 -445 -755 -443
rect -689 -443 -687 -441
rect -731 -450 -729 -448
rect -703 -447 -701 -445
rect -650 -445 -648 -443
rect -640 -445 -638 -443
rect -557 -443 -555 -441
rect -571 -448 -569 -446
rect -518 -445 -516 -443
rect -428 -442 -426 -440
rect -508 -445 -506 -443
rect -439 -447 -437 -445
rect -389 -444 -387 -442
rect -379 -444 -377 -442
rect -229 -441 -227 -439
<< ndifct1 >>
rect -286 132 -284 134
rect -211 142 -209 144
rect -116 142 -114 144
rect -250 125 -248 127
rect -222 130 -220 132
rect -72 141 -70 143
rect -127 130 -125 132
rect -28 142 -26 144
rect -83 129 -81 131
rect 25 142 27 144
rect -39 130 -37 132
rect 69 142 71 144
rect 14 130 16 132
rect 112 142 114 144
rect 58 130 60 132
rect 101 130 103 132
rect -368 20 -366 22
rect -386 10 -384 12
rect -324 10 -322 12
rect -237 20 -235 22
rect -255 10 -253 12
rect -193 10 -191 12
rect -105 20 -103 22
rect -123 10 -121 12
rect -61 10 -59 12
rect 45 20 47 22
rect 63 10 65 12
rect -339 -1 -337 1
rect -376 -18 -374 -16
rect -243 -1 -241 1
rect -321 -18 -319 -16
rect -282 -18 -280 -16
rect -111 -2 -109 0
rect -225 -18 -223 -16
rect -149 -19 -147 -17
rect 22 -2 24 0
rect -93 -19 -91 -17
rect 11 -14 13 -12
rect -448 -118 -446 -116
rect -420 -122 -418 -120
rect -308 -121 -306 -119
rect -157 -122 -155 -120
rect -409 -134 -407 -132
rect -113 -122 -111 -120
rect -297 -133 -295 -131
rect -146 -134 -144 -132
rect -102 -134 -100 -132
rect -539 -147 -537 -145
rect -521 -157 -519 -155
rect -477 -147 -475 -145
rect -407 -147 -405 -145
rect -389 -157 -387 -155
rect -345 -147 -343 -145
rect -270 -146 -268 -144
rect -252 -156 -250 -154
rect -208 -146 -206 -144
rect -139 -146 -137 -144
rect -121 -156 -119 -154
rect -500 -262 -498 -260
rect -445 -262 -443 -260
rect -407 -262 -405 -260
rect -463 -279 -461 -277
rect -351 -262 -349 -260
rect -234 -261 -232 -259
rect -369 -279 -367 -277
rect -177 -261 -175 -259
rect -139 -266 -137 -264
rect -195 -278 -193 -276
rect -128 -278 -126 -276
rect -565 -291 -563 -289
rect -576 -303 -574 -301
rect -503 -301 -501 -299
rect -379 -301 -377 -299
rect -233 -300 -231 -298
rect -699 -412 -697 -410
rect -717 -422 -715 -420
rect -655 -422 -653 -420
rect -567 -412 -565 -410
rect -585 -422 -583 -420
rect -523 -422 -521 -420
rect -435 -412 -433 -410
rect -453 -422 -451 -420
rect -391 -422 -389 -420
rect -223 -410 -221 -408
rect -205 -420 -203 -418
rect -785 -433 -783 -431
rect -678 -434 -676 -432
rect -767 -443 -765 -441
rect -717 -450 -715 -448
rect -546 -434 -544 -432
rect -660 -451 -658 -449
rect -585 -451 -583 -449
rect -417 -433 -415 -431
rect -528 -451 -526 -449
rect -453 -450 -451 -448
rect -248 -431 -246 -429
rect -399 -450 -397 -448
rect -259 -443 -257 -441
<< ntiect1 >>
rect -273 82 -271 84
rect -265 82 -263 84
rect -249 82 -247 84
rect -237 82 -235 84
rect -221 82 -219 84
rect -126 82 -124 84
rect -82 81 -80 83
rect -38 82 -36 84
rect 15 82 17 84
rect 59 82 61 84
rect 102 82 104 84
rect -269 70 -267 72
rect -138 70 -136 72
rect -6 70 -4 72
rect 43 70 45 72
rect -375 -61 -373 -59
rect -363 -61 -361 -59
rect -281 -61 -279 -59
rect -269 -61 -267 -59
rect -148 -62 -146 -60
rect -136 -62 -134 -60
rect 12 -62 14 -60
rect -447 -75 -445 -73
rect -435 -75 -433 -73
rect -419 -74 -417 -72
rect -307 -73 -305 -71
rect -156 -74 -154 -72
rect -112 -74 -110 -72
rect -422 -207 -420 -205
rect -290 -207 -288 -205
rect -153 -206 -151 -204
rect -119 -206 -117 -204
rect -499 -219 -497 -217
rect -487 -219 -485 -217
rect -406 -219 -404 -217
rect -394 -219 -392 -217
rect -233 -218 -231 -216
rect -221 -218 -219 -216
rect -138 -218 -136 -216
rect -575 -351 -573 -349
rect -490 -351 -488 -349
rect -482 -351 -480 -349
rect -366 -351 -364 -349
rect -358 -351 -356 -349
rect -220 -350 -218 -348
rect -212 -350 -210 -348
rect -600 -362 -598 -360
rect -468 -362 -466 -360
rect -336 -362 -334 -360
rect -225 -360 -223 -358
rect -765 -493 -763 -491
rect -716 -493 -714 -491
rect -704 -493 -702 -491
rect -258 -491 -256 -489
rect -584 -494 -582 -492
rect -572 -494 -570 -492
rect -452 -493 -450 -491
rect -440 -493 -438 -491
<< ptiect1 >>
rect -249 142 -247 144
rect -237 142 -235 144
rect -221 142 -219 144
rect -126 142 -124 144
rect -82 141 -80 143
rect -38 142 -36 144
rect 15 142 17 144
rect 59 142 61 144
rect 102 142 104 144
rect -269 10 -267 12
rect -138 10 -136 12
rect -6 10 -4 12
rect 10 10 12 12
rect -375 -1 -373 1
rect -363 -1 -361 1
rect -281 -1 -279 1
rect -269 -1 -267 1
rect -148 -2 -146 0
rect -136 -2 -134 0
rect 12 -2 14 0
rect -447 -135 -445 -133
rect -435 -135 -433 -133
rect -419 -134 -417 -132
rect -307 -133 -305 -131
rect -156 -134 -154 -132
rect -112 -134 -110 -132
rect -422 -147 -420 -145
rect -290 -147 -288 -145
rect -153 -146 -151 -144
rect -86 -146 -84 -144
rect -499 -279 -497 -277
rect -487 -279 -485 -277
rect -406 -279 -404 -277
rect -394 -279 -392 -277
rect -233 -278 -231 -276
rect -221 -278 -219 -276
rect -138 -278 -136 -276
rect -575 -291 -573 -289
rect -600 -422 -598 -420
rect -468 -422 -466 -420
rect -336 -422 -334 -420
rect -258 -420 -256 -418
rect -732 -433 -730 -431
rect -716 -433 -714 -431
rect -704 -433 -702 -431
rect -584 -434 -582 -432
rect -572 -434 -570 -432
rect -452 -433 -450 -431
rect -440 -433 -438 -431
rect -258 -431 -256 -429
<< pdifct0 >>
rect -286 92 -284 94
rect -275 101 -273 103
rect -275 94 -273 96
rect -264 101 -262 103
rect -264 94 -262 96
rect -239 92 -237 94
rect -212 94 -210 96
rect -202 99 -200 101
rect -202 92 -200 94
rect -192 92 -190 94
rect -117 94 -115 96
rect -107 99 -105 101
rect -107 92 -105 94
rect -97 92 -95 94
rect -73 93 -71 95
rect -63 98 -61 100
rect -63 91 -61 93
rect -53 91 -51 93
rect -29 94 -27 96
rect -19 99 -17 101
rect -19 92 -17 94
rect -9 92 -7 94
rect 24 94 26 96
rect 34 99 36 101
rect 34 92 36 94
rect 44 92 46 94
rect 68 94 70 96
rect 78 99 80 101
rect 78 92 80 94
rect 88 92 90 94
rect 111 94 113 96
rect 121 99 123 101
rect 121 92 123 94
rect 131 92 133 94
rect -386 60 -384 62
rect -366 52 -364 54
rect -366 45 -364 47
rect -356 67 -354 69
rect -346 60 -344 62
rect -336 67 -334 69
rect -336 60 -334 62
rect -326 60 -324 62
rect -316 52 -314 54
rect -306 52 -304 54
rect -306 45 -304 47
rect -296 67 -294 69
rect -285 52 -283 54
rect -275 60 -273 62
rect -255 60 -253 62
rect -235 52 -233 54
rect -235 45 -233 47
rect -225 67 -223 69
rect -215 60 -213 62
rect -205 67 -203 69
rect -205 60 -203 62
rect -195 60 -193 62
rect -185 52 -183 54
rect -175 52 -173 54
rect -175 45 -173 47
rect -165 67 -163 69
rect -154 52 -152 54
rect -144 60 -142 62
rect -123 60 -121 62
rect -103 52 -101 54
rect -103 45 -101 47
rect -93 67 -91 69
rect -83 60 -81 62
rect -73 67 -71 69
rect -73 60 -71 62
rect -63 60 -61 62
rect -53 52 -51 54
rect -43 52 -41 54
rect -43 45 -41 47
rect -33 67 -31 69
rect -22 52 -20 54
rect -12 60 -10 62
rect 17 46 19 48
rect 27 67 29 69
rect 27 60 29 62
rect 43 53 45 55
rect 43 46 45 48
rect 63 61 65 63
rect -365 -51 -363 -49
rect -347 -44 -345 -42
rect -347 -51 -345 -49
rect -337 -50 -335 -48
rect -337 -57 -335 -55
rect -310 -52 -308 -50
rect -300 -49 -298 -47
rect -271 -51 -269 -49
rect -251 -44 -249 -42
rect -251 -51 -249 -49
rect -300 -57 -298 -55
rect -241 -50 -239 -48
rect -241 -57 -239 -55
rect -214 -52 -212 -50
rect -204 -49 -202 -47
rect -204 -57 -202 -55
rect -138 -52 -136 -50
rect -119 -45 -117 -43
rect -119 -52 -117 -50
rect -109 -51 -107 -49
rect -109 -58 -107 -56
rect -82 -53 -80 -51
rect -72 -50 -70 -48
rect 21 -50 23 -48
rect 31 -45 33 -43
rect 31 -52 33 -50
rect 41 -52 43 -50
rect -72 -58 -70 -56
rect -437 -85 -435 -83
rect -410 -86 -408 -84
rect -400 -84 -398 -82
rect -400 -91 -398 -89
rect -390 -84 -388 -82
rect -298 -85 -296 -83
rect -288 -83 -286 -81
rect -288 -90 -286 -88
rect -278 -83 -276 -81
rect -147 -86 -145 -84
rect -137 -84 -135 -82
rect -137 -91 -135 -89
rect -127 -84 -125 -82
rect -103 -86 -101 -84
rect -93 -84 -91 -82
rect -93 -91 -91 -89
rect -83 -84 -81 -82
rect -539 -197 -537 -195
rect -519 -182 -517 -180
rect -519 -189 -517 -187
rect -509 -204 -507 -202
rect -499 -197 -497 -195
rect -489 -197 -487 -195
rect -479 -197 -477 -195
rect -489 -204 -487 -202
rect -469 -189 -467 -187
rect -459 -182 -457 -180
rect -459 -189 -457 -187
rect -438 -189 -436 -187
rect -428 -197 -426 -195
rect -407 -197 -405 -195
rect -449 -204 -447 -202
rect -387 -182 -385 -180
rect -387 -189 -385 -187
rect -377 -204 -375 -202
rect -367 -197 -365 -195
rect -357 -197 -355 -195
rect -347 -197 -345 -195
rect -357 -204 -355 -202
rect -337 -189 -335 -187
rect -327 -182 -325 -180
rect -327 -189 -325 -187
rect -306 -189 -304 -187
rect -296 -197 -294 -195
rect -270 -196 -268 -194
rect -317 -204 -315 -202
rect -250 -181 -248 -179
rect -250 -188 -248 -186
rect -240 -203 -238 -201
rect -230 -196 -228 -194
rect -220 -196 -218 -194
rect -210 -196 -208 -194
rect -220 -203 -218 -201
rect -200 -188 -198 -186
rect -190 -181 -188 -179
rect -190 -188 -188 -186
rect -169 -188 -167 -186
rect -159 -196 -157 -194
rect -139 -197 -137 -195
rect -180 -203 -178 -201
rect -119 -182 -117 -180
rect -119 -189 -117 -187
rect -103 -196 -101 -194
rect -103 -203 -101 -201
rect -93 -182 -91 -180
rect -489 -229 -487 -227
rect -471 -229 -469 -227
rect -471 -236 -469 -234
rect -461 -223 -459 -221
rect -461 -230 -459 -228
rect -434 -228 -432 -226
rect -424 -223 -422 -221
rect -424 -231 -422 -229
rect -396 -229 -394 -227
rect -377 -229 -375 -227
rect -377 -236 -375 -234
rect -367 -223 -365 -221
rect -367 -230 -365 -228
rect -340 -228 -338 -226
rect -330 -223 -328 -221
rect -330 -231 -328 -229
rect -223 -228 -221 -226
rect -203 -228 -201 -226
rect -203 -235 -201 -233
rect -193 -222 -191 -220
rect -193 -229 -191 -227
rect -166 -227 -164 -225
rect -156 -222 -154 -220
rect -156 -230 -154 -228
rect -129 -230 -127 -228
rect -119 -228 -117 -226
rect -119 -235 -117 -233
rect -109 -228 -107 -226
rect -566 -339 -564 -337
rect -556 -334 -554 -332
rect -556 -341 -554 -339
rect -546 -341 -544 -339
rect -503 -341 -501 -339
rect -492 -332 -490 -330
rect -492 -339 -490 -337
rect -481 -332 -479 -330
rect -481 -339 -479 -337
rect -379 -341 -377 -339
rect -368 -332 -366 -330
rect -368 -339 -366 -337
rect -357 -332 -355 -330
rect -357 -339 -355 -337
rect -233 -340 -231 -338
rect -222 -331 -220 -329
rect -222 -338 -220 -336
rect -211 -331 -209 -329
rect -211 -338 -209 -336
rect -717 -372 -715 -370
rect -697 -380 -695 -378
rect -697 -387 -695 -385
rect -687 -365 -685 -363
rect -677 -372 -675 -370
rect -667 -365 -665 -363
rect -667 -372 -665 -370
rect -657 -372 -655 -370
rect -647 -380 -645 -378
rect -637 -380 -635 -378
rect -637 -387 -635 -385
rect -627 -365 -625 -363
rect -616 -380 -614 -378
rect -606 -372 -604 -370
rect -585 -372 -583 -370
rect -565 -380 -563 -378
rect -565 -387 -563 -385
rect -555 -365 -553 -363
rect -545 -372 -543 -370
rect -535 -365 -533 -363
rect -535 -372 -533 -370
rect -525 -372 -523 -370
rect -515 -380 -513 -378
rect -505 -380 -503 -378
rect -505 -387 -503 -385
rect -495 -365 -493 -363
rect -484 -380 -482 -378
rect -474 -372 -472 -370
rect -453 -372 -451 -370
rect -433 -380 -431 -378
rect -433 -387 -431 -385
rect -423 -365 -421 -363
rect -413 -372 -411 -370
rect -403 -365 -401 -363
rect -403 -372 -401 -370
rect -393 -372 -391 -370
rect -383 -380 -381 -378
rect -373 -380 -371 -378
rect -373 -387 -371 -385
rect -363 -365 -361 -363
rect -352 -380 -350 -378
rect -342 -372 -340 -370
rect -251 -384 -249 -382
rect -241 -363 -239 -361
rect -241 -370 -239 -368
rect -225 -377 -223 -375
rect -225 -384 -223 -382
rect -205 -369 -203 -367
rect -785 -484 -783 -482
rect -765 -469 -763 -467
rect -765 -476 -763 -474
rect -739 -469 -737 -467
rect -706 -483 -704 -481
rect -686 -477 -684 -475
rect -686 -484 -684 -482
rect -676 -483 -674 -481
rect -676 -490 -674 -488
rect -649 -485 -647 -483
rect -639 -482 -637 -480
rect -574 -484 -572 -482
rect -554 -477 -552 -475
rect -554 -484 -552 -482
rect -639 -490 -637 -488
rect -544 -483 -542 -481
rect -544 -490 -542 -488
rect -517 -485 -515 -483
rect -507 -482 -505 -480
rect -442 -483 -440 -481
rect -425 -476 -423 -474
rect -425 -483 -423 -481
rect -507 -490 -505 -488
rect -415 -482 -413 -480
rect -415 -489 -413 -487
rect -388 -484 -386 -482
rect -378 -481 -376 -479
rect -249 -479 -247 -477
rect -239 -474 -237 -472
rect -239 -481 -237 -479
rect -229 -481 -227 -479
rect -378 -489 -376 -487
<< pdifct1 >>
rect -250 107 -248 109
rect -250 100 -248 102
rect -222 106 -220 108
rect -222 99 -220 101
rect -127 106 -125 108
rect -127 99 -125 101
rect -83 105 -81 107
rect -83 98 -81 100
rect -39 106 -37 108
rect -39 99 -37 101
rect 14 106 16 108
rect 14 99 16 101
rect 58 106 60 108
rect 58 99 60 101
rect 101 106 103 108
rect 101 99 103 101
rect -376 52 -374 54
rect -245 52 -243 54
rect -113 52 -111 54
rect 53 53 55 55
rect -376 -36 -374 -34
rect -376 -43 -374 -41
rect -320 -36 -318 -34
rect -320 -43 -318 -41
rect -282 -36 -280 -34
rect -282 -43 -280 -41
rect -224 -36 -222 -34
rect -224 -43 -222 -41
rect -149 -37 -147 -35
rect -149 -44 -147 -42
rect -92 -37 -90 -35
rect -92 -44 -90 -42
rect 11 -38 13 -36
rect 11 -45 13 -43
rect -448 -93 -446 -91
rect -448 -100 -446 -98
rect -420 -91 -418 -89
rect -420 -98 -418 -96
rect -308 -90 -306 -88
rect -308 -97 -306 -95
rect -157 -91 -155 -89
rect -157 -98 -155 -96
rect -113 -91 -111 -89
rect -113 -98 -111 -96
rect -529 -189 -527 -187
rect -397 -189 -395 -187
rect -260 -188 -258 -186
rect -129 -189 -127 -187
rect -500 -237 -498 -235
rect -500 -244 -498 -242
rect -444 -237 -442 -235
rect -444 -244 -442 -242
rect -407 -237 -405 -235
rect -407 -244 -405 -242
rect -350 -237 -348 -235
rect -350 -244 -348 -242
rect -234 -236 -232 -234
rect -234 -243 -232 -241
rect -176 -236 -174 -234
rect -176 -243 -174 -241
rect -139 -235 -137 -233
rect -139 -242 -137 -240
rect -576 -327 -574 -325
rect -576 -334 -574 -332
rect -707 -380 -705 -378
rect -575 -380 -573 -378
rect -443 -380 -441 -378
rect -215 -377 -213 -375
rect -775 -476 -773 -474
rect -749 -483 -747 -481
rect -749 -490 -747 -488
rect -717 -468 -715 -466
rect -717 -475 -715 -473
rect -659 -469 -657 -467
rect -659 -476 -657 -474
rect -585 -469 -583 -467
rect -585 -476 -583 -474
rect -527 -469 -525 -467
rect -527 -476 -525 -474
rect -453 -468 -451 -466
rect -453 -475 -451 -473
rect -398 -468 -396 -466
rect -398 -475 -396 -473
rect -259 -467 -257 -465
rect -259 -474 -257 -472
<< alu0 >>
rect -265 140 -261 141
rect -265 138 -264 140
rect -262 138 -261 140
rect -265 136 -261 138
rect -237 130 -233 141
rect -248 123 -247 129
rect -237 128 -236 130
rect -234 128 -233 130
rect -237 126 -233 128
rect -208 134 -188 135
rect -208 132 -192 134
rect -190 132 -188 134
rect -208 131 -188 132
rect -220 128 -219 130
rect -208 127 -204 131
rect -113 134 -93 135
rect -113 132 -97 134
rect -95 132 -93 134
rect -113 131 -93 132
rect -248 104 -247 111
rect -216 123 -204 127
rect -216 118 -212 123
rect -125 128 -124 130
rect -113 127 -109 131
rect -69 133 -49 134
rect -69 131 -53 133
rect -51 131 -49 133
rect -69 130 -49 131
rect -25 134 -5 135
rect -25 132 -9 134
rect -7 132 -5 134
rect -25 131 -5 132
rect -216 116 -215 118
rect -213 116 -212 118
rect -284 103 -271 104
rect -273 101 -271 103
rect -275 99 -271 101
rect -277 96 -271 99
rect -288 94 -282 95
rect -288 92 -286 94
rect -284 92 -282 94
rect -277 94 -275 96
rect -273 94 -271 96
rect -277 93 -271 94
rect -266 103 -260 104
rect -266 101 -264 103
rect -262 101 -260 103
rect -266 96 -260 101
rect -216 104 -212 116
rect -216 101 -199 104
rect -216 100 -202 101
rect -203 99 -202 100
rect -200 99 -199 101
rect -266 94 -264 96
rect -262 94 -260 96
rect -214 96 -208 97
rect -288 85 -282 92
rect -266 85 -260 94
rect -241 94 -235 95
rect -241 92 -239 94
rect -237 92 -235 94
rect -241 85 -235 92
rect -214 94 -212 96
rect -210 94 -208 96
rect -214 85 -208 94
rect -203 94 -199 99
rect -121 123 -109 127
rect -121 118 -117 123
rect -121 116 -120 118
rect -118 116 -117 118
rect -121 104 -117 116
rect -121 101 -104 104
rect -121 100 -107 101
rect -108 99 -107 100
rect -105 99 -104 101
rect -119 96 -113 97
rect -203 92 -202 94
rect -200 92 -199 94
rect -203 90 -199 92
rect -194 94 -188 95
rect -194 92 -192 94
rect -190 92 -188 94
rect -194 85 -188 92
rect -119 94 -117 96
rect -115 94 -113 96
rect -119 85 -113 94
rect -108 94 -104 99
rect -81 127 -80 129
rect -69 126 -65 130
rect -77 122 -65 126
rect -77 117 -73 122
rect -77 115 -76 117
rect -74 115 -73 117
rect -77 103 -73 115
rect -37 128 -36 130
rect -25 127 -21 131
rect 28 134 48 135
rect 28 132 44 134
rect 46 132 48 134
rect 28 131 48 132
rect -33 123 -21 127
rect -33 118 -29 123
rect -33 116 -32 118
rect -30 116 -29 118
rect -77 100 -60 103
rect -77 99 -63 100
rect -64 98 -63 99
rect -61 98 -60 100
rect -75 95 -69 96
rect -108 92 -107 94
rect -105 92 -104 94
rect -108 90 -104 92
rect -99 94 -93 95
rect -99 92 -97 94
rect -95 92 -93 94
rect -99 85 -93 92
rect -75 93 -73 95
rect -71 93 -69 95
rect -75 84 -69 93
rect -64 93 -60 98
rect -33 104 -29 116
rect 16 128 17 130
rect 28 127 32 131
rect 72 134 92 135
rect 72 132 88 134
rect 90 132 92 134
rect 72 131 92 132
rect -33 101 -16 104
rect -33 100 -19 101
rect -20 99 -19 100
rect -17 99 -16 101
rect -31 96 -25 97
rect -31 94 -29 96
rect -27 94 -25 96
rect -64 91 -63 93
rect -61 91 -60 93
rect -64 89 -60 91
rect -55 93 -49 94
rect -55 91 -53 93
rect -51 91 -49 93
rect -55 84 -49 91
rect -31 85 -25 94
rect -20 94 -16 99
rect 20 123 32 127
rect 20 118 24 123
rect 20 116 21 118
rect 23 116 24 118
rect 20 104 24 116
rect 60 128 61 130
rect 72 127 76 131
rect 115 134 135 135
rect 115 132 131 134
rect 133 132 135 134
rect 115 131 135 132
rect 20 101 37 104
rect 20 100 34 101
rect 33 99 34 100
rect 36 99 37 101
rect 22 96 28 97
rect -20 92 -19 94
rect -17 92 -16 94
rect -20 90 -16 92
rect -11 94 -5 95
rect -11 92 -9 94
rect -7 92 -5 94
rect -11 85 -5 92
rect 22 94 24 96
rect 26 94 28 96
rect 22 85 28 94
rect 33 94 37 99
rect 64 123 76 127
rect 64 118 68 123
rect 64 116 65 118
rect 67 116 68 118
rect 64 104 68 116
rect 64 101 81 104
rect 64 100 78 101
rect 77 99 78 100
rect 80 99 81 101
rect 66 96 72 97
rect 33 92 34 94
rect 36 92 37 94
rect 33 90 37 92
rect 42 94 48 95
rect 42 92 44 94
rect 46 92 48 94
rect 42 85 48 92
rect 66 94 68 96
rect 70 94 72 96
rect 66 85 72 94
rect 77 94 81 99
rect 103 128 104 130
rect 115 127 119 131
rect 107 123 119 127
rect 107 118 111 123
rect 107 116 108 118
rect 110 116 111 118
rect 107 104 111 116
rect 107 101 124 104
rect 107 100 121 101
rect 120 99 121 100
rect 123 99 124 101
rect 109 96 115 97
rect 77 92 78 94
rect 80 92 81 94
rect 77 90 81 92
rect 86 94 92 95
rect 86 92 88 94
rect 90 92 92 94
rect 86 85 92 92
rect 109 94 111 96
rect 113 94 115 96
rect 109 85 115 94
rect 120 94 124 99
rect 120 92 121 94
rect 123 92 124 94
rect 120 90 124 92
rect 129 94 135 95
rect 129 92 131 94
rect 133 92 135 94
rect 129 85 135 92
rect -358 67 -356 69
rect -354 67 -352 69
rect -358 66 -352 67
rect -338 67 -336 69
rect -334 67 -332 69
rect -388 62 -342 63
rect -388 60 -386 62
rect -384 60 -346 62
rect -344 60 -342 62
rect -388 59 -342 60
rect -338 62 -332 67
rect -298 67 -296 69
rect -294 67 -292 69
rect -298 66 -292 67
rect -338 60 -336 62
rect -334 60 -332 62
rect -338 59 -332 60
rect -328 62 -296 63
rect -328 60 -326 62
rect -324 60 -296 62
rect -328 59 -296 60
rect -277 62 -271 69
rect -227 67 -225 69
rect -223 67 -221 69
rect -227 66 -221 67
rect -207 67 -205 69
rect -203 67 -201 69
rect -277 60 -275 62
rect -273 60 -271 62
rect -277 59 -271 60
rect -257 62 -211 63
rect -257 60 -255 62
rect -253 60 -215 62
rect -213 60 -211 62
rect -257 59 -211 60
rect -207 62 -201 67
rect -167 67 -165 69
rect -163 67 -161 69
rect -167 66 -161 67
rect -207 60 -205 62
rect -203 60 -201 62
rect -207 59 -201 60
rect -197 62 -165 63
rect -197 60 -195 62
rect -193 60 -165 62
rect -197 59 -165 60
rect -146 62 -140 69
rect -95 67 -93 69
rect -91 67 -89 69
rect -95 66 -89 67
rect -75 67 -73 69
rect -71 67 -69 69
rect -146 60 -144 62
rect -142 60 -140 62
rect -146 59 -140 60
rect -125 62 -79 63
rect -125 60 -123 62
rect -121 60 -83 62
rect -81 60 -79 62
rect -125 59 -79 60
rect -75 62 -69 67
rect -35 67 -33 69
rect -31 67 -29 69
rect -35 66 -29 67
rect -75 60 -73 62
rect -71 60 -69 62
rect -75 59 -69 60
rect -65 62 -33 63
rect -65 60 -63 62
rect -61 60 -33 62
rect -65 59 -33 60
rect -14 62 -8 69
rect 26 67 27 69
rect 29 67 30 69
rect -14 60 -12 62
rect -10 60 -8 62
rect -14 59 -8 60
rect -368 54 -362 55
rect -368 52 -366 54
rect -364 52 -362 54
rect -368 48 -362 52
rect -380 47 -362 48
rect -380 45 -366 47
rect -364 45 -362 47
rect -380 44 -362 45
rect -380 38 -376 44
rect -358 39 -354 59
rect -300 56 -296 59
rect -380 36 -379 38
rect -377 36 -376 38
rect -380 31 -376 36
rect -371 38 -345 39
rect -371 36 -369 38
rect -367 36 -345 38
rect -371 35 -345 36
rect -380 27 -355 31
rect -359 23 -355 27
rect -359 21 -358 23
rect -356 21 -355 23
rect -359 19 -355 21
rect -349 24 -345 35
rect -328 54 -312 55
rect -328 52 -316 54
rect -314 52 -312 54
rect -328 51 -312 52
rect -307 54 -303 56
rect -307 52 -306 54
rect -304 52 -303 54
rect -328 39 -324 51
rect -307 47 -303 52
rect -331 38 -324 39
rect -331 36 -329 38
rect -327 36 -324 38
rect -331 35 -324 36
rect -349 23 -332 24
rect -349 21 -336 23
rect -334 21 -332 23
rect -349 20 -332 21
rect -328 23 -324 35
rect -320 45 -306 47
rect -304 45 -303 47
rect -320 43 -303 45
rect -300 54 -282 56
rect -300 52 -285 54
rect -283 52 -282 54
rect -320 38 -316 43
rect -300 39 -296 52
rect -286 47 -282 52
rect -286 43 -272 47
rect -320 36 -319 38
rect -317 36 -316 38
rect -320 31 -316 36
rect -311 38 -296 39
rect -311 36 -309 38
rect -307 36 -296 38
rect -311 35 -296 36
rect -320 27 -293 31
rect -276 29 -272 43
rect -237 54 -231 55
rect -237 52 -235 54
rect -233 52 -231 54
rect -276 27 -275 29
rect -273 27 -272 29
rect -297 23 -293 27
rect -276 25 -272 27
rect -237 48 -231 52
rect -249 47 -231 48
rect -249 45 -235 47
rect -233 45 -231 47
rect -249 44 -231 45
rect -249 38 -245 44
rect -227 39 -223 59
rect -169 56 -165 59
rect -249 36 -248 38
rect -246 36 -245 38
rect -249 31 -245 36
rect -240 38 -214 39
rect -240 36 -238 38
rect -236 36 -214 38
rect -240 35 -214 36
rect -249 27 -224 31
rect -228 23 -224 27
rect -328 22 -302 23
rect -328 20 -306 22
rect -304 20 -302 22
rect -328 19 -302 20
rect -297 21 -296 23
rect -294 21 -293 23
rect -297 19 -293 21
rect -287 21 -283 23
rect -287 19 -286 21
rect -284 19 -283 21
rect -228 21 -227 23
rect -225 21 -224 23
rect -228 19 -224 21
rect -218 24 -214 35
rect -197 54 -181 55
rect -197 52 -185 54
rect -183 52 -181 54
rect -197 51 -181 52
rect -176 54 -172 56
rect -176 52 -175 54
rect -173 52 -172 54
rect -197 39 -193 51
rect -176 47 -172 52
rect -200 38 -193 39
rect -200 36 -198 38
rect -196 36 -193 38
rect -200 35 -193 36
rect -218 23 -201 24
rect -218 21 -205 23
rect -203 21 -201 23
rect -218 20 -201 21
rect -197 23 -193 35
rect -189 45 -175 47
rect -173 45 -172 47
rect -189 43 -172 45
rect -169 54 -151 56
rect -169 52 -154 54
rect -152 52 -151 54
rect -189 38 -185 43
rect -169 39 -165 52
rect -155 47 -151 52
rect -155 43 -141 47
rect -189 36 -188 38
rect -186 36 -185 38
rect -189 31 -185 36
rect -180 38 -165 39
rect -180 36 -178 38
rect -176 36 -165 38
rect -180 35 -165 36
rect -189 27 -162 31
rect -145 29 -141 43
rect -105 54 -99 55
rect -105 52 -103 54
rect -101 52 -99 54
rect -145 27 -144 29
rect -142 27 -141 29
rect -166 23 -162 27
rect -145 25 -141 27
rect -105 48 -99 52
rect -117 47 -99 48
rect -117 45 -103 47
rect -101 45 -99 47
rect -117 44 -99 45
rect -117 38 -113 44
rect -95 39 -91 59
rect -37 56 -33 59
rect 26 62 30 67
rect 26 60 27 62
rect 29 60 30 62
rect 26 58 30 60
rect 34 63 67 64
rect 34 61 63 63
rect 65 61 67 63
rect 34 60 67 61
rect -117 36 -116 38
rect -114 36 -113 38
rect -117 31 -113 36
rect -108 38 -82 39
rect -108 36 -106 38
rect -104 36 -82 38
rect -108 35 -82 36
rect -117 27 -92 31
rect -96 23 -92 27
rect -197 22 -171 23
rect -197 20 -175 22
rect -173 20 -171 22
rect -197 19 -171 20
rect -166 21 -165 23
rect -163 21 -162 23
rect -166 19 -162 21
rect -156 21 -152 23
rect -156 19 -155 21
rect -153 19 -152 21
rect -96 21 -95 23
rect -93 21 -92 23
rect -96 19 -92 21
rect -86 24 -82 35
rect -65 54 -49 55
rect -65 52 -53 54
rect -51 52 -49 54
rect -65 51 -49 52
rect -44 54 -40 56
rect -44 52 -43 54
rect -41 52 -40 54
rect -65 39 -61 51
rect -44 47 -40 52
rect -68 38 -61 39
rect -68 36 -66 38
rect -64 36 -61 38
rect -68 35 -61 36
rect -86 23 -69 24
rect -86 21 -73 23
rect -71 21 -69 23
rect -86 20 -69 21
rect -65 23 -61 35
rect -57 45 -43 47
rect -41 45 -40 47
rect -57 43 -40 45
rect -37 54 -19 56
rect -37 52 -22 54
rect -20 52 -19 54
rect -57 38 -53 43
rect -37 39 -33 52
rect -23 47 -19 52
rect -23 43 -9 47
rect -57 36 -56 38
rect -54 36 -53 38
rect -57 31 -53 36
rect -48 38 -33 39
rect -48 36 -46 38
rect -44 36 -33 38
rect -48 35 -33 36
rect -57 27 -30 31
rect -13 29 -9 43
rect 34 49 38 60
rect 15 48 38 49
rect 15 46 17 48
rect 19 46 38 48
rect 15 45 38 46
rect 15 39 19 45
rect 8 35 19 39
rect -13 27 -12 29
rect -10 27 -9 29
rect -34 23 -30 27
rect -13 25 -9 27
rect 8 29 12 35
rect 34 39 38 45
rect 42 55 46 57
rect 42 53 43 55
rect 45 53 46 55
rect 42 48 46 53
rect 42 46 43 48
rect 45 47 46 48
rect 45 46 58 47
rect 42 43 58 46
rect 54 41 58 43
rect 54 39 59 41
rect 34 38 50 39
rect 34 36 46 38
rect 48 36 50 38
rect 34 35 50 36
rect 54 37 56 39
rect 58 37 59 39
rect 54 35 59 37
rect 8 27 9 29
rect 11 27 12 29
rect 8 25 12 27
rect 54 31 58 35
rect 34 27 58 31
rect 34 24 38 27
rect -65 22 -39 23
rect -65 20 -43 22
rect -41 20 -39 22
rect -65 19 -39 20
rect -34 21 -33 23
rect -31 21 -30 23
rect -34 19 -30 21
rect -24 21 -20 23
rect 34 22 35 24
rect 37 22 38 24
rect -24 19 -23 21
rect -21 19 -20 21
rect -349 15 -343 16
rect -349 13 -347 15
rect -345 13 -343 15
rect -287 13 -283 19
rect -218 15 -212 16
rect -218 13 -216 15
rect -214 13 -212 15
rect -156 13 -152 19
rect -86 15 -80 16
rect -86 13 -84 15
rect -82 13 -80 15
rect -24 13 -20 19
rect 21 21 27 22
rect 21 19 23 21
rect 25 19 27 21
rect 34 20 38 22
rect 21 13 27 19
rect -363 -13 -359 -2
rect -352 -8 -307 -7
rect -352 -10 -350 -8
rect -348 -10 -307 -8
rect -352 -11 -311 -10
rect -313 -12 -311 -11
rect -309 -12 -307 -10
rect -313 -13 -307 -12
rect -303 -10 -297 -2
rect -303 -12 -301 -10
rect -299 -12 -297 -10
rect -303 -13 -297 -12
rect -374 -20 -373 -14
rect -363 -15 -362 -13
rect -360 -15 -359 -13
rect -363 -17 -359 -15
rect -269 -13 -265 -2
rect -256 -8 -211 -7
rect -256 -10 -254 -8
rect -252 -10 -211 -8
rect -256 -11 -215 -10
rect -217 -12 -215 -11
rect -213 -12 -211 -10
rect -217 -13 -211 -12
rect -207 -10 -201 -2
rect -207 -12 -205 -10
rect -203 -12 -201 -10
rect -207 -13 -201 -12
rect -280 -20 -279 -14
rect -269 -15 -268 -13
rect -266 -15 -265 -13
rect -374 -39 -373 -32
rect -269 -17 -265 -15
rect -136 -14 -132 -3
rect -124 -9 -79 -8
rect -124 -11 -122 -9
rect -120 -11 -79 -9
rect -124 -12 -83 -11
rect -85 -13 -83 -12
rect -81 -13 -79 -11
rect -85 -14 -79 -13
rect -75 -11 -69 -3
rect -75 -13 -73 -11
rect -71 -13 -69 -11
rect -75 -14 -69 -13
rect 25 -10 45 -9
rect 25 -12 41 -10
rect 43 -12 45 -10
rect 25 -13 45 -12
rect -348 -42 -326 -40
rect -348 -44 -347 -42
rect -345 -44 -326 -42
rect -367 -49 -361 -48
rect -367 -51 -365 -49
rect -363 -51 -361 -49
rect -367 -58 -361 -51
rect -348 -49 -344 -44
rect -348 -51 -347 -49
rect -345 -51 -344 -49
rect -348 -53 -344 -51
rect -339 -48 -333 -47
rect -339 -50 -337 -48
rect -335 -50 -333 -48
rect -339 -55 -333 -50
rect -330 -49 -326 -44
rect -280 -39 -279 -32
rect -147 -21 -146 -15
rect -136 -16 -135 -14
rect -133 -16 -132 -14
rect 13 -16 14 -14
rect -252 -42 -230 -40
rect -252 -44 -251 -42
rect -249 -44 -230 -42
rect -301 -47 -297 -45
rect -301 -49 -300 -47
rect -298 -49 -297 -47
rect -330 -50 -306 -49
rect -330 -52 -310 -50
rect -308 -52 -306 -50
rect -330 -53 -306 -52
rect -339 -57 -337 -55
rect -335 -57 -333 -55
rect -339 -58 -333 -57
rect -301 -55 -297 -49
rect -301 -57 -300 -55
rect -298 -57 -297 -55
rect -301 -58 -297 -57
rect -273 -49 -267 -48
rect -273 -51 -271 -49
rect -269 -51 -267 -49
rect -273 -58 -267 -51
rect -252 -49 -248 -44
rect -252 -51 -251 -49
rect -249 -51 -248 -49
rect -252 -53 -248 -51
rect -243 -48 -237 -47
rect -243 -50 -241 -48
rect -239 -50 -237 -48
rect -243 -55 -237 -50
rect -234 -49 -230 -44
rect -136 -18 -132 -16
rect 25 -17 29 -13
rect -147 -40 -146 -33
rect -205 -47 -201 -45
rect -120 -43 -98 -41
rect -120 -45 -119 -43
rect -117 -45 -98 -43
rect -205 -49 -204 -47
rect -202 -49 -201 -47
rect -234 -50 -210 -49
rect -234 -52 -214 -50
rect -212 -52 -210 -50
rect -234 -53 -210 -52
rect -243 -57 -241 -55
rect -239 -57 -237 -55
rect -243 -58 -237 -57
rect -205 -55 -201 -49
rect -205 -57 -204 -55
rect -202 -57 -201 -55
rect -205 -58 -201 -57
rect -140 -50 -134 -49
rect -140 -52 -138 -50
rect -136 -52 -134 -50
rect -140 -59 -134 -52
rect -120 -50 -116 -45
rect -120 -52 -119 -50
rect -117 -52 -116 -50
rect -120 -54 -116 -52
rect -111 -49 -105 -48
rect -111 -51 -109 -49
rect -107 -51 -105 -49
rect -111 -56 -105 -51
rect -102 -50 -98 -45
rect 17 -21 29 -17
rect 17 -26 21 -21
rect 17 -28 18 -26
rect 20 -28 21 -26
rect 17 -40 21 -28
rect 17 -43 34 -40
rect 17 -44 31 -43
rect -73 -48 -69 -46
rect 30 -45 31 -44
rect 33 -45 34 -43
rect -73 -50 -72 -48
rect -70 -50 -69 -48
rect -102 -51 -78 -50
rect -102 -53 -82 -51
rect -80 -53 -78 -51
rect -102 -54 -78 -53
rect -111 -58 -109 -56
rect -107 -58 -105 -56
rect -111 -59 -105 -58
rect -73 -56 -69 -50
rect -73 -58 -72 -56
rect -70 -58 -69 -56
rect -73 -59 -69 -58
rect 19 -48 25 -47
rect 19 -50 21 -48
rect 23 -50 25 -48
rect 19 -59 25 -50
rect 30 -50 34 -45
rect 30 -52 31 -50
rect 33 -52 34 -50
rect 30 -54 34 -52
rect 39 -50 45 -49
rect 39 -52 41 -50
rect 43 -52 45 -50
rect 39 -59 45 -52
rect -439 -83 -433 -76
rect -439 -85 -437 -83
rect -435 -85 -433 -83
rect -439 -86 -433 -85
rect -412 -84 -406 -75
rect -412 -86 -410 -84
rect -408 -86 -406 -84
rect -412 -87 -406 -86
rect -401 -82 -397 -80
rect -401 -84 -400 -82
rect -398 -84 -397 -82
rect -401 -89 -397 -84
rect -392 -82 -386 -75
rect -392 -84 -390 -82
rect -388 -84 -386 -82
rect -392 -85 -386 -84
rect -300 -83 -294 -74
rect -300 -85 -298 -83
rect -296 -85 -294 -83
rect -300 -86 -294 -85
rect -289 -81 -285 -79
rect -289 -83 -288 -81
rect -286 -83 -285 -81
rect -401 -90 -400 -89
rect -446 -102 -445 -95
rect -414 -91 -400 -90
rect -398 -91 -397 -89
rect -414 -94 -397 -91
rect -446 -120 -445 -114
rect -435 -119 -431 -117
rect -435 -121 -434 -119
rect -432 -121 -431 -119
rect -435 -132 -431 -121
rect -414 -106 -410 -94
rect -289 -88 -285 -83
rect -280 -81 -274 -74
rect -280 -83 -278 -81
rect -276 -83 -274 -81
rect -280 -84 -274 -83
rect -149 -84 -143 -75
rect -149 -86 -147 -84
rect -145 -86 -143 -84
rect -149 -87 -143 -86
rect -138 -82 -134 -80
rect -138 -84 -137 -82
rect -135 -84 -134 -82
rect -289 -89 -288 -88
rect -302 -90 -288 -89
rect -286 -90 -285 -88
rect -302 -93 -285 -90
rect -414 -108 -413 -106
rect -411 -108 -410 -106
rect -414 -113 -410 -108
rect -414 -117 -402 -113
rect -418 -120 -417 -118
rect -406 -121 -402 -117
rect -302 -105 -298 -93
rect -138 -89 -134 -84
rect -129 -82 -123 -75
rect -129 -84 -127 -82
rect -125 -84 -123 -82
rect -129 -85 -123 -84
rect -105 -84 -99 -75
rect -105 -86 -103 -84
rect -101 -86 -99 -84
rect -105 -87 -99 -86
rect -94 -82 -90 -80
rect -94 -84 -93 -82
rect -91 -84 -90 -82
rect -138 -90 -137 -89
rect -151 -91 -137 -90
rect -135 -91 -134 -89
rect -151 -94 -134 -91
rect -302 -107 -301 -105
rect -299 -107 -298 -105
rect -302 -112 -298 -107
rect -302 -116 -290 -112
rect -306 -119 -305 -117
rect -406 -122 -386 -121
rect -406 -124 -390 -122
rect -388 -124 -386 -122
rect -406 -125 -386 -124
rect -294 -120 -290 -116
rect -151 -106 -147 -94
rect -94 -89 -90 -84
rect -85 -82 -79 -75
rect -85 -84 -83 -82
rect -81 -84 -79 -82
rect -85 -85 -79 -84
rect -94 -90 -93 -89
rect -107 -91 -93 -90
rect -91 -91 -90 -89
rect -107 -94 -90 -91
rect -151 -108 -150 -106
rect -148 -108 -147 -106
rect -151 -113 -147 -108
rect -151 -117 -139 -113
rect -155 -120 -154 -118
rect -294 -121 -274 -120
rect -294 -123 -278 -121
rect -276 -123 -274 -121
rect -294 -124 -274 -123
rect -143 -121 -139 -117
rect -107 -106 -103 -94
rect -107 -108 -106 -106
rect -104 -108 -103 -106
rect -107 -113 -103 -108
rect -107 -117 -95 -113
rect -111 -120 -110 -118
rect -143 -122 -123 -121
rect -143 -124 -127 -122
rect -125 -124 -123 -122
rect -143 -125 -123 -124
rect -99 -121 -95 -117
rect -99 -122 -79 -121
rect -99 -124 -83 -122
rect -81 -124 -79 -122
rect -99 -125 -79 -124
rect -502 -150 -500 -148
rect -498 -150 -496 -148
rect -502 -151 -496 -150
rect -440 -154 -436 -148
rect -370 -150 -368 -148
rect -366 -150 -364 -148
rect -370 -151 -364 -150
rect -308 -154 -304 -148
rect -233 -149 -231 -147
rect -229 -149 -227 -147
rect -233 -150 -227 -149
rect -171 -153 -167 -147
rect -101 -153 -95 -147
rect -512 -156 -508 -154
rect -481 -155 -455 -154
rect -512 -158 -511 -156
rect -509 -158 -508 -156
rect -512 -162 -508 -158
rect -533 -166 -508 -162
rect -502 -156 -485 -155
rect -502 -158 -489 -156
rect -487 -158 -485 -156
rect -502 -159 -485 -158
rect -481 -157 -459 -155
rect -457 -157 -455 -155
rect -481 -158 -455 -157
rect -450 -156 -446 -154
rect -450 -158 -449 -156
rect -447 -158 -446 -156
rect -440 -156 -439 -154
rect -437 -156 -436 -154
rect -440 -158 -436 -156
rect -380 -156 -376 -154
rect -349 -155 -323 -154
rect -380 -158 -379 -156
rect -377 -158 -376 -156
rect -533 -171 -529 -166
rect -502 -170 -498 -159
rect -533 -173 -532 -171
rect -530 -173 -529 -171
rect -533 -179 -529 -173
rect -524 -171 -498 -170
rect -524 -173 -522 -171
rect -520 -173 -498 -171
rect -524 -174 -498 -173
rect -481 -170 -477 -158
rect -450 -162 -446 -158
rect -429 -162 -425 -160
rect -533 -180 -515 -179
rect -533 -182 -519 -180
rect -517 -182 -515 -180
rect -533 -183 -515 -182
rect -521 -187 -515 -183
rect -521 -189 -519 -187
rect -517 -189 -515 -187
rect -521 -190 -515 -189
rect -511 -194 -507 -174
rect -484 -171 -477 -170
rect -484 -173 -482 -171
rect -480 -173 -477 -171
rect -484 -174 -477 -173
rect -481 -186 -477 -174
rect -473 -166 -446 -162
rect -473 -171 -469 -166
rect -473 -173 -472 -171
rect -470 -173 -469 -171
rect -473 -178 -469 -173
rect -464 -171 -449 -170
rect -464 -173 -462 -171
rect -460 -173 -449 -171
rect -464 -174 -449 -173
rect -473 -180 -456 -178
rect -473 -182 -459 -180
rect -457 -182 -456 -180
rect -481 -187 -465 -186
rect -481 -189 -469 -187
rect -467 -189 -465 -187
rect -481 -190 -465 -189
rect -460 -187 -456 -182
rect -460 -189 -459 -187
rect -457 -189 -456 -187
rect -460 -191 -456 -189
rect -453 -187 -449 -174
rect -429 -164 -428 -162
rect -426 -164 -425 -162
rect -429 -178 -425 -164
rect -439 -182 -425 -178
rect -439 -187 -435 -182
rect -453 -189 -438 -187
rect -436 -189 -435 -187
rect -453 -191 -435 -189
rect -380 -162 -376 -158
rect -401 -166 -376 -162
rect -370 -156 -353 -155
rect -370 -158 -357 -156
rect -355 -158 -353 -156
rect -370 -159 -353 -158
rect -349 -157 -327 -155
rect -325 -157 -323 -155
rect -349 -158 -323 -157
rect -318 -156 -314 -154
rect -318 -158 -317 -156
rect -315 -158 -314 -156
rect -308 -156 -307 -154
rect -305 -156 -304 -154
rect -308 -158 -304 -156
rect -243 -155 -239 -153
rect -212 -154 -186 -153
rect -243 -157 -242 -155
rect -240 -157 -239 -155
rect -401 -171 -397 -166
rect -370 -170 -366 -159
rect -401 -173 -400 -171
rect -398 -173 -397 -171
rect -401 -179 -397 -173
rect -392 -171 -366 -170
rect -392 -173 -390 -171
rect -388 -173 -366 -171
rect -392 -174 -366 -173
rect -349 -170 -345 -158
rect -318 -162 -314 -158
rect -297 -162 -293 -160
rect -401 -180 -383 -179
rect -401 -182 -387 -180
rect -385 -182 -383 -180
rect -401 -183 -383 -182
rect -389 -187 -383 -183
rect -389 -189 -387 -187
rect -385 -189 -383 -187
rect -389 -190 -383 -189
rect -453 -194 -449 -191
rect -379 -194 -375 -174
rect -352 -171 -345 -170
rect -352 -173 -350 -171
rect -348 -173 -345 -171
rect -352 -174 -345 -173
rect -349 -186 -345 -174
rect -341 -166 -314 -162
rect -341 -171 -337 -166
rect -341 -173 -340 -171
rect -338 -173 -337 -171
rect -341 -178 -337 -173
rect -332 -171 -317 -170
rect -332 -173 -330 -171
rect -328 -173 -317 -171
rect -332 -174 -317 -173
rect -341 -180 -324 -178
rect -341 -182 -327 -180
rect -325 -182 -324 -180
rect -349 -187 -333 -186
rect -349 -189 -337 -187
rect -335 -189 -333 -187
rect -349 -190 -333 -189
rect -328 -187 -324 -182
rect -328 -189 -327 -187
rect -325 -189 -324 -187
rect -328 -191 -324 -189
rect -321 -187 -317 -174
rect -297 -164 -296 -162
rect -294 -164 -293 -162
rect -297 -178 -293 -164
rect -307 -182 -293 -178
rect -307 -187 -303 -182
rect -321 -189 -306 -187
rect -304 -189 -303 -187
rect -321 -191 -303 -189
rect -243 -161 -239 -157
rect -264 -165 -239 -161
rect -233 -155 -216 -154
rect -233 -157 -220 -155
rect -218 -157 -216 -155
rect -233 -158 -216 -157
rect -212 -156 -190 -154
rect -188 -156 -186 -154
rect -212 -157 -186 -156
rect -181 -155 -177 -153
rect -181 -157 -180 -155
rect -178 -157 -177 -155
rect -171 -155 -170 -153
rect -168 -155 -167 -153
rect -171 -157 -167 -155
rect -112 -156 -108 -154
rect -101 -155 -99 -153
rect -97 -155 -95 -153
rect -101 -156 -95 -155
rect -264 -170 -260 -165
rect -233 -169 -229 -158
rect -264 -172 -263 -170
rect -261 -172 -260 -170
rect -264 -178 -260 -172
rect -255 -170 -229 -169
rect -255 -172 -253 -170
rect -251 -172 -229 -170
rect -255 -173 -229 -172
rect -212 -169 -208 -157
rect -181 -161 -177 -157
rect -160 -161 -156 -159
rect -264 -179 -246 -178
rect -264 -181 -250 -179
rect -248 -181 -246 -179
rect -264 -182 -246 -181
rect -252 -186 -246 -182
rect -252 -188 -250 -186
rect -248 -188 -246 -186
rect -252 -189 -246 -188
rect -321 -194 -317 -191
rect -242 -193 -238 -173
rect -215 -170 -208 -169
rect -215 -172 -213 -170
rect -211 -172 -208 -170
rect -215 -173 -208 -172
rect -212 -185 -208 -173
rect -204 -165 -177 -161
rect -204 -170 -200 -165
rect -204 -172 -203 -170
rect -201 -172 -200 -170
rect -204 -177 -200 -172
rect -195 -170 -180 -169
rect -195 -172 -193 -170
rect -191 -172 -180 -170
rect -195 -173 -180 -172
rect -204 -179 -187 -177
rect -204 -181 -190 -179
rect -188 -181 -187 -179
rect -212 -186 -196 -185
rect -212 -188 -200 -186
rect -198 -188 -196 -186
rect -212 -189 -196 -188
rect -191 -186 -187 -181
rect -191 -188 -190 -186
rect -188 -188 -187 -186
rect -191 -190 -187 -188
rect -184 -186 -180 -173
rect -160 -163 -159 -161
rect -157 -163 -156 -161
rect -160 -177 -156 -163
rect -170 -181 -156 -177
rect -170 -186 -166 -181
rect -184 -188 -169 -186
rect -167 -188 -166 -186
rect -184 -190 -166 -188
rect -112 -158 -111 -156
rect -109 -158 -108 -156
rect -112 -161 -108 -158
rect -132 -165 -108 -161
rect -132 -169 -128 -165
rect -86 -161 -82 -159
rect -86 -163 -85 -161
rect -83 -163 -82 -161
rect -133 -171 -128 -169
rect -133 -173 -132 -171
rect -130 -173 -128 -171
rect -124 -170 -108 -169
rect -124 -172 -122 -170
rect -120 -172 -108 -170
rect -124 -173 -108 -172
rect -133 -175 -128 -173
rect -132 -177 -128 -175
rect -132 -180 -116 -177
rect -132 -181 -119 -180
rect -120 -182 -119 -181
rect -117 -182 -116 -180
rect -120 -187 -116 -182
rect -120 -189 -119 -187
rect -117 -189 -116 -187
rect -184 -193 -180 -190
rect -120 -191 -116 -189
rect -112 -179 -108 -173
rect -86 -169 -82 -163
rect -93 -173 -82 -169
rect -93 -179 -89 -173
rect -112 -180 -89 -179
rect -112 -182 -93 -180
rect -91 -182 -89 -180
rect -112 -183 -89 -182
rect -272 -194 -226 -193
rect -541 -195 -495 -194
rect -541 -197 -539 -195
rect -537 -197 -499 -195
rect -497 -197 -495 -195
rect -541 -198 -495 -197
rect -491 -195 -485 -194
rect -491 -197 -489 -195
rect -487 -197 -485 -195
rect -511 -202 -505 -201
rect -511 -204 -509 -202
rect -507 -204 -505 -202
rect -491 -202 -485 -197
rect -481 -195 -449 -194
rect -481 -197 -479 -195
rect -477 -197 -449 -195
rect -481 -198 -449 -197
rect -430 -195 -424 -194
rect -430 -197 -428 -195
rect -426 -197 -424 -195
rect -491 -204 -489 -202
rect -487 -204 -485 -202
rect -451 -202 -445 -201
rect -451 -204 -449 -202
rect -447 -204 -445 -202
rect -430 -204 -424 -197
rect -409 -195 -363 -194
rect -409 -197 -407 -195
rect -405 -197 -367 -195
rect -365 -197 -363 -195
rect -409 -198 -363 -197
rect -359 -195 -353 -194
rect -359 -197 -357 -195
rect -355 -197 -353 -195
rect -379 -202 -373 -201
rect -379 -204 -377 -202
rect -375 -204 -373 -202
rect -359 -202 -353 -197
rect -349 -195 -317 -194
rect -349 -197 -347 -195
rect -345 -197 -317 -195
rect -349 -198 -317 -197
rect -298 -195 -292 -194
rect -298 -197 -296 -195
rect -294 -197 -292 -195
rect -272 -196 -270 -194
rect -268 -196 -230 -194
rect -228 -196 -226 -194
rect -272 -197 -226 -196
rect -222 -194 -216 -193
rect -222 -196 -220 -194
rect -218 -196 -216 -194
rect -359 -204 -357 -202
rect -355 -204 -353 -202
rect -319 -202 -313 -201
rect -319 -204 -317 -202
rect -315 -204 -313 -202
rect -298 -204 -292 -197
rect -242 -201 -236 -200
rect -242 -203 -240 -201
rect -238 -203 -236 -201
rect -222 -201 -216 -196
rect -212 -194 -180 -193
rect -212 -196 -210 -194
rect -208 -196 -180 -194
rect -212 -197 -180 -196
rect -161 -194 -155 -193
rect -112 -194 -108 -183
rect -161 -196 -159 -194
rect -157 -196 -155 -194
rect -222 -203 -220 -201
rect -218 -203 -216 -201
rect -182 -201 -176 -200
rect -182 -203 -180 -201
rect -178 -203 -176 -201
rect -161 -203 -155 -196
rect -141 -195 -108 -194
rect -141 -197 -139 -195
rect -137 -197 -108 -195
rect -141 -198 -108 -197
rect -104 -194 -100 -192
rect -104 -196 -103 -194
rect -101 -196 -100 -194
rect -104 -201 -100 -196
rect -104 -203 -103 -201
rect -101 -203 -100 -201
rect -491 -227 -485 -220
rect -463 -221 -457 -220
rect -463 -223 -461 -221
rect -459 -223 -457 -221
rect -491 -229 -489 -227
rect -487 -229 -485 -227
rect -491 -230 -485 -229
rect -472 -227 -468 -225
rect -472 -229 -471 -227
rect -469 -229 -468 -227
rect -472 -234 -468 -229
rect -463 -228 -457 -223
rect -425 -221 -421 -220
rect -425 -223 -424 -221
rect -422 -223 -421 -221
rect -463 -230 -461 -228
rect -459 -230 -457 -228
rect -463 -231 -457 -230
rect -454 -226 -430 -225
rect -454 -228 -434 -226
rect -432 -228 -430 -226
rect -454 -229 -430 -228
rect -425 -229 -421 -223
rect -454 -234 -450 -229
rect -425 -231 -424 -229
rect -422 -231 -421 -229
rect -398 -227 -392 -220
rect -369 -221 -363 -220
rect -369 -223 -367 -221
rect -365 -223 -363 -221
rect -398 -229 -396 -227
rect -394 -229 -392 -227
rect -398 -230 -392 -229
rect -378 -227 -374 -225
rect -378 -229 -377 -227
rect -375 -229 -374 -227
rect -425 -233 -421 -231
rect -472 -236 -471 -234
rect -469 -236 -450 -234
rect -472 -238 -450 -236
rect -498 -246 -497 -239
rect -378 -234 -374 -229
rect -369 -228 -363 -223
rect -331 -221 -327 -220
rect -331 -223 -330 -221
rect -328 -223 -327 -221
rect -369 -230 -367 -228
rect -365 -230 -363 -228
rect -369 -231 -363 -230
rect -360 -226 -336 -225
rect -360 -228 -340 -226
rect -338 -228 -336 -226
rect -360 -229 -336 -228
rect -331 -229 -327 -223
rect -225 -226 -219 -219
rect -195 -220 -189 -219
rect -195 -222 -193 -220
rect -191 -222 -189 -220
rect -360 -234 -356 -229
rect -331 -231 -330 -229
rect -328 -231 -327 -229
rect -331 -233 -327 -231
rect -225 -228 -223 -226
rect -221 -228 -219 -226
rect -225 -229 -219 -228
rect -204 -226 -200 -224
rect -204 -228 -203 -226
rect -201 -228 -200 -226
rect -378 -236 -377 -234
rect -375 -236 -356 -234
rect -378 -238 -356 -236
rect -498 -264 -497 -258
rect -487 -263 -483 -261
rect -405 -246 -404 -239
rect -487 -265 -486 -263
rect -484 -265 -483 -263
rect -487 -276 -483 -265
rect -437 -266 -431 -265
rect -437 -267 -435 -266
rect -476 -268 -435 -267
rect -433 -268 -431 -266
rect -476 -270 -474 -268
rect -472 -270 -431 -268
rect -476 -271 -431 -270
rect -427 -266 -421 -265
rect -427 -268 -425 -266
rect -423 -268 -421 -266
rect -427 -276 -421 -268
rect -405 -264 -404 -258
rect -204 -233 -200 -228
rect -195 -227 -189 -222
rect -157 -220 -153 -219
rect -157 -222 -156 -220
rect -154 -222 -153 -220
rect -195 -229 -193 -227
rect -191 -229 -189 -227
rect -195 -230 -189 -229
rect -186 -225 -162 -224
rect -186 -227 -166 -225
rect -164 -227 -162 -225
rect -186 -228 -162 -227
rect -157 -228 -153 -222
rect -186 -233 -182 -228
rect -157 -230 -156 -228
rect -154 -230 -153 -228
rect -157 -232 -153 -230
rect -131 -228 -125 -219
rect -131 -230 -129 -228
rect -127 -230 -125 -228
rect -131 -231 -125 -230
rect -120 -226 -116 -224
rect -120 -228 -119 -226
rect -117 -228 -116 -226
rect -204 -235 -203 -233
rect -201 -235 -182 -233
rect -204 -237 -182 -235
rect -232 -245 -231 -238
rect -394 -263 -390 -261
rect -120 -233 -116 -228
rect -111 -226 -105 -219
rect -111 -228 -109 -226
rect -107 -228 -105 -226
rect -111 -229 -105 -228
rect -120 -234 -119 -233
rect -394 -265 -393 -263
rect -391 -265 -390 -263
rect -394 -276 -390 -265
rect -343 -266 -337 -265
rect -343 -267 -341 -266
rect -382 -268 -341 -267
rect -339 -268 -337 -266
rect -382 -270 -380 -268
rect -378 -270 -337 -268
rect -382 -271 -337 -270
rect -333 -266 -327 -265
rect -333 -268 -331 -266
rect -329 -268 -327 -266
rect -333 -276 -327 -268
rect -232 -263 -231 -257
rect -133 -235 -119 -234
rect -117 -235 -116 -233
rect -133 -238 -116 -235
rect -221 -262 -217 -260
rect -221 -264 -220 -262
rect -218 -264 -217 -262
rect -133 -250 -129 -238
rect -133 -252 -132 -250
rect -130 -252 -129 -250
rect -133 -257 -129 -252
rect -133 -261 -121 -257
rect -137 -264 -136 -262
rect -221 -275 -217 -264
rect -169 -265 -163 -264
rect -169 -266 -167 -265
rect -208 -267 -167 -266
rect -165 -267 -163 -265
rect -208 -269 -206 -267
rect -204 -269 -163 -267
rect -208 -270 -163 -269
rect -159 -265 -153 -264
rect -159 -267 -157 -265
rect -155 -267 -153 -265
rect -159 -275 -153 -267
rect -125 -265 -121 -261
rect -125 -266 -105 -265
rect -125 -268 -109 -266
rect -107 -268 -105 -266
rect -125 -269 -105 -268
rect -212 -292 -208 -291
rect -482 -293 -478 -292
rect -482 -295 -481 -293
rect -479 -295 -478 -293
rect -482 -297 -478 -295
rect -358 -293 -354 -292
rect -358 -295 -357 -293
rect -355 -295 -354 -293
rect -358 -297 -354 -295
rect -212 -294 -211 -292
rect -209 -294 -208 -292
rect -212 -296 -208 -294
rect -562 -299 -542 -298
rect -562 -301 -546 -299
rect -544 -301 -542 -299
rect -562 -302 -542 -301
rect -574 -305 -573 -303
rect -562 -306 -558 -302
rect -570 -310 -558 -306
rect -570 -315 -566 -310
rect -570 -317 -569 -315
rect -567 -317 -566 -315
rect -570 -329 -566 -317
rect -570 -332 -553 -329
rect -570 -333 -556 -332
rect -557 -334 -556 -333
rect -554 -334 -553 -332
rect -568 -337 -562 -336
rect -568 -339 -566 -337
rect -564 -339 -562 -337
rect -568 -348 -562 -339
rect -557 -339 -553 -334
rect -501 -330 -488 -329
rect -490 -332 -488 -330
rect -492 -334 -488 -332
rect -494 -337 -488 -334
rect -557 -341 -556 -339
rect -554 -341 -553 -339
rect -557 -343 -553 -341
rect -548 -339 -542 -338
rect -548 -341 -546 -339
rect -544 -341 -542 -339
rect -548 -348 -542 -341
rect -505 -339 -499 -338
rect -505 -341 -503 -339
rect -501 -341 -499 -339
rect -494 -339 -492 -337
rect -490 -339 -488 -337
rect -494 -340 -488 -339
rect -483 -330 -477 -329
rect -483 -332 -481 -330
rect -479 -332 -477 -330
rect -483 -337 -477 -332
rect -231 -329 -218 -328
rect -377 -330 -364 -329
rect -366 -332 -364 -330
rect -368 -334 -364 -332
rect -483 -339 -481 -337
rect -479 -339 -477 -337
rect -370 -337 -364 -334
rect -505 -348 -499 -341
rect -483 -348 -477 -339
rect -381 -339 -375 -338
rect -381 -341 -379 -339
rect -377 -341 -375 -339
rect -370 -339 -368 -337
rect -366 -339 -364 -337
rect -370 -340 -364 -339
rect -359 -330 -353 -329
rect -359 -332 -357 -330
rect -355 -332 -353 -330
rect -359 -337 -353 -332
rect -220 -331 -218 -329
rect -222 -333 -218 -331
rect -224 -336 -218 -333
rect -359 -339 -357 -337
rect -355 -339 -353 -337
rect -381 -348 -375 -341
rect -359 -348 -353 -339
rect -235 -338 -229 -337
rect -235 -340 -233 -338
rect -231 -340 -229 -338
rect -224 -338 -222 -336
rect -220 -338 -218 -336
rect -224 -339 -218 -338
rect -213 -329 -207 -328
rect -213 -331 -211 -329
rect -209 -331 -207 -329
rect -213 -336 -207 -331
rect -213 -338 -211 -336
rect -209 -338 -207 -336
rect -235 -347 -229 -340
rect -213 -347 -207 -338
rect -242 -363 -241 -361
rect -239 -363 -238 -361
rect -689 -365 -687 -363
rect -685 -365 -683 -363
rect -689 -366 -683 -365
rect -669 -365 -667 -363
rect -665 -365 -663 -363
rect -719 -370 -673 -369
rect -719 -372 -717 -370
rect -715 -372 -677 -370
rect -675 -372 -673 -370
rect -719 -373 -673 -372
rect -669 -370 -663 -365
rect -629 -365 -627 -363
rect -625 -365 -623 -363
rect -629 -366 -623 -365
rect -669 -372 -667 -370
rect -665 -372 -663 -370
rect -669 -373 -663 -372
rect -659 -370 -627 -369
rect -659 -372 -657 -370
rect -655 -372 -627 -370
rect -659 -373 -627 -372
rect -608 -370 -602 -363
rect -557 -365 -555 -363
rect -553 -365 -551 -363
rect -557 -366 -551 -365
rect -537 -365 -535 -363
rect -533 -365 -531 -363
rect -608 -372 -606 -370
rect -604 -372 -602 -370
rect -608 -373 -602 -372
rect -587 -370 -541 -369
rect -587 -372 -585 -370
rect -583 -372 -545 -370
rect -543 -372 -541 -370
rect -587 -373 -541 -372
rect -537 -370 -531 -365
rect -497 -365 -495 -363
rect -493 -365 -491 -363
rect -497 -366 -491 -365
rect -537 -372 -535 -370
rect -533 -372 -531 -370
rect -537 -373 -531 -372
rect -527 -370 -495 -369
rect -527 -372 -525 -370
rect -523 -372 -495 -370
rect -527 -373 -495 -372
rect -476 -370 -470 -363
rect -425 -365 -423 -363
rect -421 -365 -419 -363
rect -425 -366 -419 -365
rect -405 -365 -403 -363
rect -401 -365 -399 -363
rect -476 -372 -474 -370
rect -472 -372 -470 -370
rect -476 -373 -470 -372
rect -455 -370 -409 -369
rect -455 -372 -453 -370
rect -451 -372 -413 -370
rect -411 -372 -409 -370
rect -455 -373 -409 -372
rect -405 -370 -399 -365
rect -365 -365 -363 -363
rect -361 -365 -359 -363
rect -365 -366 -359 -365
rect -405 -372 -403 -370
rect -401 -372 -399 -370
rect -405 -373 -399 -372
rect -395 -370 -363 -369
rect -395 -372 -393 -370
rect -391 -372 -363 -370
rect -395 -373 -363 -372
rect -344 -370 -338 -363
rect -344 -372 -342 -370
rect -340 -372 -338 -370
rect -344 -373 -338 -372
rect -242 -368 -238 -363
rect -242 -370 -241 -368
rect -239 -370 -238 -368
rect -242 -372 -238 -370
rect -234 -367 -201 -366
rect -234 -369 -205 -367
rect -203 -369 -201 -367
rect -234 -370 -201 -369
rect -699 -378 -693 -377
rect -699 -380 -697 -378
rect -695 -380 -693 -378
rect -699 -384 -693 -380
rect -711 -385 -693 -384
rect -711 -387 -697 -385
rect -695 -387 -693 -385
rect -711 -388 -693 -387
rect -711 -394 -707 -388
rect -689 -393 -685 -373
rect -631 -376 -627 -373
rect -711 -396 -710 -394
rect -708 -396 -707 -394
rect -711 -401 -707 -396
rect -702 -394 -676 -393
rect -702 -396 -700 -394
rect -698 -396 -676 -394
rect -702 -397 -676 -396
rect -711 -405 -686 -401
rect -690 -409 -686 -405
rect -690 -411 -689 -409
rect -687 -411 -686 -409
rect -690 -413 -686 -411
rect -680 -408 -676 -397
rect -659 -378 -643 -377
rect -659 -380 -647 -378
rect -645 -380 -643 -378
rect -659 -381 -643 -380
rect -638 -378 -634 -376
rect -638 -380 -637 -378
rect -635 -380 -634 -378
rect -659 -393 -655 -381
rect -638 -385 -634 -380
rect -662 -394 -655 -393
rect -662 -396 -660 -394
rect -658 -396 -655 -394
rect -662 -397 -655 -396
rect -680 -409 -663 -408
rect -680 -411 -667 -409
rect -665 -411 -663 -409
rect -680 -412 -663 -411
rect -659 -409 -655 -397
rect -651 -387 -637 -385
rect -635 -387 -634 -385
rect -651 -389 -634 -387
rect -631 -378 -613 -376
rect -631 -380 -616 -378
rect -614 -380 -613 -378
rect -651 -394 -647 -389
rect -631 -393 -627 -380
rect -617 -385 -613 -380
rect -617 -389 -603 -385
rect -651 -396 -650 -394
rect -648 -396 -647 -394
rect -651 -401 -647 -396
rect -642 -394 -627 -393
rect -642 -396 -640 -394
rect -638 -396 -627 -394
rect -642 -397 -627 -396
rect -651 -405 -624 -401
rect -607 -403 -603 -389
rect -567 -378 -561 -377
rect -567 -380 -565 -378
rect -563 -380 -561 -378
rect -607 -405 -606 -403
rect -604 -405 -603 -403
rect -628 -409 -624 -405
rect -607 -407 -603 -405
rect -567 -384 -561 -380
rect -579 -385 -561 -384
rect -579 -387 -565 -385
rect -563 -387 -561 -385
rect -579 -388 -561 -387
rect -579 -394 -575 -388
rect -557 -393 -553 -373
rect -499 -376 -495 -373
rect -579 -396 -578 -394
rect -576 -396 -575 -394
rect -579 -401 -575 -396
rect -570 -394 -544 -393
rect -570 -396 -568 -394
rect -566 -396 -544 -394
rect -570 -397 -544 -396
rect -579 -405 -554 -401
rect -558 -409 -554 -405
rect -659 -410 -633 -409
rect -659 -412 -637 -410
rect -635 -412 -633 -410
rect -659 -413 -633 -412
rect -628 -411 -627 -409
rect -625 -411 -624 -409
rect -628 -413 -624 -411
rect -618 -411 -614 -409
rect -618 -413 -617 -411
rect -615 -413 -614 -411
rect -558 -411 -557 -409
rect -555 -411 -554 -409
rect -558 -413 -554 -411
rect -548 -408 -544 -397
rect -527 -378 -511 -377
rect -527 -380 -515 -378
rect -513 -380 -511 -378
rect -527 -381 -511 -380
rect -506 -378 -502 -376
rect -506 -380 -505 -378
rect -503 -380 -502 -378
rect -527 -393 -523 -381
rect -506 -385 -502 -380
rect -530 -394 -523 -393
rect -530 -396 -528 -394
rect -526 -396 -523 -394
rect -530 -397 -523 -396
rect -548 -409 -531 -408
rect -548 -411 -535 -409
rect -533 -411 -531 -409
rect -548 -412 -531 -411
rect -527 -409 -523 -397
rect -519 -387 -505 -385
rect -503 -387 -502 -385
rect -519 -389 -502 -387
rect -499 -378 -481 -376
rect -499 -380 -484 -378
rect -482 -380 -481 -378
rect -519 -394 -515 -389
rect -499 -393 -495 -380
rect -485 -385 -481 -380
rect -485 -389 -471 -385
rect -519 -396 -518 -394
rect -516 -396 -515 -394
rect -519 -401 -515 -396
rect -510 -394 -495 -393
rect -510 -396 -508 -394
rect -506 -396 -495 -394
rect -510 -397 -495 -396
rect -519 -405 -492 -401
rect -475 -403 -471 -389
rect -435 -378 -429 -377
rect -435 -380 -433 -378
rect -431 -380 -429 -378
rect -475 -405 -474 -403
rect -472 -405 -471 -403
rect -496 -409 -492 -405
rect -475 -407 -471 -405
rect -435 -384 -429 -380
rect -447 -385 -429 -384
rect -447 -387 -433 -385
rect -431 -387 -429 -385
rect -447 -388 -429 -387
rect -447 -394 -443 -388
rect -425 -393 -421 -373
rect -367 -376 -363 -373
rect -447 -396 -446 -394
rect -444 -396 -443 -394
rect -447 -401 -443 -396
rect -438 -394 -412 -393
rect -438 -396 -436 -394
rect -434 -396 -412 -394
rect -438 -397 -412 -396
rect -447 -405 -422 -401
rect -426 -409 -422 -405
rect -527 -410 -501 -409
rect -527 -412 -505 -410
rect -503 -412 -501 -410
rect -527 -413 -501 -412
rect -496 -411 -495 -409
rect -493 -411 -492 -409
rect -496 -413 -492 -411
rect -486 -411 -482 -409
rect -486 -413 -485 -411
rect -483 -413 -482 -411
rect -426 -411 -425 -409
rect -423 -411 -422 -409
rect -426 -413 -422 -411
rect -416 -408 -412 -397
rect -395 -378 -379 -377
rect -395 -380 -383 -378
rect -381 -380 -379 -378
rect -395 -381 -379 -380
rect -374 -378 -370 -376
rect -374 -380 -373 -378
rect -371 -380 -370 -378
rect -395 -393 -391 -381
rect -374 -385 -370 -380
rect -398 -394 -391 -393
rect -398 -396 -396 -394
rect -394 -396 -391 -394
rect -398 -397 -391 -396
rect -416 -409 -399 -408
rect -416 -411 -403 -409
rect -401 -411 -399 -409
rect -416 -412 -399 -411
rect -395 -409 -391 -397
rect -387 -387 -373 -385
rect -371 -387 -370 -385
rect -387 -389 -370 -387
rect -367 -378 -349 -376
rect -367 -380 -352 -378
rect -350 -380 -349 -378
rect -387 -394 -383 -389
rect -367 -393 -363 -380
rect -353 -385 -349 -380
rect -353 -389 -339 -385
rect -387 -396 -386 -394
rect -384 -396 -383 -394
rect -387 -401 -383 -396
rect -378 -394 -363 -393
rect -378 -396 -376 -394
rect -374 -396 -363 -394
rect -378 -397 -363 -396
rect -387 -405 -360 -401
rect -343 -403 -339 -389
rect -234 -381 -230 -370
rect -253 -382 -230 -381
rect -253 -384 -251 -382
rect -249 -384 -230 -382
rect -253 -385 -230 -384
rect -253 -391 -249 -385
rect -260 -395 -249 -391
rect -343 -405 -342 -403
rect -340 -405 -339 -403
rect -260 -401 -256 -395
rect -234 -391 -230 -385
rect -226 -375 -222 -373
rect -226 -377 -225 -375
rect -223 -377 -222 -375
rect -226 -382 -222 -377
rect -226 -384 -225 -382
rect -223 -383 -222 -382
rect -223 -384 -210 -383
rect -226 -387 -210 -384
rect -214 -389 -210 -387
rect -214 -391 -209 -389
rect -234 -392 -218 -391
rect -234 -394 -222 -392
rect -220 -394 -218 -392
rect -234 -395 -218 -394
rect -214 -393 -212 -391
rect -210 -393 -209 -391
rect -214 -395 -209 -393
rect -260 -403 -259 -401
rect -257 -403 -256 -401
rect -260 -405 -256 -403
rect -214 -399 -210 -395
rect -234 -403 -210 -399
rect -364 -409 -360 -405
rect -343 -407 -339 -405
rect -234 -406 -230 -403
rect -234 -408 -233 -406
rect -231 -408 -230 -406
rect -247 -409 -241 -408
rect -395 -410 -369 -409
rect -395 -412 -373 -410
rect -371 -412 -369 -410
rect -395 -413 -369 -412
rect -364 -411 -363 -409
rect -361 -411 -360 -409
rect -364 -413 -360 -411
rect -354 -411 -350 -409
rect -354 -413 -353 -411
rect -351 -413 -350 -411
rect -680 -417 -674 -416
rect -680 -419 -678 -417
rect -676 -419 -674 -417
rect -618 -419 -614 -413
rect -548 -417 -542 -416
rect -548 -419 -546 -417
rect -544 -419 -542 -417
rect -486 -419 -482 -413
rect -416 -417 -410 -416
rect -416 -419 -414 -417
rect -412 -419 -410 -417
rect -354 -419 -350 -413
rect -247 -411 -245 -409
rect -243 -411 -241 -409
rect -234 -410 -230 -408
rect -247 -417 -241 -411
rect -758 -443 -754 -441
rect -758 -445 -757 -443
rect -755 -445 -754 -443
rect -758 -448 -754 -445
rect -778 -452 -754 -448
rect -778 -456 -774 -452
rect -732 -448 -728 -446
rect -732 -450 -731 -448
rect -729 -450 -728 -448
rect -779 -458 -774 -456
rect -779 -460 -778 -458
rect -776 -460 -774 -458
rect -770 -457 -754 -456
rect -770 -459 -768 -457
rect -766 -459 -754 -457
rect -770 -460 -754 -459
rect -779 -462 -774 -460
rect -778 -464 -774 -462
rect -778 -467 -762 -464
rect -778 -468 -765 -467
rect -766 -469 -765 -468
rect -763 -469 -762 -467
rect -766 -474 -762 -469
rect -766 -476 -765 -474
rect -763 -476 -762 -474
rect -766 -478 -762 -476
rect -758 -466 -754 -460
rect -732 -456 -728 -450
rect -739 -460 -728 -456
rect -704 -445 -700 -434
rect -691 -441 -646 -440
rect -691 -443 -689 -441
rect -687 -443 -646 -441
rect -691 -444 -650 -443
rect -739 -466 -735 -460
rect -758 -470 -749 -466
rect -745 -467 -735 -466
rect -745 -469 -739 -467
rect -737 -469 -735 -467
rect -745 -470 -735 -469
rect -758 -481 -754 -470
rect -715 -452 -714 -446
rect -704 -447 -703 -445
rect -701 -447 -700 -445
rect -652 -445 -650 -444
rect -648 -445 -646 -443
rect -652 -446 -646 -445
rect -642 -443 -636 -435
rect -642 -445 -640 -443
rect -638 -445 -636 -443
rect -642 -446 -636 -445
rect -704 -449 -700 -447
rect -572 -446 -568 -435
rect -559 -441 -514 -440
rect -559 -443 -557 -441
rect -555 -443 -514 -441
rect -559 -444 -518 -443
rect -520 -445 -518 -444
rect -516 -445 -514 -443
rect -520 -446 -514 -445
rect -510 -443 -504 -435
rect -510 -445 -508 -443
rect -506 -445 -504 -443
rect -510 -446 -504 -445
rect -715 -471 -714 -464
rect -687 -475 -665 -473
rect -687 -477 -686 -475
rect -684 -477 -665 -475
rect -787 -482 -754 -481
rect -787 -484 -785 -482
rect -783 -484 -754 -482
rect -787 -485 -754 -484
rect -750 -490 -749 -479
rect -708 -481 -702 -480
rect -708 -483 -706 -481
rect -704 -483 -702 -481
rect -708 -490 -702 -483
rect -687 -482 -683 -477
rect -687 -484 -686 -482
rect -684 -484 -683 -482
rect -687 -486 -683 -484
rect -678 -481 -672 -480
rect -678 -483 -676 -481
rect -674 -483 -672 -481
rect -678 -488 -672 -483
rect -669 -482 -665 -477
rect -583 -453 -582 -447
rect -572 -448 -571 -446
rect -569 -448 -568 -446
rect -440 -445 -436 -434
rect -430 -440 -385 -439
rect -430 -442 -428 -440
rect -426 -442 -385 -440
rect -430 -443 -389 -442
rect -391 -444 -389 -443
rect -387 -444 -385 -442
rect -391 -445 -385 -444
rect -381 -442 -375 -434
rect -381 -444 -379 -442
rect -377 -444 -375 -442
rect -381 -445 -375 -444
rect -245 -439 -225 -438
rect -245 -441 -229 -439
rect -227 -441 -225 -439
rect -245 -442 -225 -441
rect -572 -450 -568 -448
rect -583 -472 -582 -465
rect -555 -475 -533 -473
rect -555 -477 -554 -475
rect -552 -477 -533 -475
rect -640 -480 -636 -478
rect -640 -482 -639 -480
rect -637 -482 -636 -480
rect -669 -483 -645 -482
rect -669 -485 -649 -483
rect -647 -485 -645 -483
rect -669 -486 -645 -485
rect -678 -490 -676 -488
rect -674 -490 -672 -488
rect -678 -491 -672 -490
rect -640 -488 -636 -482
rect -640 -490 -639 -488
rect -637 -490 -636 -488
rect -640 -491 -636 -490
rect -576 -482 -570 -481
rect -576 -484 -574 -482
rect -572 -484 -570 -482
rect -576 -491 -570 -484
rect -555 -482 -551 -477
rect -555 -484 -554 -482
rect -552 -484 -551 -482
rect -555 -486 -551 -484
rect -546 -481 -540 -480
rect -546 -483 -544 -481
rect -542 -483 -540 -481
rect -546 -488 -540 -483
rect -537 -482 -533 -477
rect -451 -452 -450 -446
rect -440 -447 -439 -445
rect -437 -447 -436 -445
rect -440 -449 -436 -447
rect -451 -471 -450 -464
rect -426 -474 -404 -472
rect -426 -476 -425 -474
rect -423 -476 -404 -474
rect -508 -480 -504 -478
rect -508 -482 -507 -480
rect -505 -482 -504 -480
rect -537 -483 -513 -482
rect -537 -485 -517 -483
rect -515 -485 -513 -483
rect -537 -486 -513 -485
rect -546 -490 -544 -488
rect -542 -490 -540 -488
rect -546 -491 -540 -490
rect -508 -488 -504 -482
rect -508 -490 -507 -488
rect -505 -490 -504 -488
rect -444 -481 -438 -480
rect -444 -483 -442 -481
rect -440 -483 -438 -481
rect -444 -490 -438 -483
rect -426 -481 -422 -476
rect -426 -483 -425 -481
rect -423 -483 -422 -481
rect -426 -485 -422 -483
rect -417 -480 -411 -479
rect -417 -482 -415 -480
rect -413 -482 -411 -480
rect -417 -487 -411 -482
rect -408 -481 -404 -476
rect -257 -445 -256 -443
rect -245 -446 -241 -442
rect -253 -450 -241 -446
rect -253 -455 -249 -450
rect -253 -457 -252 -455
rect -250 -457 -249 -455
rect -253 -469 -249 -457
rect -253 -472 -236 -469
rect -253 -473 -239 -472
rect -240 -474 -239 -473
rect -237 -474 -236 -472
rect -251 -477 -245 -476
rect -379 -479 -375 -477
rect -379 -481 -378 -479
rect -376 -481 -375 -479
rect -408 -482 -384 -481
rect -408 -484 -388 -482
rect -386 -484 -384 -482
rect -408 -485 -384 -484
rect -417 -489 -415 -487
rect -413 -489 -411 -487
rect -417 -490 -411 -489
rect -379 -487 -375 -481
rect -379 -489 -378 -487
rect -376 -489 -375 -487
rect -251 -479 -249 -477
rect -247 -479 -245 -477
rect -251 -488 -245 -479
rect -240 -479 -236 -474
rect -240 -481 -239 -479
rect -237 -481 -236 -479
rect -240 -483 -236 -481
rect -231 -479 -225 -478
rect -231 -481 -229 -479
rect -227 -481 -225 -479
rect -231 -488 -225 -481
rect -379 -490 -375 -489
rect -508 -491 -504 -490
<< via1 >>
rect 168 143 170 145
rect -265 124 -263 126
rect -272 108 -270 110
rect -199 124 -197 126
rect -283 100 -281 102
rect -243 101 -241 103
rect -155 116 -153 118
rect -191 99 -189 101
rect -103 124 -101 126
rect -96 108 -94 110
rect -59 124 -57 126
rect -84 101 -82 103
rect -40 110 -38 112
rect -16 125 -14 127
rect -52 98 -50 100
rect 13 112 15 114
rect -8 108 -6 110
rect 37 125 39 127
rect 45 99 47 101
rect 57 110 59 112
rect 82 125 84 127
rect 80 108 82 110
rect 125 125 127 127
rect 132 99 134 101
rect -347 73 -345 75
rect -377 71 -375 73
rect 13 61 15 63
rect -347 50 -345 52
rect -387 21 -385 23
rect -283 36 -281 38
rect -267 35 -265 37
rect -216 50 -214 52
rect -245 20 -243 22
rect -153 37 -151 39
rect -136 36 -134 38
rect -83 50 -81 52
rect -110 20 -108 22
rect -25 37 -23 39
rect -4 35 -2 37
rect 25 37 27 39
rect 63 6 65 8
rect -283 -10 -281 -8
rect -364 -26 -362 -24
rect -335 -27 -333 -25
rect -351 -36 -349 -34
rect -320 -27 -318 -25
rect -239 -18 -237 -16
rect -189 -19 -187 -17
rect -267 -26 -265 -24
rect -255 -27 -253 -25
rect -404 -43 -402 -41
rect -200 -29 -198 -27
rect 0 -16 2 -14
rect -150 -29 -148 -27
rect -122 -19 -120 -17
rect -135 -27 -133 -25
rect -122 -28 -120 -26
rect -59 -29 -57 -27
rect 25 -28 27 -26
rect 42 -36 44 -34
rect -320 -61 -318 -59
rect -442 -71 -440 -69
rect -508 -108 -506 -106
rect -472 -108 -470 -106
rect -449 -126 -447 -124
rect -371 -100 -369 -98
rect -277 -92 -275 -90
rect -397 -108 -395 -106
rect -258 -92 -256 -90
rect -229 -92 -227 -90
rect -286 -99 -284 -97
rect -126 -92 -124 -90
rect -305 -123 -303 -121
rect -285 -115 -283 -113
rect -158 -111 -156 -109
rect -82 -92 -80 -90
rect -133 -108 -131 -106
rect 130 -108 132 -106
rect 151 -108 153 -106
rect -114 -119 -112 -117
rect -90 -117 -88 -115
rect -82 -139 -80 -137
rect 151 -137 153 -135
rect -492 -170 -490 -168
rect -540 -187 -538 -185
rect -438 -173 -436 -171
rect -420 -189 -418 -187
rect -360 -172 -358 -170
rect -408 -189 -406 -187
rect -305 -167 -303 -165
rect -288 -190 -286 -188
rect -223 -171 -221 -169
rect -271 -188 -269 -186
rect -167 -165 -165 -163
rect -151 -188 -149 -186
rect -100 -163 -98 -161
rect -84 -183 -82 -181
rect -517 -210 -515 -208
rect -475 -244 -473 -242
rect -435 -238 -433 -236
rect -404 -237 -402 -235
rect -271 -231 -269 -229
rect -568 -255 -566 -253
rect -485 -254 -483 -252
rect -459 -253 -457 -251
rect -444 -253 -442 -251
rect -381 -245 -379 -243
rect -333 -245 -331 -243
rect -400 -262 -398 -260
rect -342 -253 -340 -251
rect -271 -257 -269 -255
rect -235 -246 -233 -244
rect -207 -244 -205 -242
rect -364 -262 -362 -260
rect -140 -238 -138 -236
rect -158 -244 -156 -242
rect -227 -261 -225 -259
rect -168 -252 -166 -250
rect -108 -237 -106 -235
rect -190 -261 -188 -259
rect -125 -252 -123 -250
rect -113 -278 -111 -276
rect -284 -287 -282 -285
rect -259 -287 -257 -285
rect 133 -287 135 -285
rect 159 -287 161 -285
rect -577 -321 -575 -319
rect -552 -309 -550 -307
rect -531 -324 -529 -322
rect -286 -299 -284 -297
rect -258 -299 -256 -297
rect -364 -303 -362 -301
rect -480 -308 -478 -306
rect -488 -323 -486 -321
rect -503 -333 -501 -331
rect -286 -320 -284 -318
rect -248 -320 -246 -318
rect -363 -323 -361 -321
rect 134 -299 136 -297
rect 151 -299 153 -297
rect -210 -307 -208 -305
rect -225 -320 -223 -318
rect -371 -333 -369 -331
rect -234 -332 -232 -330
rect -709 -359 -707 -357
rect -260 -370 -258 -368
rect -670 -381 -668 -379
rect -615 -396 -613 -394
rect -598 -397 -596 -395
rect -538 -382 -536 -380
rect -484 -396 -482 -394
rect -466 -396 -464 -394
rect -406 -380 -404 -378
rect -355 -397 -353 -395
rect -334 -397 -332 -395
rect -244 -393 -242 -391
rect -208 -423 -206 -421
rect -747 -460 -745 -458
rect -586 -444 -584 -442
rect -642 -452 -640 -450
rect -702 -458 -700 -456
rect -686 -460 -684 -458
rect -659 -473 -657 -471
rect -642 -469 -640 -467
rect -259 -440 -257 -438
rect -514 -452 -512 -450
rect -572 -460 -570 -458
rect -554 -460 -552 -458
rect -542 -468 -540 -466
rect -380 -451 -378 -449
rect -439 -458 -437 -456
rect -428 -459 -426 -457
rect -518 -475 -516 -473
rect -397 -471 -395 -469
rect -450 -475 -448 -473
rect -381 -468 -379 -466
rect -236 -450 -234 -448
rect -228 -465 -226 -463
rect -776 -496 -774 -494
rect -748 -496 -746 -494
<< via2 >>
rect -389 71 -387 73
rect -260 108 -258 110
rect -180 99 -178 101
rect -350 36 -348 38
rect -720 -360 -718 -358
rect -451 -73 -449 -71
rect -397 -75 -395 -73
rect -351 -44 -349 -42
rect -245 10 -243 12
rect -92 108 -90 110
rect -24 112 -22 114
rect -3 109 -1 111
rect -47 99 -45 101
rect -105 12 -103 14
rect -136 -1 -134 1
rect -128 -19 -126 -17
rect 74 109 76 111
rect -166 -29 -164 -27
rect -131 -27 -129 -25
rect 49 99 51 101
rect 67 8 69 10
rect -365 -76 -363 -74
rect -245 -71 -243 -69
rect -787 -496 -785 -494
rect -525 -210 -523 -208
rect -258 -116 -256 -114
rect 143 -116 145 -114
rect 181 144 183 146
rect -19 -125 -17 -123
rect -105 -134 -103 -132
rect -82 -145 -80 -143
rect 143 -139 145 -137
rect -404 -287 -402 -285
rect -405 -323 -403 -321
rect -360 -287 -358 -285
rect -379 -323 -377 -321
rect -106 -278 -104 -276
rect -201 -423 -199 -421
<< via3 >>
rect -181 -125 -179 -123
rect -57 -125 -55 -123
<< labels >>
rlabel alu1 37 9 37 9 6 vss
rlabel alu1 37 73 37 73 6 vdd
rlabel alu1 27 -63 27 -63 8 vdd
rlabel alu1 27 1 27 1 8 vss
rlabel alu0 10 32 10 32 1 r3t1
rlabel alu0 26 47 26 47 1 r3t1
rlabel alu0 42 37 42 37 1 r3t1
rlabel alu0 50 62 50 62 1 r3t1
rlabel alu0 44 50 44 50 1 r3t11
rlabel alu1 57 53 57 53 1 Z1
rlabel alu1 65 41 65 41 1 Z1
rlabel alu1 9 53 9 53 1 X1Y0
rlabel alu1 17 61 17 61 1 X1Y0
rlabel alu1 17 29 17 29 1 X0Y1
rlabel polyct1 25 33 25 33 1 X0Y1
rlabel alu0 56 37 56 37 1 r3t11
rlabel alu0 36 25 36 25 1 r3t11
rlabel alu1 49 21 49 21 1 Z1
rlabel alu1 57 21 57 21 1 Z1
rlabel alu1 11 -27 11 -27 1 c1
rlabel alu1 19 -11 19 -11 1 c1
rlabel alu0 19 -30 19 -30 1 r4t1
rlabel alu0 32 -47 32 -47 1 r4t1
rlabel alu1 30 145 30 145 8 vss
rlabel alu1 30 81 30 81 8 vdd
rlabel alu1 38 121 38 121 1 X1
rlabel alu1 46 101 46 101 1 Y0
rlabel alu1 14 117 14 117 1 X1Y0
rlabel alu1 22 133 22 133 1 X1Y0
rlabel alu0 22 114 22 114 1 r2t1
rlabel alu0 38 133 38 133 1 r2t1
rlabel alu1 74 145 74 145 8 vss
rlabel alu1 74 81 74 81 8 vdd
rlabel alu1 27 -27 27 -27 1 X1Y0
rlabel alu1 35 -23 35 -23 1 X1Y0
rlabel alu1 35 -35 35 -35 1 X0Y1
rlabel alu1 43 -43 43 -43 1 X0Y1
rlabel alu1 58 117 58 117 1 X0Y1
rlabel alu1 66 133 66 133 1 X0Y1
rlabel alu1 74 117 74 117 1 X0
rlabel alu1 82 121 82 121 1 X0
rlabel alu1 82 109 82 109 1 Y1
rlabel alu0 66 114 66 114 1 r2t2
rlabel alu0 79 97 79 97 1 r2t2
rlabel alu0 82 133 82 133 1 r2t2
rlabel alu1 117 145 117 145 8 vss
rlabel alu1 117 81 117 81 8 vdd
rlabel alu1 101 117 101 117 1 Z0
rlabel alu1 117 117 117 117 1 X0
rlabel alu1 125 121 125 121 1 X0
rlabel alu1 125 109 125 109 1 Y0
rlabel alu1 133 101 133 101 1 Y0
rlabel alu0 109 114 109 114 1 r2t3
rlabel alu0 122 97 122 97 1 r2t3
rlabel alu1 109 133 109 133 1 Z0
rlabel alu0 125 133 125 133 1 r2t3
rlabel alu1 -63 73 -63 73 6 vdd
rlabel alu1 -11 53 -11 53 1 c1
rlabel polyct1 -3 45 -3 45 1 c1
rlabel alu0 35 -11 35 -11 1 r4t1
rlabel alu0 -11 36 -11 36 1 r3t2
rlabel alu0 -21 49 -21 49 1 r3t2
rlabel alu0 -41 37 -41 37 1 r3t2
rlabel alu0 -49 61 -49 61 1 r3t2
rlabel alu0 -42 49 -42 49 1 r3t22
rlabel polyct0 -55 37 -55 37 1 r3t22
rlabel alu0 -32 25 -32 25 1 r3t22
rlabel alu0 -93 49 -93 49 1 r3t222
rlabel alu0 -102 61 -102 61 1 r3t222
rlabel alu1 -115 53 -115 53 1 z2t1
rlabel alu1 -115 21 -115 21 1 z2t1
rlabel alu1 -107 21 -107 21 1 z2t1
rlabel alu1 -83 53 -83 53 1 X2Y0
rlabel alu1 -75 41 -75 41 1 X2Y0
rlabel alu1 -67 80 -67 80 8 vdd
rlabel alu1 -67 144 -67 144 8 vss
rlabel alu1 -83 116 -83 116 1 X2Y0
rlabel alu1 -75 132 -75 132 1 X2Y0
rlabel alu0 -75 113 -75 113 1 r2t4
rlabel alu0 -59 132 -59 132 1 r2t4
rlabel alu0 -62 96 -62 96 1 r2t4
rlabel alu1 -51 100 -51 100 1 Y0
rlabel alu1 -59 108 -59 108 1 Y0
rlabel alu1 -67 116 -67 116 1 X2
rlabel alu1 -59 120 -59 120 1 X2
rlabel polyct1 -27 37 -27 37 1 X1Y1
rlabel alu1 -19 33 -19 33 1 X1Y1
rlabel alu1 -23 145 -23 145 8 vss
rlabel alu1 -23 81 -23 81 8 vdd
rlabel alu1 -39 117 -39 117 1 X1Y1
rlabel alu1 -31 133 -31 133 1 X1Y1
rlabel alu0 -31 114 -31 114 1 r2t5
rlabel alu0 -15 133 -15 133 1 r2t5
rlabel alu1 -23 117 -23 117 1 X1
rlabel alu1 -15 121 -15 121 1 X1
rlabel alu1 -15 109 -15 109 1 Y1
rlabel alu0 -78 22 -78 22 1 r3t222
rlabel alu1 -63 9 -63 9 6 vss
rlabel alu1 -94 -63 -94 -63 8 vdd
rlabel alu1 -94 1 -94 1 8 vss
rlabel alu1 -122 -31 -122 -31 1 X2Y0
rlabel polyct1 -114 -27 -114 -27 1 X2Y0
rlabel alu1 -74 -19 -74 -19 1 c1
rlabel alu1 -74 -31 -74 -31 1 X1Y1
rlabel alu1 -82 -43 -82 -43 1 X1Y1
rlabel alu0 -90 -52 -90 -52 1 r4t2
rlabel alu0 -118 -47 -118 -47 1 r4t2
rlabel alu0 -102 -10 -102 -10 1 r4t22
rlabel alu1 -123 37 -123 37 1 z2t1
rlabel alu1 -195 9 -195 9 6 vss
rlabel alu1 -195 73 -195 73 6 vdd
rlabel alu1 -143 53 -143 53 1 c2
rlabel polyct1 -135 45 -135 45 1 c2
rlabel alu0 -153 49 -153 49 1 r3t3
rlabel alu0 -143 36 -143 36 1 r3t3
rlabel polyct1 -159 37 -159 37 1 X2Y1
rlabel alu1 -151 33 -151 33 1 X2Y1
rlabel alu0 -173 37 -173 37 1 r3t3
rlabel alu0 -164 25 -164 25 1 r3t33
rlabel polyct0 -187 37 -187 37 1 r3t33
rlabel alu0 -174 49 -174 49 1 r3t33
rlabel alu0 -181 61 -181 61 1 r3t3
rlabel alu0 -225 49 -225 49 1 r3t333
rlabel alu0 -234 61 -234 61 1 r3t333
rlabel alu0 -210 22 -210 22 1 r3t333
rlabel alu1 -247 53 -247 53 1 z2t2
rlabel alu1 -255 37 -255 37 1 z2t2
rlabel alu1 -247 21 -247 21 1 z2t2
rlabel alu1 -239 21 -239 21 1 z2t2
rlabel alu1 -111 81 -111 81 8 vdd
rlabel alu1 -127 117 -127 117 1 X2Y1
rlabel alu1 -119 133 -119 133 1 X2Y1
rlabel alu0 -119 114 -119 114 1 r2t6
rlabel alu0 -106 97 -106 97 1 r2t6
rlabel alu0 -103 133 -103 133 1 r2t6
rlabel alu1 -111 117 -111 117 1 X2
rlabel alu1 -103 121 -103 121 1 X2
rlabel alu1 -103 109 -103 109 1 Y1
rlabel alu1 -111 145 -111 145 8 vss
rlabel alu1 -206 81 -206 81 8 vdd
rlabel alu1 -206 145 -206 145 8 vss
rlabel alu1 -222 117 -222 117 1 X3Y0
rlabel alu1 -214 133 -214 133 1 X3Y0
rlabel alu0 -214 114 -214 114 1 r2t7
rlabel alu0 -201 97 -201 97 1 r2t7
rlabel alu0 -198 133 -198 133 1 r2t7
rlabel alu1 -206 117 -206 117 1 X3
rlabel alu1 -198 121 -198 121 1 X3
rlabel alu1 -198 109 -198 109 1 Y0
rlabel alu1 -190 101 -190 101 1 Y0
rlabel alu1 -242 145 -242 145 8 vss
rlabel alu1 -242 81 -242 81 8 vdd
rlabel alu1 -234 117 -234 117 5 X3Y0
rlabel alu1 -242 121 -242 121 5 X3Y0
rlabel alu1 -242 101 -242 101 5 X3Y0inv
rlabel alu1 -250 117 -250 117 5 X3Y0inv
rlabel alu1 -215 53 -215 53 1 X3Y0inv
rlabel alu1 -207 41 -207 41 1 X3Y0inv
rlabel alu1 -226 2 -226 2 8 vss
rlabel alu1 -226 -62 -226 -62 8 vdd
rlabel alu1 -254 -30 -254 -30 1 X3Y0inv
rlabel polyct1 -246 -26 -246 -26 1 X3Y0inv
rlabel alu0 -222 -51 -222 -51 1 r4t3
rlabel alu0 -250 -46 -250 -46 1 r4t3
rlabel alu0 -234 -9 -234 -9 1 r4t33
rlabel alu0 -214 -10 -214 -10 1 r4t33
rlabel alu1 -214 -42 -214 -42 1 c2
rlabel alu1 -206 -30 -206 -30 1 c2
rlabel alu1 -206 -18 -206 -18 1 X2Y1
rlabel alu1 -214 -18 -214 -18 1 X2Y1
rlabel alu1 -222 -26 -222 -26 1 X2Y1
rlabel alu0 -341 22 -341 22 1 r3t444
rlabel alu0 -356 49 -356 49 1 r3t444
rlabel alu0 -365 61 -365 61 1 r3t444
rlabel alu0 -295 25 -295 25 1 r3t44
rlabel polyct0 -318 37 -318 37 1 r3t44
rlabel alu0 -305 49 -305 49 1 r3t44
rlabel alu0 -312 61 -312 61 1 r3t4
rlabel alu0 -274 36 -274 36 1 r3t4
rlabel alu0 -284 49 -284 49 1 r3t4
rlabel alu1 -370 21 -370 21 1 z2t3
rlabel alu1 -378 21 -378 21 1 z2t3
rlabel alu1 -386 37 -386 37 1 z2t3
rlabel alu1 -378 53 -378 53 1 z2t3
rlabel alu1 -338 41 -338 41 1 vdd
rlabel alu1 -346 53 -346 53 1 vdd
rlabel alu1 -282 33 -282 33 1 X3Y1inv
rlabel polyct1 -290 37 -290 37 1 X3Y1inv
rlabel polyct1 -266 45 -266 45 1 c3
rlabel alu1 -274 53 -274 53 1 c3
rlabel alu1 -326 73 -326 73 6 vdd
rlabel alu1 -326 9 -326 9 6 vss
rlabel alu1 -286 121 -286 121 5 X3Y1inv
rlabel alu1 -278 101 -278 101 5 X3Y1inv
rlabel alu1 -262 125 -262 125 5 X3
rlabel alu1 -270 129 -270 129 5 X3
rlabel polyct1 -278 117 -278 117 5 Y1
rlabel alu1 -270 109 -270 109 5 Y1
rlabel alu1 -274 81 -274 81 8 vdd
rlabel alu1 -274 145 -274 145 8 vss
rlabel alu1 -141 1 -141 1 8 vss
rlabel alu1 -141 -63 -141 -63 8 vdd
rlabel alu1 -133 -27 -133 -27 5 c2inv
rlabel alu1 -141 -23 -141 -23 5 c2inv
rlabel alu1 -141 -43 -141 -43 5 c2
rlabel alu1 -149 -27 -149 -27 5 c2
rlabel alu1 -106 -23 -106 -23 1 c2inv
rlabel alu1 -98 -35 -98 -35 1 c2inv
rlabel alu1 -98 -19 -98 -19 1 c2inv
rlabel pdifct1 -90 -43 -90 -43 1 c2inv
rlabel alu1 -282 -26 -282 -26 5 c3
rlabel alu1 -274 -42 -274 -42 5 c3
rlabel alu1 -274 -22 -274 -22 5 c3inv
rlabel alu1 -266 -26 -266 -26 5 c3inv
rlabel alu1 -274 -62 -274 -62 8 vdd
rlabel alu1 -274 2 -274 2 8 vss
rlabel alu1 -230 -18 -230 -18 1 c3inv
rlabel alu1 -238 -22 -238 -22 1 c3inv
rlabel alu1 -230 -34 -230 -34 1 c3inv
rlabel pdifct1 -222 -42 -222 -42 1 c3inv
rlabel alu1 -376 -26 -376 -26 5 c4
rlabel alu1 -368 -42 -368 -42 5 c4
rlabel alu1 -368 -22 -368 -22 5 c4inv
rlabel alu1 -360 -26 -360 -26 5 c4inv
rlabel alu1 -368 -62 -368 -62 8 vdd
rlabel alu1 -368 2 -368 2 8 vss
rlabel alu0 -310 -10 -310 -10 5 r4t44
rlabel alu0 -330 -9 -330 -9 5 r4t44
rlabel alu0 -346 -46 -346 -46 5 r4t4
rlabel alu1 -326 -18 -326 -18 5 c4inv
rlabel alu1 -334 -22 -334 -22 5 c4inv
rlabel alu1 -326 -34 -326 -34 5 c4inv
rlabel alu1 -350 -30 -350 -30 5 X3Y1inv
rlabel polyct1 -342 -26 -342 -26 5 X3Y1inv
rlabel alu1 -302 -18 -302 -18 5 vdd
rlabel alu1 -310 -18 -310 -18 5 vdd
rlabel alu1 -302 -30 -302 -30 5 c3
rlabel alu1 -310 -42 -310 -42 5 c3
rlabel alu1 -322 -62 -322 -62 8 vdd
rlabel alu1 -322 2 -322 2 8 vss
rlabel alu1 -97 -135 -97 -135 6 vss
rlabel alu1 -97 -71 -97 -71 6 vdd
rlabel alu1 -89 -111 -89 -111 1 X0
rlabel alu1 -97 -107 -97 -107 1 X0
rlabel alu0 -105 -104 -105 -104 1 r5t1
rlabel alu0 -92 -87 -92 -87 1 r5t1
rlabel alu1 -113 -107 -113 -107 1 X0Y2
rlabel alu1 -105 -123 -105 -123 1 X0Y2
rlabel via1 -81 -91 -81 -91 1 Y2
rlabel alu1 -89 -99 -89 -99 1 Y2
rlabel alu0 -89 -123 -89 -123 1 r5t1
rlabel alu1 -91 -195 -91 -195 1 X0Y2
rlabel alu1 -83 -187 -83 -187 1 X0Y2
rlabel alu0 -84 -166 -84 -166 1 r6t11
rlabel alu1 -91 -163 -91 -163 1 z2t1
rlabel polyct1 -99 -167 -99 -167 1 z2t1
rlabel alu0 -100 -181 -100 -181 1 r6t11
rlabel alu0 -124 -196 -124 -196 1 r6t11
rlabel alu0 -118 -184 -118 -184 1 r6t1
rlabel alu0 -116 -171 -116 -171 1 r6t11
rlabel alu0 -130 -171 -130 -171 1 r6t1
rlabel alu0 -110 -159 -110 -159 1 r6t1
rlabel alu1 -111 -207 -111 -207 2 vdd
rlabel alu1 -111 -143 -111 -143 2 vss
rlabel alu1 -139 -175 -139 -175 1 Z2
rlabel alu1 -131 -155 -131 -155 1 Z2
rlabel alu1 -131 -187 -131 -187 1 Z2
rlabel alu1 -123 -279 -123 -279 6 vss
rlabel alu1 -123 -215 -123 -215 6 vdd
rlabel alu1 -107 -235 -107 -235 1 z2t1
rlabel alu1 -115 -243 -115 -243 1 z2t1
rlabel alu1 -123 -251 -123 -251 1 X0Y2
rlabel alu1 -115 -255 -115 -255 1 X0Y2
rlabel alu0 -131 -248 -131 -248 1 r7t1
rlabel alu0 -118 -231 -118 -231 1 r7t1
rlabel alu1 -139 -251 -139 -251 1 c5
rlabel alu1 -131 -267 -131 -267 1 c5
rlabel alu1 -210 -143 -210 -143 8 vss
rlabel alu1 -210 -207 -210 -207 8 vdd
rlabel alu1 -158 -187 -158 -187 5 c5
rlabel polyct1 -150 -179 -150 -179 5 c5
rlabel alu1 -166 -167 -166 -167 5 X1Y2
rlabel polyct1 -174 -171 -174 -171 5 X1Y2
rlabel alu1 -230 -187 -230 -187 5 z2t2
rlabel alu1 -222 -175 -222 -175 5 z2t2
rlabel alu1 -262 -187 -262 -187 5 z3t1
rlabel alu1 -270 -171 -270 -171 5 z3t1
rlabel alu1 -262 -155 -262 -155 5 z3t1
rlabel alu1 -254 -155 -254 -155 5 z3t1
rlabel alu0 -249 -195 -249 -195 5 r6t2
rlabel alu0 -240 -183 -240 -183 5 r6t2
rlabel alu0 -225 -156 -225 -156 5 r6t2
rlabel polyct0 -202 -171 -202 -171 5 r6t22
rlabel alu0 -189 -183 -189 -183 5 r6t22
rlabel alu0 -179 -159 -179 -159 5 r6t22
rlabel alu0 -158 -170 -158 -170 5 r6t222
rlabel alu0 -168 -183 -168 -183 5 r6t222
rlabel alu1 -141 -135 -141 -135 6 vss
rlabel alu1 -141 -71 -141 -71 6 vdd
rlabel via1 -125 -91 -125 -91 1 Y2
rlabel alu1 -133 -99 -133 -99 1 Y2
rlabel alu1 -141 -107 -141 -107 1 X1
rlabel alu1 -133 -111 -133 -111 1 X1
rlabel alu0 -136 -87 -136 -87 1 r5t2
rlabel alu0 -149 -104 -149 -104 1 r5t2
rlabel alu0 -133 -123 -133 -123 1 r5t2
rlabel alu1 -157 -107 -157 -107 1 X1Y2
rlabel alu1 -149 -123 -149 -123 1 X1Y2
rlabel alu0 -196 -195 -196 -195 5 r6t222
rlabel alu1 -178 -279 -178 -279 6 vss
rlabel alu1 -178 -215 -178 -215 6 vdd
rlabel alu1 -182 -243 -182 -243 1 c6inv
rlabel pdifct1 -174 -235 -174 -235 1 c6inv
rlabel alu1 -190 -255 -190 -255 1 c6inv
rlabel alu1 -182 -259 -182 -259 1 c6inv
rlabel alu0 -174 -226 -174 -226 1 r7t2
rlabel alu0 -202 -231 -202 -231 1 r7t2
rlabel alu0 -186 -268 -186 -268 1 r7t22
rlabel alu0 -166 -267 -166 -267 1 r7t22
rlabel alu1 -166 -235 -166 -235 1 c5
rlabel alu1 -158 -247 -158 -247 1 c5
rlabel alu1 -206 -247 -206 -247 1 z2t2
rlabel polyct1 -198 -251 -198 -251 1 z2t2
rlabel alu1 -174 -251 -174 -251 1 X1Y2
rlabel alu1 -166 -259 -166 -259 1 X1Y2
rlabel alu1 -158 -259 -158 -259 1 X1Y2
rlabel alu1 -218 -251 -218 -251 1 c6inv
rlabel alu1 -226 -255 -226 -255 1 c6inv
rlabel alu1 -226 -235 -226 -235 1 c6
rlabel alu1 -234 -251 -234 -251 1 c6
rlabel alu1 -226 -215 -226 -215 6 vdd
rlabel alu1 -226 -279 -226 -279 6 vss
rlabel alu1 -300 -122 -300 -122 1 X2Y2
rlabel alu1 -308 -106 -308 -106 1 X2Y2
rlabel alu0 -284 -122 -284 -122 1 r5t3
rlabel alu0 -287 -86 -287 -86 1 r5t3
rlabel alu0 -300 -103 -300 -103 1 r5t3
rlabel alu1 -276 -90 -276 -90 1 Y2
rlabel alu1 -284 -98 -284 -98 1 Y2
rlabel alu1 -284 -110 -284 -110 1 X2
rlabel alu1 -292 -106 -292 -106 1 X2
rlabel alu1 -292 -70 -292 -70 6 vdd
rlabel alu1 -292 -134 -292 -134 6 vss
rlabel alu1 -347 -144 -347 -144 8 vss
rlabel alu1 -347 -208 -347 -208 8 vdd
rlabel alu1 -295 -188 -295 -188 5 c6
rlabel polyct1 -287 -180 -287 -180 5 c6
rlabel alu0 -305 -184 -305 -184 5 r6t3
rlabel alu0 -295 -171 -295 -171 5 r6t3
rlabel alu0 -325 -172 -325 -172 5 r6t3
rlabel alu0 -333 -196 -333 -196 5 r6t3
rlabel alu0 -326 -184 -326 -184 5 r6t33
rlabel polyct0 -339 -172 -339 -172 5 r6t33
rlabel alu0 -316 -160 -316 -160 5 r6t33
rlabel polyct1 -311 -172 -311 -172 5 X2Y2
rlabel alu1 -303 -168 -303 -168 5 X2Y2
rlabel alu0 -386 -196 -386 -196 5 r6t333
rlabel alu0 -377 -184 -377 -184 5 r6t333
rlabel alu0 -362 -157 -362 -157 5 r6t333
rlabel alu1 -367 -188 -367 -188 5 z2t3
rlabel alu1 -359 -176 -359 -176 5 z2t3
rlabel alu1 -399 -188 -399 -188 5 z3t2
rlabel alu1 -407 -172 -407 -172 5 z3t2
rlabel alu1 -399 -156 -399 -156 5 z3t2
rlabel alu1 -391 -156 -391 -156 5 z3t2
rlabel alu1 -352 -280 -352 -280 6 vss
rlabel alu1 -352 -216 -352 -216 6 vdd
rlabel alu1 -340 -236 -340 -236 1 c6
rlabel alu1 -332 -248 -332 -248 1 c6
rlabel pdifct1 -348 -236 -348 -236 1 c7inv
rlabel alu1 -356 -244 -356 -244 1 c7inv
rlabel alu1 -364 -256 -364 -256 1 c7inv
rlabel alu1 -356 -260 -356 -260 1 c7inv
rlabel alu1 -348 -252 -348 -252 1 X2Y2
rlabel alu1 -340 -260 -340 -260 1 X2Y2
rlabel alu1 -332 -260 -332 -260 1 X2Y2
rlabel alu0 -340 -268 -340 -268 1 r7t3
rlabel alu0 -360 -269 -360 -269 1 r7t3
rlabel alu0 -376 -232 -376 -232 1 r7t33
rlabel alu0 -348 -227 -348 -227 1 r7t33
rlabel alu1 -380 -248 -380 -248 1 z2t3
rlabel polyct1 -372 -252 -372 -252 1 z2t3
rlabel alu1 -399 -280 -399 -280 6 vss
rlabel alu1 -399 -216 -399 -216 6 vdd
rlabel alu1 -391 -252 -391 -252 1 c7inv
rlabel alu1 -399 -256 -399 -256 1 c7inv
rlabel alu1 -399 -236 -399 -236 1 c7
rlabel alu1 -407 -252 -407 -252 1 c7
rlabel alu1 -479 -144 -479 -144 8 vss
rlabel alu1 -479 -208 -479 -208 8 vdd
rlabel alu1 -427 -188 -427 -188 5 c7
rlabel polyct1 -419 -180 -419 -180 5 c7
rlabel alu1 -491 -176 -491 -176 5 c4
rlabel alu1 -499 -188 -499 -188 5 c4
rlabel alu0 -437 -184 -437 -184 5 r6t4
rlabel alu0 -427 -171 -427 -171 5 r6t4
rlabel alu0 -465 -196 -465 -196 5 r6t4
rlabel alu0 -457 -172 -457 -172 5 r6t4
rlabel alu0 -458 -184 -458 -184 5 r6t44
rlabel polyct0 -471 -172 -471 -172 5 r6t44
rlabel alu0 -448 -160 -448 -160 5 r6t44
rlabel alu0 -509 -184 -509 -184 5 r6t444
rlabel alu0 -518 -196 -518 -196 5 r6t444
rlabel alu0 -494 -157 -494 -157 5 r6t444
rlabel alu1 -539 -172 -539 -172 5 z3t3
rlabel alu1 -531 -156 -531 -156 5 z3t3
rlabel alu1 -523 -156 -523 -156 5 z3t3
rlabel alu1 -531 -188 -531 -188 5 z3t3
rlabel alu1 -404 -135 -404 -135 6 vss
rlabel alu1 -404 -71 -404 -71 6 vdd
rlabel alu1 -388 -91 -388 -91 1 Y2
rlabel alu1 -396 -99 -396 -99 1 Y2
rlabel alu1 -404 -107 -404 -107 1 X3
rlabel alu1 -396 -111 -396 -111 1 X3
rlabel alu1 -420 -107 -420 -107 1 X3Y2
rlabel alu0 -399 -87 -399 -87 1 r5t4
rlabel alu0 -412 -104 -412 -104 1 r5t4
rlabel alu0 -396 -123 -396 -123 1 r5t4
rlabel alu1 -412 -123 -412 -123 1 X3Y2
rlabel alu1 -440 -136 -440 -136 6 vss
rlabel alu1 -440 -72 -440 -72 6 vdd
rlabel alu1 -432 -108 -432 -108 1 X3Y2
rlabel alu1 -440 -112 -440 -112 1 X3Y2
rlabel alu1 -440 -92 -440 -92 1 X3Y2inv
rlabel alu1 -448 -108 -448 -108 1 X3Y2inv
rlabel polyct1 -443 -172 -443 -172 1 X3Y2inv
rlabel alu1 -435 -168 -435 -168 1 X3Y2inv
rlabel alu0 -442 -227 -442 -227 1 r7t44
rlabel alu0 -470 -232 -470 -232 1 r7t44
rlabel alu0 -454 -269 -454 -269 1 r7t4
rlabel alu0 -434 -268 -434 -268 1 r7t4
rlabel polyct1 -466 -252 -466 -252 1 c4
rlabel alu1 -474 -248 -474 -248 1 c4
rlabel alu1 -426 -248 -426 -248 1 c7
rlabel alu1 -434 -236 -434 -236 1 c7
rlabel alu1 -446 -216 -446 -216 6 vdd
rlabel alu1 -446 -280 -446 -280 6 vss
rlabel alu1 -442 -252 -442 -252 1 X3Y2inv
rlabel alu1 -434 -260 -434 -260 1 X3Y2inv
rlabel alu1 -426 -260 -426 -260 1 X3Y2inv
rlabel alu1 -221 -287 -221 -287 8 vss
rlabel alu1 -221 -351 -221 -351 8 vdd
rlabel alu1 -209 -307 -209 -307 5 X0
rlabel alu1 -217 -303 -217 -303 5 X0
rlabel polyct1 -225 -315 -225 -315 5 Y3
rlabel alu1 -217 -323 -217 -323 5 Y3
rlabel alu1 -225 -331 -225 -331 5 X0Y3inv
rlabel alu1 -233 -311 -233 -311 5 X0Y3inv
rlabel alu0 -258 -398 -258 -398 1 r9t11
rlabel alu0 -218 -368 -218 -368 1 r9t11
rlabel alu0 -242 -383 -242 -383 1 r9t11
rlabel alu0 -226 -393 -226 -393 1 r9t11
rlabel alu0 -232 -405 -232 -405 1 r9t1
rlabel alu0 -224 -380 -224 -380 1 r9t1
rlabel alu0 -212 -393 -212 -393 1 r9t1
rlabel alu1 -219 -409 -219 -409 1 Z3
rlabel alu1 -211 -409 -211 -409 1 Z3
rlabel alu1 -203 -389 -203 -389 1 Z3
rlabel alu1 -211 -377 -211 -377 1 Z3
rlabel alu1 -251 -369 -251 -369 1 z3t1
rlabel alu1 -259 -377 -259 -377 1 z3t1
rlabel alu1 -251 -401 -251 -401 1 X0Y3inv
rlabel polyct1 -243 -397 -243 -397 1 X0Y3inv
rlabel alu1 -231 -357 -231 -357 6 vdd
rlabel alu1 -231 -421 -231 -421 6 vss
rlabel alu1 -243 -428 -243 -428 8 vss
rlabel alu1 -243 -492 -243 -492 8 vdd
rlabel alu1 -227 -472 -227 -472 5 X0Y3inv
rlabel alu1 -235 -464 -235 -464 5 X0Y3inv
rlabel alu1 -243 -456 -243 -456 5 z3t1
rlabel alu1 -235 -452 -235 -452 5 z3t1
rlabel alu0 -251 -459 -251 -459 5 r10t1
rlabel alu0 -238 -476 -238 -476 5 r10t1
rlabel alu1 -450 -244 -450 -244 1 c8inv
rlabel alu1 -458 -256 -458 -256 1 c8inv
rlabel alu1 -450 -260 -450 -260 1 c8inv
rlabel alu1 -492 -236 -492 -236 1 c8
rlabel alu1 -500 -252 -500 -252 1 c8
rlabel alu1 -492 -256 -492 -256 1 c8inv
rlabel alu1 -484 -252 -484 -252 1 c8inv
rlabel alu1 -492 -216 -492 -216 6 vdd
rlabel alu1 -492 -280 -492 -280 6 vss
rlabel alu1 -259 -456 -259 -456 1 c9
rlabel alu1 -251 -440 -251 -440 1 c9
rlabel alu1 -367 -288 -367 -288 8 vss
rlabel alu1 -367 -352 -367 -352 8 vdd
rlabel alu1 -363 -324 -363 -324 5 Y3
rlabel polyct1 -371 -316 -371 -316 5 Y3
rlabel alu1 -355 -308 -355 -308 5 X1
rlabel alu1 -363 -304 -363 -304 5 X1
rlabel alu1 -371 -332 -371 -332 5 X1Y3inv
rlabel alu1 -379 -312 -379 -312 5 X1Y3inv
rlabel alu1 -393 -423 -393 -423 6 vss
rlabel alu1 -393 -359 -393 -359 6 vdd
rlabel alu1 -341 -379 -341 -379 1 c9
rlabel polyct1 -333 -387 -333 -387 1 c9
rlabel polyct1 -357 -395 -357 -395 1 X1Y3inv
rlabel alu1 -349 -399 -349 -399 1 X1Y3inv
rlabel alu0 -351 -383 -351 -383 1 r9t2
rlabel alu0 -341 -396 -341 -396 1 r9t2
rlabel alu0 -379 -371 -379 -371 1 r9t2
rlabel polyct0 -385 -395 -385 -395 1 r9t22
rlabel alu0 -372 -383 -372 -383 1 r9t22
rlabel alu0 -362 -407 -362 -407 1 r9t22
rlabel alu0 -371 -395 -371 -395 1 r9t2
rlabel alu0 -432 -371 -432 -371 1 r9t222
rlabel alu0 -408 -410 -408 -410 1 r9t222
rlabel alu1 -437 -411 -437 -411 1 Z4
rlabel alu1 -445 -411 -445 -411 1 Z4
rlabel alu1 -453 -395 -453 -395 1 Z4
rlabel alu1 -413 -379 -413 -379 1 z3t2
rlabel alu1 -405 -391 -405 -391 1 z3t2
rlabel alu1 -400 -430 -400 -430 8 vss
rlabel alu1 -400 -494 -400 -494 8 vdd
rlabel alu1 -445 -430 -445 -430 8 vss
rlabel alu1 -445 -494 -445 -494 8 vdd
rlabel alu1 -380 -462 -380 -462 5 c9
rlabel alu1 -388 -474 -388 -474 5 c9
rlabel alu1 -428 -462 -428 -462 5 z3t2
rlabel polyct1 -420 -458 -420 -458 5 z3t2
rlabel alu1 -380 -450 -380 -450 5 X1Y3inv
rlabel alu1 -388 -450 -388 -450 5 X1Y3inv
rlabel alu1 -396 -458 -396 -458 5 X1Y3inv
rlabel pdifct1 -396 -474 -396 -474 5 c10inv
rlabel alu1 -404 -466 -404 -466 5 c10inv
rlabel alu1 -412 -454 -412 -454 5 c10inv
rlabel alu1 -404 -450 -404 -450 5 c10inv
rlabel alu0 -396 -483 -396 -483 5 r10t2
rlabel alu0 -424 -478 -424 -478 5 r10t2
rlabel alu0 -408 -441 -408 -441 5 r10t22
rlabel alu0 -388 -442 -388 -442 5 r10t22
rlabel alu1 -445 -454 -445 -454 5 c10inv
rlabel alu1 -437 -458 -437 -458 5 c10inv
rlabel alu1 -453 -458 -453 -458 5 c10
rlabel alu1 -445 -474 -445 -474 5 c10
rlabel alu1 -479 -308 -479 -308 5 X2
rlabel alu1 -487 -304 -487 -304 5 X2
rlabel alu1 -487 -324 -487 -324 5 Y3
rlabel polyct1 -495 -316 -495 -316 5 Y3
rlabel alu1 -491 -352 -491 -352 8 vdd
rlabel alu1 -491 -288 -491 -288 8 vss
rlabel alu1 -503 -312 -503 -312 1 X2Y3inv
rlabel alu1 -495 -332 -495 -332 1 X2Y3inv
rlabel alu1 -445 -379 -445 -379 1 Z4
rlabel alu0 -423 -383 -423 -383 1 r9t222
rlabel alu0 -564 -371 -564 -371 1 r9t333
rlabel alu0 -540 -410 -540 -410 1 r9t333
rlabel alu0 -555 -383 -555 -383 1 r9t333
rlabel alu0 -504 -383 -504 -383 1 r9t33
rlabel polyct0 -517 -395 -517 -395 1 r9t33
rlabel alu0 -494 -407 -494 -407 1 r9t33
rlabel alu0 -503 -395 -503 -395 1 r9t3
rlabel alu0 -511 -371 -511 -371 1 r9t3
rlabel alu0 -483 -383 -483 -383 1 r9t3
rlabel alu0 -473 -396 -473 -396 1 r9t3
rlabel alu1 -569 -411 -569 -411 1 Z5
rlabel alu1 -577 -411 -577 -411 1 Z5
rlabel alu1 -585 -395 -585 -395 1 Z5
rlabel alu1 -577 -379 -577 -379 1 Z5
rlabel alu1 -545 -379 -545 -379 1 z3t3
rlabel alu1 -537 -391 -537 -391 1 z3t3
rlabel alu1 -481 -399 -481 -399 1 X2Y3inv
rlabel polyct1 -489 -395 -489 -395 1 X2Y3inv
rlabel alu1 -473 -379 -473 -379 1 c10
rlabel polyct1 -465 -387 -465 -387 1 c10
rlabel alu1 -525 -359 -525 -359 6 vdd
rlabel alu1 -525 -423 -525 -423 6 vss
rlabel alu0 -517 -443 -517 -443 5 r10t33
rlabel alu0 -537 -442 -537 -442 5 r10t33
rlabel alu0 -553 -479 -553 -479 5 r10t3
rlabel alu0 -525 -484 -525 -484 5 r10t3
rlabel alu1 -585 -459 -585 -459 5 c11
rlabel alu1 -577 -475 -577 -475 5 c11
rlabel alu1 -577 -455 -577 -455 5 c11inv
rlabel alu1 -569 -459 -569 -459 5 c11inv
rlabel alu1 -533 -451 -533 -451 5 c11inv
rlabel alu1 -541 -455 -541 -455 5 c11inv
rlabel alu1 -533 -467 -533 -467 5 c11inv
rlabel pdifct1 -525 -475 -525 -475 5 c11inv
rlabel alu1 -557 -463 -557 -463 5 z3t3
rlabel polyct1 -549 -459 -549 -459 5 z3t3
rlabel alu1 -509 -451 -509 -451 5 X2Y3inv
rlabel alu1 -517 -451 -517 -451 5 X2Y3inv
rlabel alu1 -525 -459 -525 -459 5 X2Y3inv
rlabel alu1 -517 -475 -517 -475 5 c10
rlabel alu1 -509 -463 -509 -463 5 c10
rlabel alu1 -577 -495 -577 -495 8 vdd
rlabel alu1 -577 -431 -577 -431 8 vss
rlabel alu1 -529 -495 -529 -495 8 vdd
rlabel alu1 -529 -431 -529 -431 8 vss
rlabel alu1 -560 -288 -560 -288 8 vss
rlabel alu1 -560 -352 -560 -352 8 vdd
rlabel alu1 -544 -332 -544 -332 5 Y3
rlabel alu1 -552 -324 -552 -324 5 Y3
rlabel alu1 -552 -312 -552 -312 5 X3
rlabel alu1 -560 -316 -560 -316 5 X3
rlabel alu1 -576 -316 -576 -316 5 X3Y3
rlabel alu1 -568 -300 -568 -300 5 X3Y3
rlabel alu0 -555 -336 -555 -336 5 r8t1
rlabel alu0 -568 -319 -568 -319 5 r8t1
rlabel alu0 -552 -300 -552 -300 1 r8t1
rlabel alu1 -657 -423 -657 -423 6 vss
rlabel alu1 -657 -359 -657 -359 6 vdd
rlabel alu1 -605 -379 -605 -379 1 c11
rlabel polyct1 -597 -387 -597 -387 1 c11
rlabel alu1 -613 -399 -613 -399 1 X3Y3
rlabel polyct1 -621 -395 -621 -395 1 X3Y3
rlabel alu1 -677 -379 -677 -379 1 c8
rlabel alu1 -669 -391 -669 -391 1 c8
rlabel alu1 -709 -379 -709 -379 1 Z6
rlabel alu1 -717 -395 -717 -395 1 Z6
rlabel alu1 -709 -411 -709 -411 1 Z6
rlabel alu1 -701 -411 -701 -411 1 Z6
rlabel alu0 -605 -396 -605 -396 1 r9t4
rlabel alu0 -615 -383 -615 -383 1 r9t4
rlabel alu0 -643 -371 -643 -371 1 r9t4
rlabel alu0 -635 -395 -635 -395 1 r9t4
rlabel alu0 -636 -383 -636 -383 1 r9t44
rlabel polyct0 -649 -395 -649 -395 1 r9t44
rlabel alu0 -626 -407 -626 -407 1 r9t44
rlabel alu0 -687 -383 -687 -383 1 r9t444
rlabel alu0 -696 -371 -696 -371 1 r9t444
rlabel alu0 -672 -410 -672 -410 1 r9t444
rlabel alu1 -661 -431 -661 -431 8 vss
rlabel alu1 -661 -495 -661 -495 8 vdd
rlabel alu1 -709 -494 -709 -494 8 vdd
rlabel alu1 -709 -430 -709 -430 8 vss
rlabel alu1 -649 -475 -649 -475 5 c11
rlabel alu1 -641 -463 -641 -463 5 c11
rlabel alu1 -657 -459 -657 -459 5 X3Y3
rlabel alu1 -649 -451 -649 -451 5 X3Y3
rlabel via1 -641 -451 -641 -451 5 X3Y3
rlabel alu1 -689 -463 -689 -463 5 c8
rlabel polyct1 -681 -459 -681 -459 5 c8
rlabel pdifct1 -657 -475 -657 -475 5 c12inv
rlabel alu1 -665 -467 -665 -467 5 c12inv
rlabel alu1 -673 -455 -673 -455 5 c12inv
rlabel alu1 -665 -451 -665 -451 5 c12inv
rlabel alu0 -657 -484 -657 -484 5 r10t4
rlabel alu0 -685 -479 -685 -479 5 r10t4
rlabel alu0 -649 -443 -649 -443 5 r10t44
rlabel alu0 -669 -442 -669 -442 5 r10t44
rlabel alu1 -701 -458 -701 -458 5 c12inv
rlabel alu1 -709 -454 -709 -454 5 c12inv
rlabel alu1 -709 -474 -709 -474 5 c12
rlabel alu1 -717 -458 -717 -458 5 c12
rlabel alu1 -757 -430 -757 -430 2 vss
rlabel alu1 -757 -494 -757 -494 2 vdd
rlabel alu1 -737 -450 -737 -450 1 vdd
rlabel polyct1 -745 -454 -745 -454 1 vdd
rlabel alu1 -729 -474 -729 -474 1 c12
rlabel alu1 -737 -482 -737 -482 1 c12
rlabel alu0 -730 -453 -730 -453 1 r10t5
rlabel alu0 -762 -458 -762 -458 1 r10t5
rlabel alu0 -770 -483 -770 -483 1 r10t5
rlabel alu0 -776 -458 -776 -458 1 r10t55
rlabel alu0 -764 -471 -764 -471 1 r10t55
rlabel alu0 -756 -446 -756 -446 1 r10t55
rlabel alu1 -769 -442 -769 -442 1 Z7
rlabel alu1 -777 -442 -777 -442 1 Z7
rlabel alu1 -785 -462 -785 -462 1 Z7
rlabel alu1 -777 -474 -777 -474 1 Z7
<< end >>
