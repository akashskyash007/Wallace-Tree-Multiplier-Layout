magic
tech scmos
timestamp 1199202065
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 9 56 11 61
rect 21 56 23 61
rect 9 35 11 38
rect 21 35 23 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 21 33 27 35
rect 21 31 23 33
rect 25 31 27 33
rect 21 29 27 31
rect 9 22 11 29
rect 21 26 23 29
rect 9 8 11 13
rect 21 12 23 17
<< ndif >>
rect 13 22 21 26
rect 4 19 9 22
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 11 17 21 22
rect 23 24 30 26
rect 23 22 26 24
rect 28 22 30 24
rect 23 20 30 22
rect 23 17 28 20
rect 11 15 15 17
rect 17 15 19 17
rect 11 13 19 15
<< pdif >>
rect 13 67 19 69
rect 13 65 15 67
rect 17 65 19 67
rect 13 56 19 65
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 4 38 9 43
rect 11 38 21 56
rect 23 51 28 56
rect 23 49 30 51
rect 23 47 26 49
rect 28 47 30 49
rect 23 45 30 47
rect 23 38 28 45
<< alu1 >>
rect -2 67 34 72
rect -2 65 5 67
rect 7 65 15 67
rect 17 65 25 67
rect 27 65 34 67
rect -2 64 34 65
rect 2 54 14 59
rect 2 52 4 54
rect 6 53 14 54
rect 2 47 6 52
rect 2 45 4 47
rect 2 19 6 45
rect 26 35 30 43
rect 18 33 30 35
rect 18 31 23 33
rect 25 31 30 33
rect 18 29 30 31
rect 2 17 7 19
rect 2 15 4 17
rect 6 15 7 17
rect 2 13 7 15
rect -2 7 34 8
rect -2 5 22 7
rect 24 5 34 7
rect -2 0 34 5
<< ptie >>
rect 17 7 29 9
rect 17 5 22 7
rect 24 5 29 7
rect 17 3 29 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
rect 23 67 29 69
rect 23 65 25 67
rect 27 65 29 67
rect 23 63 29 65
<< nmos >>
rect 9 13 11 22
rect 21 17 23 26
<< pmos >>
rect 9 38 11 56
rect 21 38 23 56
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 23 31 25 33
<< ndifct0 >>
rect 26 22 28 24
rect 15 15 17 17
<< ndifct1 >>
rect 4 15 6 17
<< ntiect1 >>
rect 5 65 7 67
rect 25 65 27 67
<< ptiect1 >>
rect 22 5 24 7
<< pdifct0 >>
rect 26 47 28 49
<< pdifct1 >>
rect 15 65 17 67
rect 4 52 6 54
rect 4 45 6 47
<< alu0 >>
rect 6 43 7 53
rect 10 49 30 50
rect 10 47 26 49
rect 28 47 30 49
rect 10 46 30 47
rect 10 33 14 46
rect 10 31 11 33
rect 13 31 14 33
rect 10 25 14 31
rect 10 24 30 25
rect 10 22 26 24
rect 28 22 30 24
rect 10 21 30 22
rect 13 17 19 18
rect 13 15 15 17
rect 17 15 19 17
rect 13 8 19 15
<< labels >>
rlabel alu0 12 35 12 35 6 an
rlabel alu0 20 23 20 23 6 an
rlabel alu0 20 48 20 48 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 12 56 12 56 6 z
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 20 32 20 32 6 a
rlabel alu1 28 36 28 36 6 a
<< end >>
