magic
tech scmos
timestamp 1199203552
<< ab >>
rect 0 0 96 72
<< nwell >>
rect -5 32 101 77
<< pwell >>
rect -5 -5 101 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 65 31 70
rect 36 68 64 70
rect 36 65 38 68
rect 55 60 57 64
rect 62 60 64 68
rect 74 66 76 70
rect 9 35 11 38
rect 19 35 21 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 29 30 31 38
rect 36 34 38 38
rect 55 35 57 38
rect 51 33 57 35
rect 51 31 53 33
rect 55 31 57 33
rect 51 30 57 31
rect 10 20 12 29
rect 19 25 21 29
rect 29 28 57 30
rect 62 34 64 38
rect 74 35 76 38
rect 62 32 70 34
rect 62 30 66 32
rect 68 30 70 32
rect 62 28 70 30
rect 74 33 81 35
rect 74 31 77 33
rect 79 31 81 33
rect 74 29 81 31
rect 17 23 21 25
rect 37 24 39 28
rect 62 25 64 28
rect 74 25 76 29
rect 17 20 19 23
rect 27 20 29 24
rect 37 8 39 12
rect 62 8 64 12
rect 10 2 12 7
rect 17 2 19 7
rect 27 4 29 7
rect 74 4 76 12
rect 27 2 76 4
<< ndif >>
rect 32 20 37 24
rect 2 7 10 20
rect 12 7 17 20
rect 19 17 27 20
rect 19 15 22 17
rect 24 15 27 17
rect 19 7 27 15
rect 29 18 37 20
rect 29 16 32 18
rect 34 16 37 18
rect 29 12 37 16
rect 39 16 46 24
rect 39 14 42 16
rect 44 14 46 16
rect 39 12 46 14
rect 55 23 62 25
rect 55 21 57 23
rect 59 21 62 23
rect 55 16 62 21
rect 55 14 57 16
rect 59 14 62 16
rect 55 12 62 14
rect 64 16 74 25
rect 64 14 69 16
rect 71 14 74 16
rect 64 12 74 14
rect 76 18 81 25
rect 76 16 83 18
rect 76 14 79 16
rect 81 14 83 16
rect 76 12 83 14
rect 29 7 34 12
rect 2 5 4 7
rect 6 5 8 7
rect 2 3 8 5
<< pdif >>
rect 4 60 9 66
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 54 9 56
rect 4 38 9 54
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 38 19 47
rect 21 65 26 66
rect 21 49 29 65
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 38 36 65
rect 38 63 46 65
rect 38 61 41 63
rect 43 61 46 63
rect 38 50 46 61
rect 66 64 74 66
rect 66 62 69 64
rect 71 62 74 64
rect 66 60 74 62
rect 38 38 44 50
rect 50 44 55 60
rect 48 42 55 44
rect 48 40 50 42
rect 52 40 55 42
rect 48 38 55 40
rect 57 38 62 60
rect 64 38 74 60
rect 76 59 81 66
rect 76 57 83 59
rect 76 55 79 57
rect 81 55 83 57
rect 76 53 83 55
rect 76 38 81 53
<< alu1 >>
rect -2 67 98 72
rect -2 65 89 67
rect 91 65 98 67
rect -2 64 98 65
rect 2 49 18 50
rect 2 47 14 49
rect 16 47 18 49
rect 2 46 18 47
rect 2 18 6 46
rect 58 35 62 51
rect 66 45 78 51
rect 50 33 62 35
rect 50 31 53 33
rect 55 31 62 33
rect 50 29 62 31
rect 66 32 70 35
rect 68 30 70 32
rect 74 34 78 45
rect 74 33 81 34
rect 74 31 77 33
rect 79 31 81 33
rect 74 30 81 31
rect 66 26 70 30
rect 66 21 79 26
rect 2 17 26 18
rect 2 15 22 17
rect 24 15 26 17
rect 2 14 26 15
rect -2 7 98 8
rect -2 5 4 7
rect 6 5 89 7
rect 91 5 98 7
rect -2 0 98 5
<< ptie >>
rect 87 7 93 24
rect 87 5 89 7
rect 91 5 93 7
rect 87 3 93 5
<< ntie >>
rect 87 67 93 69
rect 87 65 89 67
rect 91 65 93 67
rect 87 40 93 65
<< nmos >>
rect 10 7 12 20
rect 17 7 19 20
rect 27 7 29 20
rect 37 12 39 24
rect 62 12 64 25
rect 74 12 76 25
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 65
rect 36 38 38 65
rect 55 38 57 60
rect 62 38 64 60
rect 74 38 76 66
<< polyct0 >>
rect 11 31 13 33
rect 21 31 23 33
<< polyct1 >>
rect 53 31 55 33
rect 66 30 68 32
rect 77 31 79 33
<< ndifct0 >>
rect 32 16 34 18
rect 42 14 44 16
rect 57 21 59 23
rect 57 14 59 16
rect 69 14 71 16
rect 79 14 81 16
<< ndifct1 >>
rect 22 15 24 17
rect 4 5 6 7
<< ntiect1 >>
rect 89 65 91 67
<< ptiect1 >>
rect 89 5 91 7
<< pdifct0 >>
rect 4 56 6 58
rect 24 47 26 49
rect 24 40 26 42
rect 41 61 43 63
rect 69 62 71 64
rect 50 40 52 42
rect 79 55 81 57
<< pdifct1 >>
rect 14 47 16 49
<< alu0 >>
rect 40 63 44 64
rect 40 61 41 63
rect 43 61 44 63
rect 67 62 69 64
rect 71 62 73 64
rect 67 61 73 62
rect 40 59 44 61
rect 2 58 36 59
rect 2 56 4 58
rect 6 56 36 58
rect 2 55 36 56
rect 50 57 89 58
rect 50 55 79 57
rect 81 55 89 57
rect 32 54 89 55
rect 32 51 54 54
rect 23 49 27 51
rect 23 47 24 49
rect 26 47 27 49
rect 23 42 27 47
rect 10 40 24 42
rect 26 40 27 42
rect 10 38 27 40
rect 10 33 14 38
rect 32 34 36 51
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 19 33 36 34
rect 19 31 21 33
rect 23 31 36 33
rect 19 30 36 31
rect 42 42 54 43
rect 42 40 50 42
rect 52 40 54 42
rect 42 39 54 40
rect 10 25 35 26
rect 42 25 46 39
rect 65 28 66 34
rect 10 23 61 25
rect 10 22 57 23
rect 31 21 57 22
rect 59 21 61 23
rect 31 18 35 21
rect 31 16 32 18
rect 34 16 35 18
rect 31 14 35 16
rect 40 16 46 17
rect 40 14 42 16
rect 44 14 46 16
rect 40 8 46 14
rect 55 16 61 21
rect 85 17 89 54
rect 55 14 57 16
rect 59 14 61 16
rect 55 13 61 14
rect 67 16 73 17
rect 67 14 69 16
rect 71 14 73 16
rect 67 8 73 14
rect 77 16 89 17
rect 77 14 79 16
rect 81 14 89 16
rect 77 13 89 14
<< labels >>
rlabel polyct0 12 32 12 32 6 an
rlabel alu0 33 20 33 20 6 an
rlabel alu0 27 32 27 32 6 bn
rlabel alu0 25 44 25 44 6 an
rlabel alu0 19 57 19 57 6 bn
rlabel alu0 58 19 58 19 6 an
rlabel alu0 48 41 48 41 6 an
rlabel alu0 83 15 83 15 6 bn
rlabel alu0 69 56 69 56 6 bn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 48 4 48 4 6 vss
rlabel alu1 52 32 52 32 6 a2
rlabel alu1 68 28 68 28 6 a1
rlabel alu1 60 40 60 40 6 a2
rlabel alu1 68 48 68 48 6 b
rlabel alu1 48 68 48 68 6 vdd
rlabel alu1 76 24 76 24 6 a1
rlabel alu1 76 44 76 44 6 b
<< end >>
