magic
tech scmos
timestamp 1199203187
<< ab >>
rect 0 0 136 80
<< nwell >>
rect -5 36 141 88
<< pwell >>
rect -5 -8 141 36
<< poly >>
rect 31 70 33 74
rect 39 70 41 74
rect 47 70 49 74
rect 57 70 59 74
rect 65 70 67 74
rect 73 70 75 74
rect 83 70 85 74
rect 91 70 93 74
rect 99 70 101 74
rect 109 70 111 74
rect 116 70 118 74
rect 123 70 125 74
rect 9 61 11 65
rect 19 63 21 68
rect 9 39 11 42
rect 19 39 21 42
rect 31 39 33 42
rect 39 39 41 42
rect 47 39 49 42
rect 57 39 59 42
rect 65 39 67 42
rect 73 39 75 42
rect 83 39 85 42
rect 91 39 93 42
rect 99 39 101 42
rect 109 39 111 42
rect 9 37 21 39
rect 9 35 14 37
rect 16 35 21 37
rect 9 33 21 35
rect 26 37 33 39
rect 26 35 28 37
rect 30 35 33 37
rect 26 33 33 35
rect 37 37 43 39
rect 47 37 59 39
rect 63 37 69 39
rect 37 35 39 37
rect 41 35 43 37
rect 37 33 43 35
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 63 35 65 37
rect 67 35 69 37
rect 63 33 69 35
rect 73 37 85 39
rect 89 37 95 39
rect 73 35 75 37
rect 77 35 79 37
rect 73 33 79 35
rect 89 35 91 37
rect 93 35 95 37
rect 89 33 95 35
rect 99 37 111 39
rect 99 36 105 37
rect 99 34 101 36
rect 103 34 105 36
rect 9 30 11 33
rect 19 30 21 33
rect 29 29 33 33
rect 51 30 53 33
rect 29 27 43 29
rect 29 24 31 27
rect 41 24 43 27
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 67 28 69 33
rect 89 28 91 33
rect 67 26 91 28
rect 67 23 69 26
rect 77 23 79 26
rect 89 23 91 26
rect 99 32 105 34
rect 116 33 118 42
rect 123 39 125 42
rect 123 37 134 39
rect 123 35 130 37
rect 132 35 134 37
rect 123 33 134 35
rect 99 23 101 32
rect 113 31 119 33
rect 113 29 115 31
rect 117 29 119 31
rect 113 27 119 29
rect 125 23 127 33
rect 41 6 43 10
rect 51 6 53 10
rect 67 8 69 13
rect 77 8 79 13
rect 125 12 127 17
rect 89 6 91 11
rect 99 6 101 11
<< ndif >>
rect 4 23 9 30
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 12 9 17
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 12 19 26
rect 21 24 26 30
rect 46 24 51 30
rect 21 21 29 24
rect 21 19 24 21
rect 26 19 29 21
rect 21 12 29 19
rect 31 14 41 24
rect 31 12 35 14
rect 37 12 41 14
rect 33 10 41 12
rect 43 21 51 24
rect 43 19 46 21
rect 48 19 51 21
rect 43 10 51 19
rect 53 23 65 30
rect 53 14 67 23
rect 53 12 59 14
rect 61 13 67 14
rect 69 21 77 23
rect 69 19 72 21
rect 74 19 77 21
rect 69 13 77 19
rect 79 13 89 23
rect 61 12 65 13
rect 53 10 65 12
rect 81 11 89 13
rect 91 21 99 23
rect 91 19 94 21
rect 96 19 99 21
rect 91 11 99 19
rect 101 11 109 23
rect 118 21 125 23
rect 118 19 120 21
rect 122 19 125 21
rect 118 17 125 19
rect 127 21 134 23
rect 127 19 130 21
rect 132 19 134 21
rect 127 17 134 19
rect 81 9 83 11
rect 85 9 87 11
rect 81 7 87 9
rect 103 9 105 11
rect 107 9 109 11
rect 103 7 109 9
<< pdif >>
rect 23 68 31 70
rect 23 66 25 68
rect 27 66 31 68
rect 23 63 31 66
rect 14 61 19 63
rect 2 59 9 61
rect 2 57 4 59
rect 6 57 9 59
rect 2 42 9 57
rect 11 59 19 61
rect 11 57 14 59
rect 16 57 19 59
rect 11 52 19 57
rect 11 50 14 52
rect 16 50 19 52
rect 11 42 19 50
rect 21 42 31 63
rect 33 42 39 70
rect 41 42 47 70
rect 49 61 57 70
rect 49 59 52 61
rect 54 59 57 61
rect 49 42 57 59
rect 59 42 65 70
rect 67 42 73 70
rect 75 68 83 70
rect 75 66 78 68
rect 80 66 83 68
rect 75 42 83 66
rect 85 42 91 70
rect 93 42 99 70
rect 101 61 109 70
rect 101 59 104 61
rect 106 59 109 61
rect 101 42 109 59
rect 111 42 116 70
rect 118 42 123 70
rect 125 68 134 70
rect 125 66 130 68
rect 132 66 134 68
rect 125 61 134 66
rect 125 59 130 61
rect 132 59 134 61
rect 125 42 134 59
<< alu1 >>
rect -2 81 138 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 138 81
rect -2 68 138 79
rect 16 61 108 62
rect 16 59 52 61
rect 54 59 104 61
rect 106 59 108 61
rect 16 58 108 59
rect 2 29 6 51
rect 25 50 134 54
rect 17 39 23 46
rect 10 37 23 39
rect 10 35 14 37
rect 16 35 23 37
rect 10 33 23 35
rect 41 42 69 46
rect 41 39 45 42
rect 34 37 45 39
rect 34 35 39 37
rect 41 35 45 37
rect 34 34 45 35
rect 49 37 55 38
rect 49 35 51 37
rect 53 35 55 37
rect 2 28 18 29
rect 2 26 14 28
rect 16 26 18 28
rect 2 25 18 26
rect 34 25 38 34
rect 49 30 55 35
rect 63 37 69 42
rect 63 35 65 37
rect 67 35 69 37
rect 63 34 69 35
rect 73 37 79 50
rect 73 35 75 37
rect 77 35 79 37
rect 73 34 79 35
rect 89 42 119 46
rect 89 37 95 42
rect 89 35 91 37
rect 93 35 95 37
rect 89 34 95 35
rect 102 36 106 38
rect 103 34 106 36
rect 102 30 106 34
rect 49 26 106 30
rect 113 31 119 42
rect 129 37 134 50
rect 129 35 130 37
rect 132 35 134 37
rect 129 33 134 35
rect 113 29 115 31
rect 117 29 119 31
rect 113 26 119 29
rect -2 11 138 12
rect -2 9 83 11
rect 85 9 105 11
rect 107 9 138 11
rect -2 1 138 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 138 1
rect -2 -2 138 -1
<< ptie >>
rect 0 1 136 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 136 1
rect 0 -3 136 -1
<< ntie >>
rect 0 81 136 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 136 81
rect 0 77 136 79
<< nmos >>
rect 9 12 11 30
rect 19 12 21 30
rect 29 12 31 24
rect 41 10 43 24
rect 51 10 53 30
rect 67 13 69 23
rect 77 13 79 23
rect 89 11 91 23
rect 99 11 101 23
rect 125 17 127 23
<< pmos >>
rect 9 42 11 61
rect 19 42 21 63
rect 31 42 33 70
rect 39 42 41 70
rect 47 42 49 70
rect 57 42 59 70
rect 65 42 67 70
rect 73 42 75 70
rect 83 42 85 70
rect 91 42 93 70
rect 99 42 101 70
rect 109 42 111 70
rect 116 42 118 70
rect 123 42 125 70
<< polyct0 >>
rect 28 35 30 37
rect 101 34 102 36
<< polyct1 >>
rect 14 35 16 37
rect 39 35 41 37
rect 51 35 53 37
rect 65 35 67 37
rect 75 35 77 37
rect 91 35 93 37
rect 102 34 103 36
rect 130 35 132 37
rect 115 29 117 31
<< ndifct0 >>
rect 4 19 6 21
rect 24 19 26 21
rect 35 12 37 14
rect 46 19 48 21
rect 59 12 61 14
rect 72 19 74 21
rect 94 19 96 21
rect 120 19 122 21
rect 130 19 132 21
<< ndifct1 >>
rect 14 26 16 28
rect 83 9 85 11
rect 105 9 107 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
<< pdifct0 >>
rect 25 66 27 68
rect 4 57 6 59
rect 14 57 16 59
rect 14 50 16 52
rect 78 66 80 68
rect 130 66 132 68
rect 130 59 132 61
<< pdifct1 >>
rect 52 59 54 61
rect 104 59 106 61
<< alu0 >>
rect 2 59 8 68
rect 23 66 25 68
rect 27 66 29 68
rect 23 65 29 66
rect 76 66 78 68
rect 80 66 82 68
rect 76 65 82 66
rect 128 66 130 68
rect 132 66 134 68
rect 2 57 4 59
rect 6 57 8 59
rect 2 56 8 57
rect 13 59 16 62
rect 13 57 14 59
rect 128 61 134 66
rect 128 59 130 61
rect 132 59 134 61
rect 128 58 134 59
rect 16 57 18 58
rect 13 53 18 57
rect 2 52 18 53
rect 2 51 14 52
rect 6 50 14 51
rect 16 50 18 52
rect 6 49 18 50
rect 27 37 31 50
rect 27 35 28 37
rect 30 35 31 37
rect 27 33 31 35
rect 100 36 102 38
rect 100 34 101 36
rect 100 30 102 34
rect 2 21 124 22
rect 2 19 4 21
rect 6 19 24 21
rect 26 19 46 21
rect 48 19 72 21
rect 74 19 94 21
rect 96 19 120 21
rect 122 19 124 21
rect 2 18 124 19
rect 129 21 133 23
rect 129 19 130 21
rect 132 19 133 21
rect 33 14 39 15
rect 33 12 35 14
rect 37 12 39 14
rect 57 14 63 15
rect 57 12 59 14
rect 61 12 63 14
rect 129 12 133 19
<< labels >>
rlabel alu0 63 20 63 20 6 n3
rlabel alu1 12 36 12 36 6 b
rlabel alu1 20 40 20 40 6 b
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 36 32 36 32 6 a2
rlabel alu1 44 44 44 44 6 a2
rlabel alu1 36 52 36 52 6 a1
rlabel alu1 44 52 44 52 6 a1
rlabel alu1 28 52 28 52 6 a1
rlabel alu1 28 60 28 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 68 6 68 6 6 vss
rlabel alu1 60 28 60 28 6 a3
rlabel alu1 68 28 68 28 6 a3
rlabel alu1 76 28 76 28 6 a3
rlabel alu1 52 32 52 32 6 a3
rlabel alu1 52 44 52 44 6 a2
rlabel alu1 76 44 76 44 6 a1
rlabel alu1 60 44 60 44 6 a2
rlabel alu1 60 52 60 52 6 a1
rlabel alu1 68 52 68 52 6 a1
rlabel alu1 52 52 52 52 6 a1
rlabel alu1 52 60 52 60 6 z
rlabel alu1 60 60 60 60 6 z
rlabel alu1 68 60 68 60 6 z
rlabel alu1 76 60 76 60 6 z
rlabel alu1 68 74 68 74 6 vdd
rlabel alu1 84 28 84 28 6 a3
rlabel alu1 100 28 100 28 6 a3
rlabel alu1 92 28 92 28 6 a3
rlabel alu1 100 44 100 44 6 a2
rlabel alu1 108 44 108 44 6 a2
rlabel alu1 92 40 92 40 6 a2
rlabel alu1 100 52 100 52 6 a1
rlabel alu1 108 52 108 52 6 a1
rlabel alu1 92 52 92 52 6 a1
rlabel alu1 84 52 84 52 6 a1
rlabel alu1 84 60 84 60 6 z
rlabel alu1 100 60 100 60 6 z
rlabel alu1 92 60 92 60 6 z
rlabel alu1 132 40 132 40 6 a1
rlabel alu1 116 36 116 36 6 a2
rlabel alu1 116 52 116 52 6 a1
rlabel alu1 124 52 124 52 6 a1
<< end >>
