magic
tech scmos
timestamp 1199201770
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 78 61 84 63
rect 78 59 80 61
rect 82 59 84 61
rect 78 57 84 59
rect 71 45 77 47
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 24 39
rect 9 35 20 37
rect 22 35 24 37
rect 29 35 31 44
rect 39 41 41 44
rect 49 41 51 44
rect 38 39 44 41
rect 38 37 40 39
rect 42 37 44 39
rect 38 35 44 37
rect 48 39 55 41
rect 48 37 51 39
rect 53 37 55 39
rect 48 35 55 37
rect 59 39 61 44
rect 71 43 73 45
rect 75 43 77 45
rect 71 41 77 43
rect 59 37 66 39
rect 59 35 62 37
rect 64 35 66 37
rect 9 33 24 35
rect 28 33 34 35
rect 9 30 11 33
rect 19 30 21 33
rect 28 31 30 33
rect 32 31 34 33
rect 9 15 11 19
rect 28 29 35 31
rect 33 26 35 29
rect 40 26 42 35
rect 48 31 50 35
rect 59 31 66 35
rect 47 29 50 31
rect 54 29 66 31
rect 47 26 49 29
rect 54 26 56 29
rect 64 26 66 29
rect 71 26 73 41
rect 82 37 84 57
rect 78 35 84 37
rect 78 26 80 35
rect 88 33 94 35
rect 88 31 90 33
rect 92 31 94 33
rect 85 29 94 31
rect 85 26 87 29
rect 19 9 21 13
rect 33 6 35 10
rect 40 6 42 10
rect 47 6 49 10
rect 54 6 56 10
rect 64 6 66 10
rect 71 6 73 10
rect 78 6 80 10
rect 85 6 87 10
<< ndif >>
rect 2 23 9 30
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 19 19 26
rect 14 13 19 19
rect 21 26 26 30
rect 21 14 33 26
rect 21 13 26 14
rect 23 12 26 13
rect 28 12 33 14
rect 23 10 33 12
rect 35 10 40 26
rect 42 10 47 26
rect 49 10 54 26
rect 56 21 64 26
rect 56 19 59 21
rect 61 19 64 21
rect 56 10 64 19
rect 66 10 71 26
rect 73 10 78 26
rect 80 10 85 26
rect 87 21 94 26
rect 87 19 90 21
rect 92 19 94 21
rect 87 14 94 19
rect 87 12 90 14
rect 92 12 94 14
rect 87 10 94 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 60 29 66
rect 21 58 24 60
rect 26 58 29 60
rect 21 44 29 58
rect 31 57 39 70
rect 31 55 34 57
rect 36 55 39 57
rect 31 49 39 55
rect 31 47 34 49
rect 36 47 39 49
rect 31 44 39 47
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 44 49 66
rect 51 61 59 70
rect 51 59 54 61
rect 56 59 59 61
rect 51 44 59 59
rect 61 68 69 70
rect 61 66 64 68
rect 66 66 69 68
rect 61 44 69 66
rect 21 42 27 44
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 65 61 87 62
rect 65 59 80 61
rect 82 59 87 61
rect 65 58 87 59
rect 10 47 14 55
rect 65 54 69 58
rect 2 41 14 47
rect 10 30 14 41
rect 42 50 69 54
rect 73 50 87 54
rect 42 40 46 50
rect 73 46 77 50
rect 38 39 46 40
rect 38 37 40 39
rect 42 37 46 39
rect 38 36 46 37
rect 50 45 77 46
rect 50 43 73 45
rect 75 43 77 45
rect 50 42 77 43
rect 81 42 87 46
rect 50 39 54 42
rect 50 37 51 39
rect 53 37 54 39
rect 81 38 86 42
rect 50 35 54 37
rect 60 37 86 38
rect 60 35 62 37
rect 64 35 86 37
rect 10 28 17 30
rect 10 26 14 28
rect 16 26 17 28
rect 10 24 17 26
rect 29 33 33 35
rect 60 34 86 35
rect 29 31 30 33
rect 32 31 33 33
rect 29 30 33 31
rect 90 33 94 35
rect 92 31 94 33
rect 90 30 94 31
rect 29 26 94 30
rect 74 25 94 26
rect 74 17 78 25
rect -2 1 98 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 9 19 11 30
rect 19 13 21 30
rect 33 10 35 26
rect 40 10 42 26
rect 47 10 49 26
rect 54 10 56 26
rect 64 10 66 26
rect 71 10 73 26
rect 78 10 80 26
rect 85 10 87 26
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 44 31 70
rect 39 44 41 70
rect 49 44 51 70
rect 59 44 61 70
<< polyct0 >>
rect 20 35 22 37
<< polyct1 >>
rect 80 59 82 61
rect 40 37 42 39
rect 51 37 53 39
rect 73 43 75 45
rect 62 35 64 37
rect 30 31 32 33
rect 90 31 92 33
<< ndifct0 >>
rect 4 21 6 23
rect 26 12 28 14
rect 59 19 61 21
rect 90 19 92 21
rect 90 12 92 14
<< ndifct1 >>
rect 14 26 16 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 59 16 61
rect 14 52 16 54
rect 24 66 26 68
rect 24 58 26 60
rect 34 55 36 57
rect 34 47 36 49
rect 44 66 46 68
rect 54 59 56 61
rect 64 66 66 68
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 23 66 24 68
rect 26 66 27 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 55 17 59
rect 23 60 27 66
rect 42 66 44 68
rect 46 66 48 68
rect 42 65 48 66
rect 62 66 64 68
rect 66 66 68 68
rect 62 65 68 66
rect 23 58 24 60
rect 26 58 27 60
rect 23 56 27 58
rect 33 61 58 62
rect 33 59 54 61
rect 56 59 58 61
rect 33 58 58 59
rect 33 57 37 58
rect 14 54 17 55
rect 16 52 17 54
rect 14 50 17 52
rect 33 55 34 57
rect 36 55 37 57
rect 33 49 37 55
rect 21 47 34 49
rect 36 47 37 49
rect 21 45 37 47
rect 21 38 25 45
rect 18 37 25 38
rect 18 35 20 37
rect 22 35 25 37
rect 18 34 25 35
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 12 7 21
rect 21 22 25 34
rect 89 30 90 35
rect 21 21 63 22
rect 21 19 59 21
rect 61 19 63 21
rect 21 18 63 19
rect 88 21 94 22
rect 88 19 90 21
rect 92 19 94 21
rect 24 14 30 15
rect 24 12 26 14
rect 28 12 30 14
rect 88 14 94 19
rect 88 12 90 14
rect 92 12 94 14
<< labels >>
rlabel alu0 23 33 23 33 6 zn
rlabel alu0 35 53 35 53 6 zn
rlabel alu0 42 20 42 20 6 zn
rlabel alu0 45 60 45 60 6 zn
rlabel alu1 12 40 12 40 6 z
rlabel alu1 4 44 4 44 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 36 28 36 28 6 a
rlabel alu1 52 28 52 28 6 a
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 44 44 44 6 b
rlabel alu1 52 52 52 52 6 b
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 60 28 60 28 6 a
rlabel alu1 76 24 76 24 6 a
rlabel alu1 68 28 68 28 6 a
rlabel alu1 60 44 60 44 6 c
rlabel alu1 76 36 76 36 6 d
rlabel alu1 68 44 68 44 6 c
rlabel alu1 68 36 68 36 6 d
rlabel alu1 76 52 76 52 6 c
rlabel alu1 60 52 60 52 6 b
rlabel alu1 76 60 76 60 6 b
rlabel alu1 68 60 68 60 6 b
rlabel alu1 92 28 92 28 6 a
rlabel alu1 84 28 84 28 6 a
rlabel alu1 84 44 84 44 6 d
rlabel alu1 84 52 84 52 6 c
rlabel alu1 84 60 84 60 6 b
<< end >>
