magic
tech scmos
timestamp 1199203081
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 19 62 21 67
rect 26 62 28 67
rect 9 54 11 59
rect 40 58 42 63
rect 9 34 11 46
rect 9 32 15 34
rect 9 30 11 32
rect 13 30 15 32
rect 9 28 15 30
rect 19 28 21 46
rect 26 43 28 46
rect 40 43 42 46
rect 26 41 33 43
rect 40 41 55 43
rect 26 39 28 41
rect 30 39 33 41
rect 26 37 33 39
rect 49 39 51 41
rect 53 39 55 41
rect 49 37 55 39
rect 9 19 11 28
rect 19 26 25 28
rect 19 24 21 26
rect 23 24 25 26
rect 19 22 25 24
rect 19 19 21 22
rect 31 19 33 37
rect 51 26 53 37
rect 51 15 53 20
rect 9 7 11 12
rect 19 7 21 12
rect 31 7 33 12
<< ndif >>
rect 44 24 51 26
rect 44 22 46 24
rect 48 22 51 24
rect 44 20 51 22
rect 53 24 60 26
rect 53 22 56 24
rect 58 22 60 24
rect 53 20 60 22
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 12 9 15
rect 11 16 19 19
rect 11 14 14 16
rect 16 14 19 16
rect 11 12 19 14
rect 21 12 31 19
rect 33 16 40 19
rect 33 14 36 16
rect 38 14 40 16
rect 33 12 40 14
rect 23 7 29 12
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< pdif >>
rect 14 54 19 62
rect 2 52 9 54
rect 2 50 4 52
rect 6 50 9 52
rect 2 46 9 50
rect 11 50 19 54
rect 11 48 14 50
rect 16 48 19 50
rect 11 46 19 48
rect 21 46 26 62
rect 28 58 38 62
rect 28 56 40 58
rect 28 54 35 56
rect 37 54 40 56
rect 28 46 40 54
rect 42 52 47 58
rect 42 50 49 52
rect 42 48 45 50
rect 47 48 49 50
rect 42 46 49 48
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 57 67
rect 59 65 66 67
rect -2 64 66 65
rect 10 50 22 51
rect 10 48 14 50
rect 16 48 22 50
rect 10 45 22 48
rect 10 43 14 45
rect 2 39 14 43
rect 26 42 30 51
rect 26 41 39 42
rect 26 39 28 41
rect 30 39 39 41
rect 2 17 6 39
rect 26 38 39 39
rect 10 32 23 34
rect 10 30 11 32
rect 13 30 23 32
rect 10 21 14 30
rect 50 41 62 43
rect 50 39 51 41
rect 53 39 62 41
rect 50 37 62 39
rect 58 29 62 37
rect 2 15 4 17
rect 2 13 6 15
rect -2 7 66 8
rect -2 5 25 7
rect 27 5 49 7
rect 51 5 57 7
rect 59 5 66 7
rect -2 0 66 5
<< ptie >>
rect 47 7 61 9
rect 47 5 49 7
rect 51 5 57 7
rect 59 5 61 7
rect 47 3 61 5
<< ntie >>
rect 3 67 9 69
rect 55 67 61 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
rect 55 65 57 67
rect 59 65 61 67
rect 55 46 61 65
<< nmos >>
rect 51 20 53 26
rect 9 12 11 19
rect 19 12 21 19
rect 31 12 33 19
<< pmos >>
rect 9 46 11 54
rect 19 46 21 62
rect 26 46 28 62
rect 40 46 42 58
<< polyct0 >>
rect 21 24 23 26
<< polyct1 >>
rect 11 30 13 32
rect 28 39 30 41
rect 51 39 53 41
<< ndifct0 >>
rect 46 22 48 24
rect 56 22 58 24
rect 14 14 16 16
rect 36 14 38 16
<< ndifct1 >>
rect 4 15 6 17
rect 25 5 27 7
<< ntiect1 >>
rect 5 65 7 67
rect 57 65 59 67
<< ptiect1 >>
rect 49 5 51 7
rect 57 5 59 7
<< pdifct0 >>
rect 4 50 6 52
rect 35 54 37 56
rect 45 48 47 50
<< pdifct1 >>
rect 14 48 16 50
<< alu0 >>
rect 3 52 7 64
rect 34 56 38 64
rect 34 54 35 56
rect 37 54 38 56
rect 34 52 38 54
rect 3 50 4 52
rect 6 50 7 52
rect 3 48 7 50
rect 42 50 49 51
rect 42 48 45 50
rect 47 48 49 50
rect 42 47 49 48
rect 42 27 46 47
rect 19 26 46 27
rect 19 24 21 26
rect 23 25 46 26
rect 23 24 50 25
rect 19 23 46 24
rect 42 22 46 23
rect 48 22 50 24
rect 42 21 50 22
rect 54 24 60 25
rect 54 22 56 24
rect 58 22 60 24
rect 6 13 7 19
rect 12 16 40 17
rect 12 14 14 16
rect 16 14 36 16
rect 38 14 40 16
rect 12 13 40 14
rect 54 8 60 22
<< labels >>
rlabel alu0 26 15 26 15 6 n1
rlabel alu0 32 25 32 25 6 a2n
rlabel alu0 45 49 45 49 6 a2n
rlabel alu0 44 36 44 36 6 a2n
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 24 12 24 6 b
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 32 20 32 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 a1
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 40 36 40 6 a1
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 60 36 60 36 6 a2
rlabel polyct1 52 40 52 40 6 a2
<< end >>
