magic
tech scmos
timestamp 1199201720
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 70 11 74
rect 19 67 21 72
rect 29 67 31 72
rect 41 67 43 72
rect 9 39 11 42
rect 19 39 21 50
rect 29 47 31 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 29 11 33
rect 22 29 24 33
rect 29 29 31 41
rect 41 39 43 50
rect 41 37 47 39
rect 41 35 43 37
rect 45 35 47 37
rect 36 33 47 35
rect 36 29 38 33
rect 9 10 11 15
rect 22 7 24 12
rect 29 7 31 12
rect 36 7 38 12
<< ndif >>
rect 4 23 9 29
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 15 9 17
rect 11 15 22 29
rect 13 12 22 15
rect 24 12 29 29
rect 31 12 36 29
rect 38 22 43 29
rect 38 20 45 22
rect 38 18 41 20
rect 43 18 45 20
rect 38 16 45 18
rect 38 12 43 16
rect 13 11 20 12
rect 13 9 16 11
rect 18 9 20 11
rect 13 7 20 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 67 17 70
rect 33 71 39 73
rect 33 69 35 71
rect 37 69 39 71
rect 33 67 39 69
rect 11 65 19 67
rect 11 63 14 65
rect 16 63 19 65
rect 11 50 19 63
rect 21 61 29 67
rect 21 59 24 61
rect 26 59 29 61
rect 21 54 29 59
rect 21 52 24 54
rect 26 52 29 54
rect 21 50 29 52
rect 31 50 41 67
rect 43 64 48 67
rect 43 62 50 64
rect 43 60 46 62
rect 48 60 50 62
rect 43 58 50 60
rect 43 50 48 58
rect 11 42 17 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 35 71
rect 37 69 58 71
rect -2 68 58 69
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 2 22 6 42
rect 18 38 22 47
rect 42 46 46 55
rect 29 45 46 46
rect 29 43 31 45
rect 33 43 46 45
rect 29 42 46 43
rect 18 37 31 38
rect 18 35 21 37
rect 23 35 31 37
rect 18 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 30 47 35
rect 33 26 47 30
rect 2 21 15 22
rect 2 19 4 21
rect 6 19 15 21
rect 2 17 15 19
rect -2 11 58 12
rect -2 9 16 11
rect 18 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 15 11 29
rect 22 12 24 29
rect 29 12 31 29
rect 36 12 38 29
<< pmos >>
rect 9 42 11 70
rect 19 50 21 67
rect 29 50 31 67
rect 41 50 43 67
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 21 35 23 37
rect 43 35 45 37
<< ndifct0 >>
rect 41 18 43 20
<< ndifct1 >>
rect 4 19 6 21
rect 16 9 18 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 14 63 16 65
rect 24 59 26 61
rect 24 52 26 54
rect 46 60 48 62
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 35 69 37 71
<< alu0 >>
rect 13 65 17 68
rect 13 63 14 65
rect 16 63 17 65
rect 13 61 17 63
rect 23 62 50 63
rect 23 61 46 62
rect 23 59 24 61
rect 26 60 46 61
rect 48 60 50 62
rect 26 59 50 60
rect 23 55 28 59
rect 10 54 28 55
rect 10 52 24 54
rect 26 52 28 54
rect 10 51 28 52
rect 10 37 14 51
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 10 26 26 30
rect 22 21 26 26
rect 22 20 45 21
rect 22 18 41 20
rect 43 18 45 20
rect 22 17 45 18
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 19 53 19 53 6 zn
rlabel alu0 25 57 25 57 6 zn
rlabel alu0 33 19 33 19 6 zn
rlabel alu0 36 61 36 61 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 44 20 44 6 a
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 36 28 36 6 a
rlabel alu1 36 28 36 28 6 c
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 c
rlabel alu1 44 52 44 52 6 b
<< end >>
