magic
tech scmos
timestamp 1199203165
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 11 63 13 68
rect 18 63 20 68
rect 28 63 30 68
rect 35 63 37 68
rect 47 62 49 67
rect 57 62 59 67
rect 11 44 13 47
rect 3 42 13 44
rect 3 40 5 42
rect 7 40 9 42
rect 3 38 9 40
rect 18 37 20 47
rect 28 43 30 47
rect 35 44 37 47
rect 47 44 49 49
rect 57 46 59 49
rect 57 44 64 46
rect 13 35 20 37
rect 25 41 31 43
rect 25 39 27 41
rect 29 39 31 41
rect 25 37 31 39
rect 35 42 53 44
rect 13 34 15 35
rect 9 32 15 34
rect 9 30 11 32
rect 13 30 15 32
rect 25 31 27 37
rect 35 31 37 42
rect 47 40 49 42
rect 51 40 53 42
rect 57 42 60 44
rect 62 42 64 44
rect 57 40 64 42
rect 47 38 53 40
rect 51 35 53 38
rect 9 28 15 30
rect 13 25 15 28
rect 23 28 27 31
rect 33 28 37 31
rect 41 32 47 34
rect 51 33 56 35
rect 41 30 43 32
rect 45 30 47 32
rect 41 28 47 30
rect 23 25 25 28
rect 33 25 35 28
rect 43 25 45 28
rect 54 25 56 33
rect 61 25 63 40
rect 13 13 15 18
rect 23 13 25 18
rect 33 13 35 18
rect 43 13 45 18
rect 54 9 56 14
rect 61 9 63 14
<< ndif >>
rect 4 18 13 25
rect 15 22 23 25
rect 15 20 18 22
rect 20 20 23 22
rect 15 18 23 20
rect 25 23 33 25
rect 25 21 28 23
rect 30 21 33 23
rect 25 18 33 21
rect 35 22 43 25
rect 35 20 38 22
rect 40 20 43 22
rect 35 18 43 20
rect 45 18 54 25
rect 4 7 11 18
rect 47 16 49 18
rect 51 16 54 18
rect 47 14 54 16
rect 56 14 61 25
rect 63 23 70 25
rect 63 21 66 23
rect 68 21 70 23
rect 63 19 70 21
rect 63 14 68 19
rect 4 5 7 7
rect 9 5 11 7
rect 4 3 11 5
<< pdif >>
rect 39 67 45 69
rect 61 67 68 69
rect 39 65 41 67
rect 43 65 45 67
rect 39 63 45 65
rect 2 61 11 63
rect 2 59 4 61
rect 6 59 11 61
rect 2 54 11 59
rect 2 52 4 54
rect 6 52 11 54
rect 2 47 11 52
rect 13 47 18 63
rect 20 51 28 63
rect 20 49 23 51
rect 25 49 28 51
rect 20 47 28 49
rect 30 47 35 63
rect 37 62 45 63
rect 61 65 63 67
rect 65 65 68 67
rect 61 62 68 65
rect 37 49 47 62
rect 49 58 57 62
rect 49 56 52 58
rect 54 56 57 58
rect 49 49 57 56
rect 59 49 68 62
rect 37 47 45 49
<< alu1 >>
rect -2 67 74 72
rect -2 65 41 67
rect 43 65 63 67
rect 65 65 74 67
rect -2 64 74 65
rect 18 51 27 52
rect 18 49 23 51
rect 25 49 27 51
rect 18 48 27 49
rect 10 32 14 35
rect 10 30 11 32
rect 13 30 14 32
rect 10 27 14 30
rect 18 33 22 48
rect 33 46 63 50
rect 33 43 38 46
rect 59 44 63 46
rect 26 41 38 43
rect 26 39 27 41
rect 29 39 38 41
rect 26 37 38 39
rect 59 42 60 44
rect 62 42 63 44
rect 51 40 55 42
rect 59 40 63 42
rect 49 38 55 40
rect 51 34 55 38
rect 18 29 32 33
rect 51 30 63 34
rect 2 21 14 27
rect 2 13 6 21
rect 26 23 32 29
rect 26 21 28 23
rect 30 21 32 23
rect 26 20 32 21
rect -2 7 74 8
rect -2 5 7 7
rect 9 5 27 7
rect 29 5 35 7
rect 37 5 74 7
rect -2 0 74 5
<< ptie >>
rect 25 7 39 9
rect 25 5 27 7
rect 29 5 35 7
rect 37 5 39 7
rect 25 3 39 5
<< nmos >>
rect 13 18 15 25
rect 23 18 25 25
rect 33 18 35 25
rect 43 18 45 25
rect 54 14 56 25
rect 61 14 63 25
<< pmos >>
rect 11 47 13 63
rect 18 47 20 63
rect 28 47 30 63
rect 35 47 37 63
rect 47 49 49 62
rect 57 49 59 62
<< polyct0 >>
rect 5 40 7 42
rect 43 30 45 32
<< polyct1 >>
rect 27 39 29 41
rect 11 30 13 32
rect 49 40 51 42
rect 60 42 62 44
<< ndifct0 >>
rect 18 20 20 22
rect 38 20 40 22
rect 49 16 51 18
rect 66 21 68 23
<< ndifct1 >>
rect 28 21 30 23
rect 7 5 9 7
<< ptiect1 >>
rect 27 5 29 7
rect 35 5 37 7
<< pdifct0 >>
rect 4 59 6 61
rect 4 52 6 54
rect 52 56 54 58
<< pdifct1 >>
rect 41 65 43 67
rect 23 49 25 51
rect 63 65 65 67
<< alu0 >>
rect 3 61 7 64
rect 3 59 4 61
rect 6 59 7 61
rect 3 54 7 59
rect 3 52 4 54
rect 6 52 7 54
rect 3 50 7 52
rect 10 58 70 59
rect 10 56 52 58
rect 54 56 70 58
rect 10 55 70 56
rect 10 43 14 55
rect 3 42 14 43
rect 3 40 5 42
rect 7 40 14 42
rect 3 39 14 40
rect 47 42 53 43
rect 47 38 49 42
rect 47 37 51 38
rect 41 32 48 33
rect 41 30 43 32
rect 45 30 48 32
rect 41 29 48 30
rect 17 22 21 24
rect 17 20 18 22
rect 20 20 21 22
rect 44 26 48 29
rect 66 26 70 55
rect 37 22 41 24
rect 44 23 70 26
rect 44 22 66 23
rect 37 20 38 22
rect 40 20 41 22
rect 64 21 66 22
rect 68 21 70 23
rect 64 20 70 21
rect 17 17 21 20
rect 37 17 41 20
rect 17 13 41 17
rect 47 18 53 19
rect 47 16 49 18
rect 51 16 53 18
rect 47 8 53 16
<< labels >>
rlabel alu0 8 41 8 41 6 b
rlabel alu0 19 18 19 18 6 n4
rlabel alu0 39 18 39 18 6 n4
rlabel alu0 40 57 40 57 6 b
rlabel alu0 68 39 68 39 6 b
rlabel alu1 4 20 4 20 6 a3
rlabel alu1 12 28 12 28 6 a3
rlabel alu1 28 24 28 24 6 z
rlabel polyct1 28 40 28 40 6 b2
rlabel alu1 20 40 20 40 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 52 40 52 40 6 b1
rlabel alu1 36 44 36 44 6 b2
rlabel alu1 52 48 52 48 6 b2
rlabel alu1 44 48 44 48 6 b2
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 32 60 32 6 b1
rlabel alu1 60 48 60 48 6 b2
<< end >>
