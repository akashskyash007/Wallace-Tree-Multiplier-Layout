magic
tech scmos
timestamp 1199203511
<< ab >>
rect 0 0 128 80
<< nwell >>
rect -5 36 133 88
<< pwell >>
rect -5 -8 133 36
<< poly >>
rect 37 69 39 74
rect 47 69 49 74
rect 54 69 56 74
rect 9 61 11 65
rect 19 61 21 65
rect 85 65 87 70
rect 97 65 99 70
rect 107 65 109 70
rect 117 65 119 70
rect 9 39 11 42
rect 19 39 21 42
rect 37 39 39 50
rect 47 39 49 50
rect 54 47 56 50
rect 72 48 78 50
rect 53 45 59 47
rect 53 43 55 45
rect 57 43 59 45
rect 72 46 74 48
rect 76 46 78 48
rect 85 46 87 49
rect 72 44 87 46
rect 53 41 59 43
rect 9 37 15 39
rect 19 37 39 39
rect 43 37 49 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 25 35 27 37
rect 29 35 35 37
rect 25 33 35 35
rect 43 35 45 37
rect 47 35 49 37
rect 43 33 49 35
rect 13 25 15 33
rect 33 30 35 33
rect 45 30 47 33
rect 57 30 59 41
rect 97 40 99 49
rect 63 38 99 40
rect 107 39 109 49
rect 117 40 119 49
rect 63 36 65 38
rect 67 36 69 38
rect 63 34 69 36
rect 73 32 79 34
rect 73 30 75 32
rect 77 30 79 32
rect 73 28 79 30
rect 77 25 79 28
rect 33 16 35 21
rect 45 16 47 21
rect 57 16 59 21
rect 89 23 91 38
rect 103 37 109 39
rect 103 35 105 37
rect 107 35 109 37
rect 103 33 109 35
rect 113 38 119 40
rect 113 36 115 38
rect 117 36 119 38
rect 113 34 119 36
rect 107 29 109 33
rect 99 23 101 28
rect 107 26 111 29
rect 109 23 111 26
rect 116 23 118 34
rect 13 11 15 16
rect 77 8 79 18
rect 89 12 91 16
rect 99 8 101 16
rect 109 11 111 16
rect 116 11 118 16
rect 77 6 101 8
<< ndif >>
rect 17 25 33 30
rect 8 22 13 25
rect 6 20 13 22
rect 6 18 8 20
rect 10 18 13 20
rect 6 16 13 18
rect 15 21 33 25
rect 35 28 45 30
rect 35 26 38 28
rect 40 26 45 28
rect 35 21 45 26
rect 47 28 57 30
rect 47 26 52 28
rect 54 26 57 28
rect 47 21 57 26
rect 59 27 64 30
rect 59 25 66 27
rect 59 23 62 25
rect 64 23 66 25
rect 59 21 66 23
rect 70 23 77 25
rect 70 21 72 23
rect 74 21 77 23
rect 15 16 31 21
rect 70 18 77 21
rect 79 23 87 25
rect 79 18 89 23
rect 17 11 31 16
rect 17 9 19 11
rect 21 9 27 11
rect 29 9 31 11
rect 17 7 31 9
rect 81 16 89 18
rect 91 21 99 23
rect 91 19 94 21
rect 96 19 99 21
rect 91 16 99 19
rect 101 21 109 23
rect 101 19 104 21
rect 106 19 109 21
rect 101 16 109 19
rect 111 16 116 23
rect 118 16 126 23
rect 81 15 87 16
rect 81 13 83 15
rect 85 13 87 15
rect 81 11 87 13
rect 120 11 126 16
rect 120 9 122 11
rect 124 9 126 11
rect 120 7 126 9
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 89 71 95 73
rect 13 67 19 69
rect 13 61 17 67
rect 32 64 37 69
rect 30 62 37 64
rect 2 59 9 61
rect 2 57 4 59
rect 6 57 9 59
rect 2 52 9 57
rect 2 50 4 52
rect 6 50 9 52
rect 2 48 9 50
rect 4 42 9 48
rect 11 42 19 61
rect 21 54 26 61
rect 30 60 32 62
rect 34 60 37 62
rect 30 58 37 60
rect 21 52 28 54
rect 21 50 24 52
rect 26 50 28 52
rect 32 50 37 58
rect 39 61 47 69
rect 39 59 42 61
rect 44 59 47 61
rect 39 50 47 59
rect 49 50 54 69
rect 56 67 64 69
rect 56 65 59 67
rect 61 65 64 67
rect 89 69 91 71
rect 93 69 95 71
rect 89 65 95 69
rect 56 60 64 65
rect 56 58 59 60
rect 61 58 64 60
rect 78 62 85 65
rect 78 60 80 62
rect 82 60 85 62
rect 78 58 85 60
rect 56 50 64 58
rect 21 48 28 50
rect 21 42 26 48
rect 80 49 85 58
rect 87 49 97 65
rect 99 53 107 65
rect 99 51 102 53
rect 104 51 107 53
rect 99 49 107 51
rect 109 54 117 65
rect 109 52 112 54
rect 114 52 117 54
rect 109 49 117 52
rect 119 62 126 65
rect 119 60 122 62
rect 124 60 126 62
rect 119 58 126 60
rect 119 49 124 58
<< alu1 >>
rect -2 81 130 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 130 81
rect -2 71 130 79
rect -2 69 15 71
rect 17 69 91 71
rect 93 69 130 71
rect -2 68 130 69
rect 74 50 87 54
rect 10 42 23 46
rect 10 37 14 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 25 14 35
rect 25 37 31 38
rect 25 35 27 37
rect 29 35 31 37
rect 25 31 31 35
rect 18 25 31 31
rect 74 48 78 50
rect 76 46 78 48
rect 74 32 78 46
rect 110 54 126 55
rect 110 52 112 54
rect 114 52 126 54
rect 110 50 126 52
rect 74 30 75 32
rect 77 30 78 32
rect 74 28 78 30
rect 122 22 126 50
rect 102 21 126 22
rect 102 19 104 21
rect 106 19 126 21
rect 102 18 126 19
rect -2 11 130 12
rect -2 9 19 11
rect 21 9 27 11
rect 29 9 122 11
rect 124 9 130 11
rect -2 1 130 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 130 1
rect -2 -2 130 -1
<< ptie >>
rect 0 1 128 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 128 1
rect 0 -3 128 -1
<< ntie >>
rect 0 81 128 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 128 81
rect 0 77 128 79
<< nmos >>
rect 13 16 15 25
rect 33 21 35 30
rect 45 21 47 30
rect 57 21 59 30
rect 77 18 79 25
rect 89 16 91 23
rect 99 16 101 23
rect 109 16 111 23
rect 116 16 118 23
<< pmos >>
rect 9 42 11 61
rect 19 42 21 61
rect 37 50 39 69
rect 47 50 49 69
rect 54 50 56 69
rect 85 49 87 65
rect 97 49 99 65
rect 107 49 109 65
rect 117 49 119 65
<< polyct0 >>
rect 55 43 57 45
rect 45 35 47 37
rect 65 36 67 38
rect 105 35 107 37
rect 115 36 117 38
<< polyct1 >>
rect 74 46 76 48
rect 11 35 13 37
rect 27 35 29 37
rect 75 30 77 32
<< ndifct0 >>
rect 8 18 10 20
rect 38 26 40 28
rect 52 26 54 28
rect 62 23 64 25
rect 72 21 74 23
rect 94 19 96 21
rect 83 13 85 15
<< ndifct1 >>
rect 19 9 21 11
rect 27 9 29 11
rect 104 19 106 21
rect 122 9 124 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
<< pdifct0 >>
rect 4 57 6 59
rect 4 50 6 52
rect 32 60 34 62
rect 24 50 26 52
rect 42 59 44 61
rect 59 65 61 67
rect 59 58 61 60
rect 80 60 82 62
rect 102 51 104 53
rect 122 60 124 62
<< pdifct1 >>
rect 15 69 17 71
rect 91 69 93 71
rect 112 52 114 54
<< alu0 >>
rect 57 67 63 68
rect 57 65 59 67
rect 61 65 63 67
rect 2 62 36 63
rect 2 60 32 62
rect 34 60 36 62
rect 2 59 36 60
rect 40 61 51 62
rect 40 59 42 61
rect 44 59 51 61
rect 2 57 4 59
rect 6 57 7 59
rect 40 58 51 59
rect 2 52 7 57
rect 47 54 51 58
rect 57 60 63 65
rect 57 58 59 60
rect 61 58 63 60
rect 78 62 126 63
rect 78 60 80 62
rect 82 60 122 62
rect 124 60 126 62
rect 78 59 126 60
rect 57 57 63 58
rect 2 50 4 52
rect 6 50 7 52
rect 2 48 7 50
rect 22 52 41 53
rect 22 50 24 52
rect 26 50 41 52
rect 47 50 68 54
rect 22 49 41 50
rect 2 21 6 48
rect 37 46 41 49
rect 37 45 59 46
rect 37 43 55 45
rect 57 43 59 45
rect 37 42 59 43
rect 37 28 41 42
rect 37 26 38 28
rect 40 26 41 28
rect 37 24 41 26
rect 44 37 48 39
rect 44 35 45 37
rect 47 35 48 37
rect 64 38 68 50
rect 73 44 74 50
rect 64 36 65 38
rect 67 36 68 38
rect 44 21 48 35
rect 51 32 68 36
rect 92 38 96 59
rect 101 53 105 55
rect 101 51 102 53
rect 104 51 105 53
rect 101 46 105 51
rect 101 42 118 46
rect 114 38 118 42
rect 51 28 55 32
rect 84 37 109 38
rect 84 35 105 37
rect 107 35 109 37
rect 84 34 109 35
rect 114 36 115 38
rect 117 36 118 38
rect 51 26 52 28
rect 54 26 55 28
rect 51 24 55 26
rect 61 25 65 27
rect 61 23 62 25
rect 64 23 65 25
rect 84 24 88 34
rect 114 30 118 36
rect 61 21 65 23
rect 2 20 65 21
rect 70 23 88 24
rect 70 21 72 23
rect 74 21 88 23
rect 70 20 88 21
rect 93 26 118 30
rect 93 21 97 26
rect 2 18 8 20
rect 10 18 65 20
rect 2 17 65 18
rect 93 19 94 21
rect 96 19 97 21
rect 93 17 97 19
rect 81 15 87 16
rect 81 13 83 15
rect 85 13 87 15
rect 81 12 87 13
<< labels >>
rlabel alu0 4 40 4 40 6 an
rlabel alu0 46 28 46 28 6 an
rlabel alu0 31 51 31 51 6 bn
rlabel alu0 39 38 39 38 6 bn
rlabel alu0 19 61 19 61 6 an
rlabel alu0 33 19 33 19 6 an
rlabel alu0 63 22 63 22 6 an
rlabel alu0 53 30 53 30 6 iz
rlabel alu0 48 44 48 44 6 bn
rlabel alu0 66 43 66 43 6 iz
rlabel alu0 45 60 45 60 6 iz
rlabel alu0 79 22 79 22 6 cn
rlabel alu0 95 23 95 23 6 zn
rlabel alu0 116 36 116 36 6 zn
rlabel alu0 96 36 96 36 6 cn
rlabel alu0 103 48 103 48 6 zn
rlabel alu0 102 61 102 61 6 cn
rlabel alu1 28 32 28 32 6 b
rlabel alu1 20 28 20 28 6 b
rlabel alu1 12 32 12 32 6 a
rlabel alu1 20 44 20 44 6 a
rlabel alu1 64 6 64 6 6 vss
rlabel alu1 76 40 76 40 6 c
rlabel alu1 84 52 84 52 6 c
rlabel alu1 64 74 64 74 6 vdd
rlabel alu1 116 20 116 20 6 z
rlabel alu1 108 20 108 20 6 z
rlabel alu1 124 40 124 40 6 z
rlabel alu1 116 52 116 52 6 z
<< end >>
