magic
tech scmos
timestamp 1199203279
<< ab >>
rect 0 0 104 80
<< nwell >>
rect -5 36 109 88
<< pwell >>
rect -5 -8 109 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 31 70 33 74
rect 38 70 40 74
rect 45 70 47 74
rect 55 70 57 74
rect 62 70 64 74
rect 69 70 71 74
rect 79 58 81 63
rect 86 58 88 63
rect 93 58 95 63
rect 9 39 11 42
rect 19 39 21 42
rect 31 39 33 42
rect 9 37 21 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 28 37 34 39
rect 28 35 30 37
rect 32 35 34 37
rect 28 33 34 35
rect 38 33 40 42
rect 45 39 47 42
rect 55 39 57 42
rect 45 37 57 39
rect 9 30 11 33
rect 19 30 21 33
rect 29 24 31 33
rect 38 31 47 33
rect 38 29 43 31
rect 45 29 47 31
rect 38 27 47 29
rect 39 24 41 27
rect 51 24 53 37
rect 62 31 64 42
rect 69 39 71 42
rect 79 39 81 42
rect 69 37 81 39
rect 73 35 75 37
rect 77 35 79 37
rect 73 33 79 35
rect 62 29 68 31
rect 86 29 88 42
rect 62 27 64 29
rect 66 27 88 29
rect 93 39 95 42
rect 93 37 99 39
rect 93 35 95 37
rect 97 35 99 37
rect 93 33 99 35
rect 62 25 68 27
rect 9 11 11 16
rect 19 11 21 16
rect 93 23 95 33
rect 86 21 95 23
rect 29 6 31 11
rect 39 6 41 11
rect 51 8 53 11
rect 86 8 88 21
rect 51 6 88 8
<< ndif >>
rect 2 20 9 30
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 16 19 19
rect 21 24 27 30
rect 21 20 29 24
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 23 11 29 16
rect 31 20 39 24
rect 31 18 34 20
rect 36 18 39 20
rect 31 11 39 18
rect 41 11 51 24
rect 53 22 58 24
rect 53 20 60 22
rect 53 18 56 20
rect 58 18 60 20
rect 53 16 60 18
rect 53 11 58 16
rect 43 9 45 11
rect 47 9 49 11
rect 43 7 49 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 31 70
rect 21 66 25 68
rect 27 66 31 68
rect 21 61 31 66
rect 21 59 25 61
rect 27 59 31 61
rect 21 42 31 59
rect 33 42 38 70
rect 40 42 45 70
rect 47 60 55 70
rect 47 58 50 60
rect 52 58 55 60
rect 47 53 55 58
rect 47 51 50 53
rect 52 51 55 53
rect 47 42 55 51
rect 57 42 62 70
rect 64 42 69 70
rect 71 58 77 70
rect 71 56 79 58
rect 71 54 74 56
rect 76 54 79 56
rect 71 42 79 54
rect 81 42 86 58
rect 88 42 93 58
rect 95 55 100 58
rect 95 53 102 55
rect 95 51 98 53
rect 100 51 102 53
rect 95 46 102 51
rect 95 44 98 46
rect 100 44 102 46
rect 95 42 102 44
<< alu1 >>
rect -2 81 106 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 106 81
rect -2 68 106 79
rect 2 46 6 55
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 13 46 17 51
rect 2 44 14 46
rect 16 44 17 46
rect 2 42 17 44
rect 2 30 6 42
rect 33 42 55 46
rect 33 39 38 42
rect 2 28 17 30
rect 2 26 14 28
rect 16 26 17 28
rect 2 25 17 26
rect 29 37 38 39
rect 29 35 30 37
rect 32 35 38 37
rect 29 33 38 35
rect 51 38 55 42
rect 51 37 79 38
rect 51 35 75 37
rect 77 35 79 37
rect 51 34 79 35
rect 89 37 102 39
rect 89 35 95 37
rect 97 35 102 37
rect 89 33 102 35
rect 42 31 46 33
rect 42 29 43 31
rect 45 30 46 31
rect 45 29 71 30
rect 42 27 64 29
rect 66 27 71 29
rect 42 26 71 27
rect 89 26 95 33
rect 13 21 17 25
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect 65 18 71 26
rect -2 11 106 12
rect -2 9 45 11
rect 47 9 106 11
rect -2 1 106 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 106 1
rect -2 -2 106 -1
<< ptie >>
rect 0 1 104 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 104 1
rect 0 -3 104 -1
<< ntie >>
rect 0 81 104 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 104 81
rect 0 77 104 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 11 31 24
rect 39 11 41 24
rect 51 11 53 24
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 31 42 33 70
rect 38 42 40 70
rect 45 42 47 70
rect 55 42 57 70
rect 62 42 64 70
rect 69 42 71 70
rect 79 42 81 58
rect 86 42 88 58
rect 93 42 95 58
<< polyct0 >>
rect 17 35 19 37
<< polyct1 >>
rect 30 35 32 37
rect 43 29 45 31
rect 75 35 77 37
rect 64 27 66 29
rect 95 35 97 37
<< ndifct0 >>
rect 4 18 6 20
rect 24 18 26 20
rect 34 18 36 20
rect 56 18 58 20
<< ndifct1 >>
rect 14 26 16 28
rect 14 19 16 21
rect 45 9 47 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 25 66 27 68
rect 25 59 27 61
rect 50 58 52 60
rect 50 51 52 53
rect 74 54 76 56
rect 98 51 100 53
rect 98 44 100 46
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 23 66 25 68
rect 27 66 29 68
rect 23 61 29 66
rect 23 59 25 61
rect 27 59 29 61
rect 23 58 29 59
rect 49 60 53 62
rect 49 58 50 60
rect 52 58 53 60
rect 49 54 53 58
rect 73 56 77 68
rect 73 54 74 56
rect 76 54 77 56
rect 21 53 67 54
rect 21 51 50 53
rect 52 51 67 53
rect 73 52 77 54
rect 96 53 102 54
rect 21 50 67 51
rect 21 38 25 50
rect 63 47 67 50
rect 96 51 98 53
rect 100 51 102 53
rect 96 47 102 51
rect 63 46 102 47
rect 63 44 98 46
rect 100 44 102 46
rect 63 43 102 44
rect 15 37 25 38
rect 15 35 17 37
rect 19 35 25 37
rect 15 34 25 35
rect 21 29 25 34
rect 21 25 36 29
rect 32 21 36 25
rect 2 20 8 21
rect 2 18 4 20
rect 6 18 8 20
rect 2 12 8 18
rect 22 20 28 21
rect 22 18 24 20
rect 26 18 28 20
rect 22 12 28 18
rect 32 20 60 21
rect 32 18 34 20
rect 36 18 56 20
rect 58 18 60 20
rect 32 17 60 18
<< labels >>
rlabel alu0 20 36 20 36 6 zn
rlabel alu0 46 19 46 19 6 zn
rlabel alu0 44 52 44 52 6 zn
rlabel alu0 51 56 51 56 6 zn
rlabel alu0 82 45 82 45 6 zn
rlabel alu0 99 48 99 48 6 zn
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 36 40 36 40 6 a
rlabel alu1 44 44 44 44 6 a
rlabel alu1 52 6 52 6 6 vss
rlabel alu1 52 28 52 28 6 b
rlabel alu1 68 36 68 36 6 a
rlabel polyct1 76 36 76 36 6 a
rlabel alu1 68 24 68 24 6 b
rlabel alu1 60 36 60 36 6 a
rlabel alu1 60 28 60 28 6 b
rlabel alu1 52 44 52 44 6 a
rlabel alu1 52 74 52 74 6 vdd
rlabel alu1 100 36 100 36 6 c
rlabel alu1 92 32 92 32 6 c
<< end >>
