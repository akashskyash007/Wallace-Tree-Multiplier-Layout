magic
tech scmos
timestamp 1199201969
<< ab >>
rect 0 0 104 80
<< nwell >>
rect -5 36 109 88
<< pwell >>
rect -5 -8 109 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 65 61 70
rect 69 61 71 65
rect 79 61 81 65
rect 89 61 91 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 41 39
rect 29 35 37 37
rect 39 35 41 37
rect 29 33 41 35
rect 29 30 31 33
rect 39 30 41 33
rect 49 39 51 42
rect 59 39 61 42
rect 49 37 61 39
rect 49 35 54 37
rect 56 35 61 37
rect 49 33 61 35
rect 49 30 51 33
rect 59 30 61 33
rect 69 39 71 42
rect 79 39 81 42
rect 89 39 91 42
rect 69 37 91 39
rect 69 35 83 37
rect 85 35 91 37
rect 69 33 91 35
rect 69 30 71 33
rect 79 30 81 33
rect 29 6 31 10
rect 39 6 41 10
rect 49 6 51 10
rect 59 6 61 10
rect 69 9 71 14
rect 79 9 81 14
<< ndif >>
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 14 29 19
rect 21 12 24 14
rect 26 12 29 14
rect 21 10 29 12
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 21 39 26
rect 31 19 34 21
rect 36 19 39 21
rect 31 10 39 19
rect 41 21 49 30
rect 41 19 44 21
rect 46 19 49 21
rect 41 14 49 19
rect 41 12 44 14
rect 46 12 49 14
rect 41 10 49 12
rect 51 28 59 30
rect 51 26 54 28
rect 56 26 59 28
rect 51 21 59 26
rect 51 19 54 21
rect 56 19 59 21
rect 51 10 59 19
rect 61 27 69 30
rect 61 25 64 27
rect 66 25 69 27
rect 61 19 69 25
rect 61 17 64 19
rect 66 17 69 19
rect 61 14 69 17
rect 71 28 79 30
rect 71 26 74 28
rect 76 26 79 28
rect 71 21 79 26
rect 71 19 74 21
rect 76 19 79 21
rect 71 14 79 19
rect 81 26 88 30
rect 81 24 84 26
rect 86 24 88 26
rect 81 18 88 24
rect 81 16 84 18
rect 86 16 88 18
rect 81 14 88 16
rect 61 10 67 14
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 42 9 52
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 60 29 66
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 53 39 70
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 60 49 66
rect 41 58 44 60
rect 46 58 49 60
rect 41 42 49 58
rect 51 65 56 70
rect 51 53 59 65
rect 51 51 54 53
rect 56 51 59 53
rect 51 46 59 51
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 61 67 65
rect 61 59 69 61
rect 61 57 64 59
rect 66 57 69 59
rect 61 52 69 57
rect 61 50 64 52
rect 66 50 69 52
rect 61 42 69 50
rect 71 53 79 61
rect 71 51 74 53
rect 76 51 79 53
rect 71 46 79 51
rect 71 44 74 46
rect 76 44 79 46
rect 71 42 79 44
rect 81 59 89 61
rect 81 57 84 59
rect 86 57 89 59
rect 81 52 89 57
rect 81 50 84 52
rect 86 50 89 52
rect 81 42 89 50
rect 91 55 96 61
rect 91 53 98 55
rect 91 51 94 53
rect 96 51 98 53
rect 91 46 98 51
rect 91 44 94 46
rect 96 44 98 46
rect 91 42 98 44
<< alu1 >>
rect -2 81 106 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 106 81
rect -2 68 106 79
rect 33 53 38 55
rect 33 51 34 53
rect 36 51 38 53
rect 33 46 38 51
rect 53 53 57 55
rect 53 51 54 53
rect 56 51 57 53
rect 53 46 57 51
rect 9 44 14 46
rect 16 44 34 46
rect 36 44 54 46
rect 56 44 57 46
rect 9 42 57 44
rect 26 30 30 42
rect 81 37 95 38
rect 81 35 83 37
rect 85 35 95 37
rect 81 34 95 35
rect 26 28 57 30
rect 26 26 34 28
rect 36 26 54 28
rect 56 26 57 28
rect 33 21 38 26
rect 33 19 34 21
rect 36 19 38 21
rect 33 17 38 19
rect 53 21 57 26
rect 53 19 54 21
rect 56 19 57 21
rect 53 17 57 19
rect 90 25 95 34
rect -2 1 106 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 106 1
rect -2 -2 106 -1
<< ptie >>
rect 0 1 104 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 104 1
rect 0 -3 104 -1
<< ntie >>
rect 0 81 104 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 104 81
rect 0 77 104 79
<< nmos >>
rect 29 10 31 30
rect 39 10 41 30
rect 49 10 51 30
rect 59 10 61 30
rect 69 14 71 30
rect 79 14 81 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 65
rect 69 42 71 61
rect 79 42 81 61
rect 89 42 91 61
<< polyct0 >>
rect 37 35 39 37
rect 54 35 56 37
<< polyct1 >>
rect 83 35 85 37
<< ndifct0 >>
rect 24 19 26 21
rect 24 12 26 14
rect 44 19 46 21
rect 44 12 46 14
rect 64 25 66 27
rect 64 17 66 19
rect 74 26 76 28
rect 74 19 76 21
rect 84 24 86 26
rect 84 16 86 18
<< ndifct1 >>
rect 34 26 36 28
rect 34 19 36 21
rect 54 26 56 28
rect 54 19 56 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 4 52 6 54
rect 14 51 16 53
rect 24 66 26 68
rect 24 58 26 60
rect 44 66 46 68
rect 44 58 46 60
rect 64 57 66 59
rect 64 50 66 52
rect 74 51 76 53
rect 74 44 76 46
rect 84 57 86 59
rect 84 50 86 52
rect 94 51 96 53
rect 94 44 96 46
<< pdifct1 >>
rect 14 44 16 46
rect 34 51 36 53
rect 34 44 36 46
rect 54 51 56 53
rect 54 44 56 46
<< alu0 >>
rect 3 66 4 68
rect 6 66 7 68
rect 3 61 7 66
rect 3 59 4 61
rect 6 59 7 61
rect 3 54 7 59
rect 23 66 24 68
rect 26 66 27 68
rect 23 60 27 66
rect 23 58 24 60
rect 26 58 27 60
rect 23 56 27 58
rect 43 66 44 68
rect 46 66 47 68
rect 43 60 47 66
rect 43 58 44 60
rect 46 58 47 60
rect 43 56 47 58
rect 62 59 68 68
rect 62 57 64 59
rect 66 57 68 59
rect 3 52 4 54
rect 6 52 7 54
rect 3 50 7 52
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 13 46 17 51
rect 62 52 68 57
rect 82 59 88 68
rect 82 57 84 59
rect 86 57 88 59
rect 62 50 64 52
rect 66 50 68 52
rect 62 49 68 50
rect 73 53 77 55
rect 73 51 74 53
rect 76 51 77 53
rect 73 46 77 51
rect 82 52 88 57
rect 82 50 84 52
rect 86 50 88 52
rect 82 49 88 50
rect 93 53 97 55
rect 93 51 94 53
rect 96 51 97 53
rect 93 46 97 51
rect 73 44 74 46
rect 76 44 94 46
rect 96 44 97 46
rect 73 42 97 44
rect 73 38 77 42
rect 35 37 77 38
rect 35 35 37 37
rect 39 35 54 37
rect 56 35 77 37
rect 35 34 77 35
rect 22 21 28 22
rect 22 19 24 21
rect 26 19 28 21
rect 22 14 28 19
rect 42 21 48 22
rect 42 19 44 21
rect 46 19 48 21
rect 22 12 24 14
rect 26 12 28 14
rect 42 14 48 19
rect 63 27 67 29
rect 63 25 64 27
rect 66 25 67 27
rect 63 19 67 25
rect 63 17 64 19
rect 66 17 67 19
rect 73 28 77 34
rect 73 26 74 28
rect 76 26 77 28
rect 73 21 77 26
rect 73 19 74 21
rect 76 19 77 21
rect 73 17 77 19
rect 83 26 87 28
rect 83 24 84 26
rect 86 24 87 26
rect 83 18 87 24
rect 42 12 44 14
rect 46 12 48 14
rect 63 12 67 17
rect 83 16 84 18
rect 86 16 87 18
rect 83 12 87 16
<< labels >>
rlabel alu0 56 36 56 36 6 an
rlabel alu0 75 36 75 36 6 an
rlabel alu0 95 48 95 48 6 an
rlabel alu1 20 44 20 44 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 44 28 44 28 6 z
rlabel alu1 36 24 36 24 6 z
rlabel alu1 44 44 44 44 6 z
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 52 6 52 6 6 vss
rlabel alu1 52 28 52 28 6 z
rlabel alu1 52 44 52 44 6 z
rlabel alu1 52 74 52 74 6 vdd
rlabel alu1 92 32 92 32 6 a
rlabel polyct1 84 36 84 36 6 a
<< end >>
