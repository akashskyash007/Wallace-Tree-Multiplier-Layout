magic
tech scmos
timestamp 1199469712
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -2 48 62 104
<< pwell >>
rect -2 -4 62 48
<< poly >>
rect 7 81 13 83
rect 7 79 9 81
rect 11 79 13 81
rect 7 77 13 79
rect 11 73 13 77
rect 23 75 25 80
rect 35 75 37 80
rect 47 73 49 78
rect 11 39 13 55
rect 23 52 25 55
rect 17 50 25 52
rect 17 48 19 50
rect 21 48 25 50
rect 17 46 29 48
rect 11 25 13 30
rect 27 24 29 46
rect 35 42 37 55
rect 47 52 49 55
rect 42 50 49 52
rect 42 48 44 50
rect 46 48 49 50
rect 42 46 49 48
rect 35 40 43 42
rect 35 38 39 40
rect 41 38 43 40
rect 35 36 43 38
rect 35 24 37 36
rect 47 33 49 46
rect 47 19 49 24
rect 27 2 29 7
rect 35 2 37 7
<< ndif >>
rect 3 34 11 39
rect 3 32 5 34
rect 7 32 11 34
rect 3 30 11 32
rect 13 37 21 39
rect 13 35 17 37
rect 19 35 21 37
rect 13 33 21 35
rect 13 30 18 33
rect 39 31 47 33
rect 39 29 41 31
rect 43 29 47 31
rect 39 24 47 29
rect 49 31 57 33
rect 49 29 53 31
rect 55 29 57 31
rect 49 27 57 29
rect 49 24 54 27
rect 19 22 27 24
rect 19 20 21 22
rect 23 20 27 22
rect 19 18 27 20
rect 22 7 27 18
rect 29 7 35 24
rect 37 21 45 24
rect 37 19 41 21
rect 43 19 45 21
rect 37 11 45 19
rect 37 9 41 11
rect 43 9 45 11
rect 37 7 45 9
<< pdif >>
rect 15 81 21 83
rect 15 79 17 81
rect 19 79 21 81
rect 39 81 45 83
rect 15 75 21 79
rect 39 79 41 81
rect 43 79 45 81
rect 39 75 45 79
rect 15 73 23 75
rect 6 61 11 73
rect 3 59 11 61
rect 3 57 5 59
rect 7 57 11 59
rect 3 55 11 57
rect 13 55 23 73
rect 25 71 35 75
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 73 45 75
rect 37 55 47 73
rect 49 61 54 73
rect 49 59 57 61
rect 49 57 53 59
rect 55 57 57 59
rect 49 55 57 57
<< alu1 >>
rect -2 95 62 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 62 95
rect -2 88 62 93
rect 8 81 12 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 73 12 79
rect 16 81 20 88
rect 16 79 17 81
rect 19 79 20 81
rect 16 77 20 79
rect 40 81 44 88
rect 40 79 41 81
rect 43 79 44 81
rect 40 77 44 79
rect 8 67 22 73
rect 4 59 8 61
rect 4 57 5 59
rect 7 57 8 59
rect 18 57 22 67
rect 28 71 32 73
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 4 51 8 57
rect 4 50 23 51
rect 4 48 19 50
rect 21 48 23 50
rect 4 47 23 48
rect 16 37 20 47
rect 4 34 8 36
rect 4 32 5 34
rect 7 32 8 34
rect 16 35 17 37
rect 19 35 20 37
rect 16 33 20 35
rect 4 12 8 32
rect 28 23 32 59
rect 38 68 53 73
rect 38 51 42 68
rect 52 59 56 61
rect 52 57 53 59
rect 55 57 56 59
rect 38 50 48 51
rect 38 48 44 50
rect 46 48 48 50
rect 38 47 48 48
rect 52 41 56 57
rect 37 40 56 41
rect 37 38 39 40
rect 41 38 56 40
rect 37 37 56 38
rect 18 22 32 23
rect 18 20 21 22
rect 23 20 32 22
rect 18 17 32 20
rect 40 31 44 33
rect 40 29 41 31
rect 43 29 44 31
rect 40 21 44 29
rect 52 31 56 37
rect 52 29 53 31
rect 55 29 56 31
rect 52 27 56 29
rect 40 19 41 21
rect 43 19 44 21
rect 40 12 44 19
rect -2 11 62 12
rect -2 9 41 11
rect 43 9 62 11
rect -2 7 62 9
rect -2 5 9 7
rect 11 5 62 7
rect -2 0 62 5
<< ptie >>
rect 7 7 13 9
rect 7 5 9 7
rect 11 5 13 7
rect 7 3 13 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 11 30 13 39
rect 47 24 49 33
rect 27 7 29 24
rect 35 7 37 24
<< pmos >>
rect 11 55 13 73
rect 23 55 25 75
rect 35 55 37 75
rect 47 55 49 73
<< polyct1 >>
rect 9 79 11 81
rect 19 48 21 50
rect 44 48 46 50
rect 39 38 41 40
<< ndifct1 >>
rect 5 32 7 34
rect 17 35 19 37
rect 41 29 43 31
rect 53 29 55 31
rect 21 20 23 22
rect 41 19 43 21
rect 41 9 43 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
<< pdifct1 >>
rect 17 79 19 81
rect 41 79 43 81
rect 5 57 7 59
rect 29 69 31 71
rect 29 59 31 61
rect 53 57 55 59
<< labels >>
rlabel alu1 6 54 6 54 6 bn
rlabel alu1 10 75 10 75 6 b
rlabel alu1 20 20 20 20 6 z
rlabel alu1 18 42 18 42 6 bn
rlabel alu1 13 49 13 49 6 bn
rlabel alu1 20 65 20 65 6 b
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 30 45 30 45 6 z
rlabel alu1 40 60 40 60 6 a
rlabel alu1 30 94 30 94 6 vdd
rlabel alu1 46 39 46 39 6 an
rlabel alu1 54 44 54 44 6 an
rlabel alu1 50 70 50 70 6 a
<< end >>
