magic
tech scmos
timestamp 1199203569
<< ab >>
rect 0 0 200 80
<< nwell >>
rect -5 36 205 88
<< pwell >>
rect -5 -8 205 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 79 70 81 74
rect 89 70 91 74
rect 99 70 101 74
rect 109 70 111 74
rect 119 70 121 74
rect 126 70 128 74
rect 136 70 138 74
rect 143 70 145 74
rect 153 70 155 74
rect 160 70 162 74
rect 170 70 172 74
rect 177 70 179 74
rect 79 47 81 50
rect 89 47 91 50
rect 99 47 101 50
rect 79 45 101 47
rect 79 43 81 45
rect 83 43 85 45
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 31 39
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 41 85 43
rect 99 43 101 45
rect 109 43 111 46
rect 99 41 111 43
rect 79 39 81 41
rect 39 37 64 39
rect 9 30 11 37
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 58 35 60 37
rect 62 35 64 37
rect 58 33 64 35
rect 19 30 21 33
rect 42 29 44 33
rect 52 29 54 33
rect 62 29 64 33
rect 69 37 81 39
rect 69 29 71 37
rect 79 29 81 37
rect 89 38 95 40
rect 89 36 91 38
rect 93 36 95 38
rect 119 37 121 42
rect 126 39 128 42
rect 136 39 138 42
rect 126 37 138 39
rect 143 39 145 42
rect 153 39 155 42
rect 143 37 155 39
rect 86 34 95 36
rect 114 35 121 37
rect 86 29 88 34
rect 114 33 116 35
rect 118 33 121 35
rect 129 35 131 37
rect 133 35 135 37
rect 129 33 135 35
rect 114 31 121 33
rect 133 27 135 33
rect 143 35 147 37
rect 149 35 155 37
rect 143 33 155 35
rect 160 39 162 42
rect 170 39 172 42
rect 160 37 172 39
rect 160 35 163 37
rect 165 35 167 37
rect 160 33 167 35
rect 143 27 145 33
rect 153 27 155 33
rect 163 27 165 33
rect 177 31 179 42
rect 177 29 183 31
rect 177 27 179 29
rect 181 27 183 29
rect 9 10 11 13
rect 19 10 21 13
rect 42 10 44 13
rect 52 10 54 13
rect 9 8 54 10
rect 62 8 64 13
rect 69 8 71 13
rect 79 8 81 13
rect 86 8 88 13
rect 177 25 183 27
rect 133 6 135 10
rect 143 6 145 10
rect 153 6 155 10
rect 163 6 165 10
<< ndif >>
rect 2 25 9 30
rect 2 23 4 25
rect 6 23 9 25
rect 2 17 9 23
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 13 19 19
rect 21 17 29 30
rect 21 15 24 17
rect 26 15 29 17
rect 35 27 42 29
rect 35 25 37 27
rect 39 25 42 27
rect 35 20 42 25
rect 35 18 37 20
rect 39 18 42 20
rect 35 16 42 18
rect 21 13 29 15
rect 37 13 42 16
rect 44 27 52 29
rect 44 25 47 27
rect 49 25 52 27
rect 44 13 52 25
rect 54 27 62 29
rect 54 25 57 27
rect 59 25 62 27
rect 54 20 62 25
rect 54 18 57 20
rect 59 18 62 20
rect 54 13 62 18
rect 64 13 69 29
rect 71 17 79 29
rect 71 15 74 17
rect 76 15 79 17
rect 71 13 79 15
rect 81 13 86 29
rect 88 27 95 29
rect 88 25 91 27
rect 93 25 95 27
rect 88 20 95 25
rect 88 18 91 20
rect 93 18 95 20
rect 88 16 95 18
rect 124 21 133 27
rect 124 19 127 21
rect 129 19 133 21
rect 88 13 93 16
rect 124 14 133 19
rect 124 12 127 14
rect 129 12 133 14
rect 124 10 133 12
rect 135 21 143 27
rect 135 19 138 21
rect 140 19 143 21
rect 135 10 143 19
rect 145 14 153 27
rect 145 12 148 14
rect 150 12 153 14
rect 145 10 153 12
rect 155 21 163 27
rect 155 19 158 21
rect 160 19 163 21
rect 155 10 163 19
rect 165 14 173 27
rect 165 12 168 14
rect 170 12 173 14
rect 165 10 173 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 54 19 70
rect 11 52 14 54
rect 16 52 19 54
rect 11 47 19 52
rect 11 45 14 47
rect 16 45 19 47
rect 11 42 19 45
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 42 39 52
rect 41 62 49 70
rect 41 60 44 62
rect 46 60 49 62
rect 41 46 49 60
rect 41 44 44 46
rect 46 44 49 46
rect 41 42 49 44
rect 51 53 59 70
rect 51 51 54 53
rect 56 51 59 53
rect 51 46 59 51
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 62 69 70
rect 61 60 64 62
rect 66 60 69 62
rect 61 55 69 60
rect 61 53 64 55
rect 66 53 69 55
rect 61 42 69 53
rect 71 54 79 70
rect 71 52 74 54
rect 76 52 79 54
rect 71 50 79 52
rect 81 62 89 70
rect 81 60 84 62
rect 86 60 89 62
rect 81 50 89 60
rect 91 54 99 70
rect 91 52 94 54
rect 96 52 99 54
rect 91 50 99 52
rect 101 62 109 70
rect 101 60 104 62
rect 106 60 109 62
rect 101 50 109 60
rect 71 42 76 50
rect 104 46 109 50
rect 111 61 119 70
rect 111 59 114 61
rect 116 59 119 61
rect 111 54 119 59
rect 111 52 114 54
rect 116 52 119 54
rect 111 46 119 52
rect 114 42 119 46
rect 121 42 126 70
rect 128 68 136 70
rect 128 66 131 68
rect 133 66 136 68
rect 128 61 136 66
rect 128 59 131 61
rect 133 59 136 61
rect 128 42 136 59
rect 138 42 143 70
rect 145 61 153 70
rect 145 59 148 61
rect 150 59 153 61
rect 145 54 153 59
rect 145 52 148 54
rect 150 52 153 54
rect 145 42 153 52
rect 155 42 160 70
rect 162 68 170 70
rect 162 66 165 68
rect 167 66 170 68
rect 162 61 170 66
rect 162 59 165 61
rect 167 59 170 61
rect 162 42 170 59
rect 172 42 177 70
rect 179 55 184 70
rect 179 53 186 55
rect 179 51 182 53
rect 184 51 186 53
rect 179 46 186 51
rect 179 44 182 46
rect 184 44 186 46
rect 179 42 186 44
<< alu1 >>
rect -2 81 202 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 202 81
rect -2 68 202 79
rect 26 39 30 47
rect 18 37 30 39
rect 18 35 21 37
rect 23 35 30 37
rect 18 33 30 35
rect 26 25 30 33
rect 34 46 48 47
rect 34 44 44 46
rect 46 44 48 46
rect 34 42 48 44
rect 34 27 38 42
rect 129 42 167 46
rect 113 35 119 38
rect 34 25 37 27
rect 34 21 38 25
rect 113 33 116 35
rect 118 33 119 35
rect 129 37 135 42
rect 129 35 131 37
rect 133 35 135 37
rect 129 34 135 35
rect 113 30 119 33
rect 146 37 150 38
rect 146 35 147 37
rect 149 35 150 37
rect 146 30 150 35
rect 161 37 167 42
rect 161 35 163 37
rect 165 35 167 37
rect 161 34 167 35
rect 56 27 95 30
rect 56 25 57 27
rect 59 26 91 27
rect 59 25 61 26
rect 56 21 61 25
rect 34 20 61 21
rect 34 18 37 20
rect 39 18 57 20
rect 59 18 61 20
rect 89 25 91 26
rect 93 25 95 27
rect 89 20 95 25
rect 34 17 61 18
rect 89 18 91 20
rect 93 18 95 20
rect 113 29 183 30
rect 113 27 179 29
rect 181 27 183 29
rect 113 26 183 27
rect 113 18 119 26
rect 89 17 95 18
rect -2 1 202 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 202 1
rect -2 -2 202 -1
<< ptie >>
rect 0 1 200 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 171 1
rect 173 -1 179 1
rect 181 -1 187 1
rect 189 -1 195 1
rect 197 -1 200 1
rect 0 -3 200 -1
<< ntie >>
rect 0 81 200 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 171 81
rect 173 79 179 81
rect 181 79 187 81
rect 189 79 195 81
rect 197 79 200 81
rect 0 77 200 79
<< nmos >>
rect 9 13 11 30
rect 19 13 21 30
rect 42 13 44 29
rect 52 13 54 29
rect 62 13 64 29
rect 69 13 71 29
rect 79 13 81 29
rect 86 13 88 29
rect 133 10 135 27
rect 143 10 145 27
rect 153 10 155 27
rect 163 10 165 27
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 79 50 81 70
rect 89 50 91 70
rect 99 50 101 70
rect 109 46 111 70
rect 119 42 121 70
rect 126 42 128 70
rect 136 42 138 70
rect 143 42 145 70
rect 153 42 155 70
rect 160 42 162 70
rect 170 42 172 70
rect 177 42 179 70
<< polyct0 >>
rect 81 43 83 45
rect 60 35 62 37
rect 91 36 93 38
<< polyct1 >>
rect 21 35 23 37
rect 116 33 118 35
rect 131 35 133 37
rect 147 35 149 37
rect 163 35 165 37
rect 179 27 181 29
<< ndifct0 >>
rect 4 23 6 25
rect 4 15 6 17
rect 14 26 16 28
rect 14 19 16 21
rect 24 15 26 17
rect 38 25 39 27
rect 47 25 49 27
rect 74 15 76 17
rect 127 19 129 21
rect 127 12 129 14
rect 138 19 140 21
rect 148 12 150 14
rect 158 19 160 21
rect 168 12 170 14
<< ndifct1 >>
rect 37 25 38 27
rect 37 18 39 20
rect 57 25 59 27
rect 57 18 59 20
rect 91 25 93 27
rect 91 18 93 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
rect 171 79 173 81
rect 179 79 181 81
rect 187 79 189 81
rect 195 79 197 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
rect 171 -1 173 1
rect 179 -1 181 1
rect 187 -1 189 1
rect 195 -1 197 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 52 16 54
rect 14 45 16 47
rect 24 66 26 68
rect 24 59 26 61
rect 34 59 36 61
rect 34 52 36 54
rect 44 60 46 62
rect 54 51 56 53
rect 54 44 56 46
rect 64 60 66 62
rect 64 53 66 55
rect 74 52 76 54
rect 84 60 86 62
rect 94 52 96 54
rect 104 60 106 62
rect 114 59 116 61
rect 114 52 116 54
rect 131 66 133 68
rect 131 59 133 61
rect 148 59 150 61
rect 148 52 150 54
rect 165 66 167 68
rect 165 59 167 61
rect 182 51 184 53
rect 182 44 184 46
<< pdifct1 >>
rect 44 44 46 46
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 129 66 131 68
rect 133 66 135 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 33 61 37 63
rect 33 59 34 61
rect 36 59 37 61
rect 42 62 108 63
rect 42 60 44 62
rect 46 60 64 62
rect 66 60 84 62
rect 86 60 104 62
rect 106 60 108 62
rect 42 59 108 60
rect 113 61 117 63
rect 113 59 114 61
rect 116 59 117 61
rect 33 55 37 59
rect 63 55 67 59
rect 113 55 117 59
rect 129 61 135 66
rect 163 66 165 68
rect 167 66 169 68
rect 129 59 131 61
rect 133 59 135 61
rect 129 58 135 59
rect 147 61 151 63
rect 147 59 148 61
rect 150 59 151 61
rect 147 55 151 59
rect 163 61 169 66
rect 163 59 165 61
rect 167 59 169 61
rect 189 59 193 68
rect 163 58 169 59
rect 12 54 57 55
rect 12 52 14 54
rect 16 52 34 54
rect 36 53 57 54
rect 36 52 54 53
rect 12 51 54 52
rect 56 51 57 53
rect 63 53 64 55
rect 66 53 67 55
rect 63 51 67 53
rect 72 54 185 55
rect 72 52 74 54
rect 76 52 94 54
rect 96 52 114 54
rect 116 52 148 54
rect 150 53 185 54
rect 150 52 182 53
rect 72 51 182 52
rect 184 51 185 53
rect 12 47 17 51
rect 10 45 14 47
rect 16 45 17 47
rect 10 43 17 45
rect 10 29 14 43
rect 10 28 18 29
rect 3 25 7 27
rect 10 26 14 28
rect 16 26 18 28
rect 10 25 18 26
rect 53 46 57 51
rect 53 44 54 46
rect 56 45 85 46
rect 56 44 81 45
rect 53 43 81 44
rect 83 43 85 45
rect 53 42 85 43
rect 90 38 94 51
rect 181 46 185 51
rect 181 44 182 46
rect 184 44 190 46
rect 181 42 190 44
rect 45 37 91 38
rect 45 35 60 37
rect 62 36 91 37
rect 93 36 94 38
rect 62 35 94 36
rect 45 34 94 35
rect 38 27 40 29
rect 39 25 40 27
rect 3 23 4 25
rect 6 23 7 25
rect 3 17 7 23
rect 12 21 18 25
rect 12 19 14 21
rect 16 19 18 21
rect 38 21 40 25
rect 45 27 51 34
rect 145 30 146 38
rect 150 30 151 38
rect 45 25 47 27
rect 49 25 51 27
rect 45 24 51 25
rect 12 18 18 19
rect 3 15 4 17
rect 6 15 7 17
rect 3 12 7 15
rect 23 17 27 19
rect 73 17 77 19
rect 126 21 130 23
rect 186 22 190 42
rect 126 19 127 21
rect 129 19 130 21
rect 23 15 24 17
rect 26 15 27 17
rect 23 12 27 15
rect 73 15 74 17
rect 76 15 77 17
rect 73 12 77 15
rect 126 14 130 19
rect 136 21 190 22
rect 136 19 138 21
rect 140 19 158 21
rect 160 19 190 21
rect 136 18 190 19
rect 126 12 127 14
rect 129 12 130 14
rect 146 14 152 15
rect 146 12 148 14
rect 150 12 152 14
rect 166 14 172 15
rect 166 12 168 14
rect 170 12 172 14
<< labels >>
rlabel alu0 15 23 15 23 6 bn
rlabel alu0 14 49 14 49 6 bn
rlabel alu0 35 57 35 57 6 bn
rlabel alu0 48 31 48 31 6 an
rlabel alu0 55 48 55 48 6 bn
rlabel alu0 34 53 34 53 6 bn
rlabel alu0 69 44 69 44 6 bn
rlabel alu0 115 57 115 57 6 an
rlabel alu0 149 57 149 57 6 an
rlabel alu0 163 20 163 20 6 an
rlabel alu0 183 48 183 48 6 an
rlabel alu0 128 53 128 53 6 an
rlabel alu1 20 36 20 36 6 b
rlabel alu1 28 36 28 36 6 b
rlabel alu1 60 28 60 28 6 z
rlabel alu1 68 28 68 28 6 z
rlabel alu1 76 28 76 28 6 z
rlabel alu1 36 32 36 32 6 z
rlabel alu1 44 44 44 44 6 z
rlabel alu1 100 6 100 6 6 vss
rlabel alu1 116 28 116 28 6 a2
rlabel alu1 84 28 84 28 6 z
rlabel alu1 92 24 92 24 6 z
rlabel alu1 100 74 100 74 6 vdd
rlabel alu1 124 28 124 28 6 a2
rlabel alu1 132 28 132 28 6 a2
rlabel alu1 140 28 140 28 6 a2
rlabel alu1 156 28 156 28 6 a2
rlabel alu1 148 32 148 32 6 a2
rlabel alu1 132 40 132 40 6 a1
rlabel alu1 140 44 140 44 6 a1
rlabel alu1 148 44 148 44 6 a1
rlabel alu1 156 44 156 44 6 a1
rlabel alu1 164 28 164 28 6 a2
rlabel alu1 172 28 172 28 6 a2
rlabel polyct1 180 28 180 28 6 a2
rlabel alu1 164 40 164 40 6 a1
rlabel alu1 164 44 164 44 6 a1
<< end >>
