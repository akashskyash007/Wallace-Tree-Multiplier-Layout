magic
tech scmos
timestamp 1199202389
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 10 66 12 71
rect 20 58 22 63
rect 10 39 12 42
rect 20 39 22 42
rect 9 37 23 39
rect 9 35 19 37
rect 21 35 23 37
rect 9 33 23 35
rect 9 30 11 33
rect 9 10 11 15
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 15 9 17
rect 11 27 19 30
rect 11 25 14 27
rect 16 25 19 27
rect 11 19 19 25
rect 11 17 14 19
rect 16 17 19 19
rect 11 15 19 17
<< pdif >>
rect 2 64 10 66
rect 2 62 5 64
rect 7 62 10 64
rect 2 56 10 62
rect 2 54 5 56
rect 7 54 10 56
rect 2 42 10 54
rect 12 58 17 66
rect 12 53 20 58
rect 12 51 15 53
rect 17 51 20 53
rect 12 46 20 51
rect 12 44 15 46
rect 17 44 20 46
rect 12 42 20 44
rect 22 56 30 58
rect 22 54 25 56
rect 27 54 30 56
rect 22 42 30 54
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 41 14 47
rect 2 30 6 41
rect 26 39 30 47
rect 18 37 30 39
rect 18 35 19 37
rect 21 35 30 37
rect 18 33 30 35
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 15 11 30
<< pmos >>
rect 10 42 12 66
rect 20 42 22 58
<< polyct1 >>
rect 19 35 21 37
<< ndifct0 >>
rect 14 25 16 27
rect 14 17 16 19
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 5 62 7 64
rect 5 54 7 56
rect 15 51 17 53
rect 15 44 17 46
rect 25 54 27 56
<< alu0 >>
rect 4 64 8 68
rect 4 62 5 64
rect 7 62 8 64
rect 4 56 8 62
rect 4 54 5 56
rect 7 54 8 56
rect 24 56 28 68
rect 24 54 25 56
rect 27 54 28 56
rect 4 52 8 54
rect 13 53 19 54
rect 13 51 15 53
rect 17 51 19 53
rect 24 52 28 54
rect 13 47 19 51
rect 14 46 19 47
rect 14 44 15 46
rect 17 44 19 46
rect 14 43 19 44
rect 13 27 17 29
rect 13 25 14 27
rect 16 25 17 27
rect 13 19 17 25
rect 13 17 14 19
rect 16 17 17 19
rect 13 12 17 17
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 12 44 12 44 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel polyct1 20 36 20 36 6 a
rlabel alu1 28 40 28 40 6 a
<< end >>
