magic
tech scmos
timestamp 1199202256
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 9 35 11 38
rect 19 35 21 38
rect 9 33 22 35
rect 9 31 18 33
rect 20 31 22 33
rect 9 29 22 31
rect 9 26 11 29
rect 19 26 21 29
rect 19 10 21 15
rect 9 4 11 9
<< ndif >>
rect 2 13 9 26
rect 2 11 4 13
rect 6 11 9 13
rect 2 9 9 11
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 15 19 22
rect 21 20 29 26
rect 21 18 24 20
rect 26 18 29 20
rect 21 15 29 18
rect 11 9 16 15
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
<< alu1 >>
rect -2 64 34 72
rect 2 48 14 50
rect 16 48 23 50
rect 2 46 23 48
rect 2 25 6 46
rect 17 35 23 42
rect 17 33 30 35
rect 17 31 18 33
rect 20 31 30 33
rect 17 29 30 31
rect 2 24 18 25
rect 2 22 14 24
rect 16 22 18 24
rect 2 21 18 22
rect -2 7 34 8
rect -2 5 25 7
rect 27 5 34 7
rect -2 0 34 5
<< ptie >>
rect 23 7 29 9
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< nmos >>
rect 9 9 11 26
rect 19 15 21 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
<< polyct1 >>
rect 18 31 20 33
<< ndifct0 >>
rect 4 11 6 13
rect 24 18 26 20
<< ndifct1 >>
rect 14 22 16 24
<< ptiect1 >>
rect 25 5 27 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 55 16 57
rect 24 62 26 64
rect 24 55 26 57
<< pdifct1 >>
rect 14 48 16 50
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 50 17 55
rect 22 57 28 62
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 23 20 27 22
rect 23 18 24 20
rect 26 18 27 20
rect 3 13 7 15
rect 3 11 4 13
rect 6 11 7 13
rect 3 8 7 11
rect 23 8 27 18
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 20 48 20 48 6 z
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 32 28 32 6 a
<< end >>
