magic
tech scmos
timestamp 1199203016
<< ab >>
rect 0 0 88 72
<< nwell >>
rect -5 32 93 77
<< pwell >>
rect -5 -5 93 32
<< poly >>
rect 11 66 13 70
rect 18 66 20 70
rect 25 66 27 70
rect 35 66 37 70
rect 42 66 44 70
rect 49 66 51 70
rect 59 66 61 70
rect 66 66 68 70
rect 73 66 75 70
rect 11 30 13 39
rect 18 36 20 39
rect 25 36 27 39
rect 35 36 37 39
rect 18 34 21 36
rect 25 34 37 36
rect 19 30 21 34
rect 29 33 35 34
rect 29 31 31 33
rect 33 31 35 33
rect 9 28 15 30
rect 9 26 11 28
rect 13 26 15 28
rect 9 24 15 26
rect 19 28 25 30
rect 19 26 21 28
rect 23 26 25 28
rect 19 24 25 26
rect 29 29 35 31
rect 9 21 11 24
rect 19 21 21 24
rect 29 21 31 29
rect 42 26 44 39
rect 49 36 51 39
rect 59 36 61 39
rect 49 34 62 36
rect 56 32 58 34
rect 60 32 62 34
rect 56 30 62 32
rect 66 26 68 39
rect 42 24 68 26
rect 73 27 75 39
rect 73 25 79 27
rect 42 17 48 24
rect 73 23 75 25
rect 77 23 79 25
rect 73 21 79 23
rect 42 15 44 17
rect 46 15 48 17
rect 42 13 48 15
rect 9 2 11 6
rect 19 2 21 6
rect 29 2 31 6
<< ndif >>
rect 4 19 9 21
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 6 9 13
rect 11 10 19 21
rect 11 8 14 10
rect 16 8 19 10
rect 11 6 19 8
rect 21 17 29 21
rect 21 15 24 17
rect 26 15 29 17
rect 21 6 29 15
rect 31 17 39 21
rect 31 15 34 17
rect 36 15 39 17
rect 31 10 39 15
rect 31 8 34 10
rect 36 8 39 10
rect 31 6 39 8
<< pdif >>
rect 6 58 11 66
rect 4 56 11 58
rect 4 54 6 56
rect 8 54 11 56
rect 4 49 11 54
rect 4 47 6 49
rect 8 47 11 49
rect 4 45 11 47
rect 6 39 11 45
rect 13 39 18 66
rect 20 39 25 66
rect 27 64 35 66
rect 27 62 30 64
rect 32 62 35 64
rect 27 57 35 62
rect 27 55 30 57
rect 32 55 35 57
rect 27 39 35 55
rect 37 39 42 66
rect 44 39 49 66
rect 51 57 59 66
rect 51 55 54 57
rect 56 55 59 57
rect 51 50 59 55
rect 51 48 54 50
rect 56 48 59 50
rect 51 39 59 48
rect 61 39 66 66
rect 68 39 73 66
rect 75 64 82 66
rect 75 62 78 64
rect 80 62 82 64
rect 75 57 82 62
rect 75 55 78 57
rect 80 55 82 57
rect 75 39 82 55
<< alu1 >>
rect -2 64 90 72
rect 2 50 6 51
rect 2 49 54 50
rect 2 47 6 49
rect 8 48 54 49
rect 56 48 63 50
rect 8 47 63 48
rect 2 46 63 47
rect 2 18 6 46
rect 10 38 63 42
rect 10 28 14 38
rect 57 34 63 38
rect 29 33 53 34
rect 29 31 31 33
rect 33 31 53 33
rect 29 30 53 31
rect 57 32 58 34
rect 60 32 63 34
rect 57 30 63 32
rect 10 26 11 28
rect 13 26 14 28
rect 10 24 14 26
rect 20 28 24 30
rect 20 26 21 28
rect 23 26 24 28
rect 49 26 53 30
rect 20 22 45 26
rect 49 25 79 26
rect 49 23 75 25
rect 77 23 79 25
rect 49 22 79 23
rect 41 18 45 22
rect 2 17 28 18
rect 2 15 4 17
rect 6 15 24 17
rect 26 15 28 17
rect 2 14 28 15
rect 41 17 55 18
rect 41 15 44 17
rect 46 15 55 17
rect 41 14 55 15
rect -2 7 90 8
rect -2 5 69 7
rect 71 5 77 7
rect 79 5 90 7
rect -2 0 90 5
<< ptie >>
rect 67 7 81 18
rect 67 5 69 7
rect 71 5 77 7
rect 79 5 81 7
rect 67 3 81 5
<< nmos >>
rect 9 6 11 21
rect 19 6 21 21
rect 29 6 31 21
<< pmos >>
rect 11 39 13 66
rect 18 39 20 66
rect 25 39 27 66
rect 35 39 37 66
rect 42 39 44 66
rect 49 39 51 66
rect 59 39 61 66
rect 66 39 68 66
rect 73 39 75 66
<< polyct1 >>
rect 31 31 33 33
rect 11 26 13 28
rect 21 26 23 28
rect 58 32 60 34
rect 75 23 77 25
rect 44 15 46 17
<< ndifct0 >>
rect 14 8 16 10
rect 34 15 36 17
rect 34 8 36 10
<< ndifct1 >>
rect 4 15 6 17
rect 24 15 26 17
<< ptiect1 >>
rect 69 5 71 7
rect 77 5 79 7
<< pdifct0 >>
rect 6 54 8 56
rect 30 62 32 64
rect 30 55 32 57
rect 54 55 56 57
rect 78 62 80 64
rect 78 55 80 57
<< pdifct1 >>
rect 6 47 8 49
rect 54 48 56 50
<< alu0 >>
rect 28 62 30 64
rect 32 62 34 64
rect 5 56 9 58
rect 5 54 6 56
rect 8 54 9 56
rect 28 57 34 62
rect 76 62 78 64
rect 80 62 82 64
rect 28 55 30 57
rect 32 55 34 57
rect 28 54 34 55
rect 53 57 57 59
rect 53 55 54 57
rect 56 55 57 57
rect 5 51 9 54
rect 6 50 9 51
rect 53 50 57 55
rect 76 57 82 62
rect 76 55 78 57
rect 80 55 82 57
rect 76 54 82 55
rect 32 17 38 18
rect 32 15 34 17
rect 36 15 38 17
rect 12 10 18 11
rect 12 8 14 10
rect 16 8 18 10
rect 32 10 38 15
rect 32 8 34 10
rect 36 8 38 10
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel alu1 12 32 12 32 6 c
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 24 28 24 6 b
rlabel alu1 20 40 20 40 6 c
rlabel alu1 28 40 28 40 6 c
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 44 4 44 4 6 vss
rlabel alu1 44 16 44 16 6 b
rlabel alu1 36 24 36 24 6 b
rlabel alu1 44 32 44 32 6 a
rlabel alu1 36 32 36 32 6 a
rlabel alu1 36 40 36 40 6 c
rlabel alu1 44 40 44 40 6 c
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 44 68 44 68 6 vdd
rlabel alu1 52 16 52 16 6 b
rlabel alu1 52 24 52 24 6 a
rlabel alu1 60 24 60 24 6 a
rlabel alu1 68 24 68 24 6 a
rlabel alu1 52 40 52 40 6 c
rlabel alu1 60 36 60 36 6 c
rlabel alu1 52 48 52 48 6 z
rlabel alu1 60 48 60 48 6 z
rlabel polyct1 76 24 76 24 6 a
<< end >>
