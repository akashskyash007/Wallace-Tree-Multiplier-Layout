magic
tech scmos
timestamp 1199203124
<< ab >>
rect 0 0 104 72
<< nwell >>
rect -5 32 109 77
<< pwell >>
rect -5 -5 109 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 36 66 38 70
rect 46 66 48 70
rect 53 66 55 70
rect 63 66 65 70
rect 70 66 72 70
rect 80 58 82 63
rect 87 58 89 63
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 33 21 35
rect 9 31 11 33
rect 13 31 21 33
rect 9 29 21 31
rect 25 33 31 35
rect 25 31 27 33
rect 29 31 31 33
rect 25 29 31 31
rect 36 29 38 38
rect 46 29 48 38
rect 53 35 55 38
rect 63 35 65 38
rect 70 35 72 38
rect 80 35 82 38
rect 53 33 65 35
rect 69 33 82 35
rect 87 35 89 38
rect 87 33 95 35
rect 55 31 57 33
rect 59 31 61 33
rect 55 29 61 31
rect 9 26 11 29
rect 19 26 21 29
rect 36 27 51 29
rect 39 24 41 27
rect 49 24 51 27
rect 59 24 61 29
rect 69 31 71 33
rect 73 31 75 33
rect 69 29 75 31
rect 87 31 91 33
rect 93 31 95 33
rect 87 29 95 31
rect 69 24 71 29
rect 79 27 95 29
rect 79 24 81 27
rect 91 24 93 27
rect 29 18 31 23
rect 59 8 61 12
rect 9 2 11 7
rect 19 4 21 7
rect 29 4 31 7
rect 19 2 31 4
rect 39 2 41 7
rect 49 4 51 7
rect 69 4 71 12
rect 49 2 71 4
rect 79 2 81 7
rect 91 2 93 7
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 7 9 13
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 7 19 22
rect 21 18 26 26
rect 34 18 39 24
rect 21 16 29 18
rect 21 14 24 16
rect 26 14 29 16
rect 21 7 29 14
rect 31 16 39 18
rect 31 14 34 16
rect 36 14 39 16
rect 31 7 39 14
rect 41 11 49 24
rect 41 9 44 11
rect 46 9 49 11
rect 41 7 49 9
rect 51 21 59 24
rect 51 19 54 21
rect 56 19 59 21
rect 51 12 59 19
rect 61 16 69 24
rect 61 14 64 16
rect 66 14 69 16
rect 61 12 69 14
rect 71 21 79 24
rect 71 19 74 21
rect 76 19 79 21
rect 71 12 79 19
rect 51 7 56 12
rect 74 7 79 12
rect 81 7 91 24
rect 93 18 98 24
rect 93 16 100 18
rect 93 14 96 16
rect 98 14 100 16
rect 93 12 100 14
rect 93 7 98 12
rect 83 5 85 7
rect 87 5 89 7
rect 83 3 89 5
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 56 19 66
rect 11 54 14 56
rect 16 54 19 56
rect 11 49 19 54
rect 11 47 14 49
rect 16 47 19 49
rect 11 38 19 47
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 38 36 66
rect 38 56 46 66
rect 38 54 41 56
rect 43 54 46 56
rect 38 49 46 54
rect 38 47 41 49
rect 43 47 46 49
rect 38 38 46 47
rect 48 38 53 66
rect 55 64 63 66
rect 55 62 58 64
rect 60 62 63 64
rect 55 57 63 62
rect 55 55 58 57
rect 60 55 63 57
rect 55 38 63 55
rect 65 38 70 66
rect 72 58 77 66
rect 72 56 80 58
rect 72 54 75 56
rect 77 54 80 56
rect 72 49 80 54
rect 72 47 75 49
rect 77 47 80 49
rect 72 38 80 47
rect 82 38 87 58
rect 89 56 97 58
rect 89 54 92 56
rect 94 54 97 56
rect 89 49 97 54
rect 89 47 92 49
rect 94 47 97 49
rect 89 38 97 47
<< alu1 >>
rect -2 67 106 72
rect -2 65 97 67
rect 99 65 106 67
rect -2 64 106 65
rect 40 56 46 59
rect 40 54 41 56
rect 43 54 46 56
rect 73 56 79 59
rect 73 54 75 56
rect 77 54 79 56
rect 40 50 46 54
rect 73 50 79 54
rect 2 49 79 50
rect 2 47 14 49
rect 16 47 41 49
rect 43 47 75 49
rect 77 47 79 49
rect 2 46 79 47
rect 2 24 6 46
rect 10 38 23 42
rect 57 38 95 42
rect 10 33 14 38
rect 57 34 61 38
rect 10 31 11 33
rect 13 31 14 33
rect 10 29 14 31
rect 25 33 61 34
rect 25 31 27 33
rect 29 31 57 33
rect 59 31 61 33
rect 25 30 61 31
rect 65 33 85 34
rect 65 31 71 33
rect 73 31 85 33
rect 65 30 85 31
rect 89 33 95 38
rect 89 31 91 33
rect 93 31 95 33
rect 89 30 95 31
rect 81 26 85 30
rect 2 22 4 24
rect 2 17 6 22
rect 81 22 95 26
rect 2 15 4 17
rect 6 16 28 17
rect 6 15 24 16
rect 2 14 24 15
rect 26 14 28 16
rect 2 13 28 14
rect -2 7 106 8
rect -2 5 85 7
rect 87 5 106 7
rect -2 0 106 5
<< ntie >>
rect 95 67 101 69
rect 95 65 97 67
rect 99 65 101 67
rect 95 63 101 65
<< nmos >>
rect 9 7 11 26
rect 19 7 21 26
rect 29 7 31 18
rect 39 7 41 24
rect 49 7 51 24
rect 59 12 61 24
rect 69 12 71 24
rect 79 7 81 24
rect 91 7 93 24
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 36 38 38 66
rect 46 38 48 66
rect 53 38 55 66
rect 63 38 65 66
rect 70 38 72 66
rect 80 38 82 58
rect 87 38 89 58
<< polyct1 >>
rect 11 31 13 33
rect 27 31 29 33
rect 57 31 59 33
rect 71 31 73 33
rect 91 31 93 33
<< ndifct0 >>
rect 14 22 16 24
rect 34 14 36 16
rect 44 9 46 11
rect 54 19 56 21
rect 64 14 66 16
rect 74 19 76 21
rect 96 14 98 16
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
rect 24 14 26 16
rect 85 5 87 7
<< ntiect1 >>
rect 97 65 99 67
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 54 16 56
rect 24 62 26 64
rect 24 55 26 57
rect 58 62 60 64
rect 58 55 60 57
rect 92 54 94 56
rect 92 47 94 49
<< pdifct1 >>
rect 14 47 16 49
rect 41 54 43 56
rect 41 47 43 49
rect 75 54 77 56
rect 75 47 77 49
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 56 17 58
rect 13 54 14 56
rect 16 54 17 56
rect 22 57 28 62
rect 56 62 58 64
rect 60 62 62 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 56 57 62 62
rect 56 55 58 57
rect 60 55 62 57
rect 56 54 62 55
rect 13 50 17 54
rect 90 56 96 64
rect 90 54 92 56
rect 94 54 96 56
rect 90 49 96 54
rect 90 47 92 49
rect 94 47 96 49
rect 90 46 96 47
rect 6 17 8 25
rect 12 24 77 25
rect 12 22 14 24
rect 16 22 77 24
rect 12 21 77 22
rect 32 16 38 21
rect 53 19 54 21
rect 56 19 57 21
rect 53 17 57 19
rect 73 19 74 21
rect 76 19 77 21
rect 73 17 77 19
rect 32 14 34 16
rect 36 14 38 16
rect 32 13 38 14
rect 62 16 68 17
rect 62 14 64 16
rect 66 14 68 16
rect 43 11 47 13
rect 43 9 44 11
rect 46 9 47 11
rect 43 8 47 9
rect 62 8 68 14
rect 73 16 100 17
rect 73 14 96 16
rect 98 14 100 16
rect 73 13 100 14
<< labels >>
rlabel alu0 35 19 35 19 6 n1
rlabel alu0 86 15 86 15 6 n1
rlabel alu0 75 19 75 19 6 n1
rlabel alu0 44 23 44 23 6 n1
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 36 32 36 32 6 a1
rlabel polyct1 28 32 28 32 6 a1
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 52 4 52 4 6 vss
rlabel alu1 52 32 52 32 6 a1
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 60 40 60 40 6 a1
rlabel alu1 44 52 44 52 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 52 68 52 68 6 vdd
rlabel alu1 76 32 76 32 6 a2
rlabel alu1 68 32 68 32 6 a2
rlabel alu1 76 40 76 40 6 a1
rlabel alu1 68 40 68 40 6 a1
rlabel alu1 76 52 76 52 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 84 24 84 24 6 a2
rlabel alu1 92 24 92 24 6 a2
rlabel alu1 84 40 84 40 6 a1
rlabel alu1 92 36 92 36 6 a1
<< end >>
