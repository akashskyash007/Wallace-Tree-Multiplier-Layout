magic
tech scmos
timestamp 1199540192
<< ab >>
rect -12 0 314 100
<< alu1 >>
rect -10 81 -6 92
rect -10 79 -9 81
rect -7 79 -6 81
rect -10 61 -6 79
rect -10 59 -9 61
rect -7 59 -6 61
rect -10 41 -6 59
rect -10 39 -9 41
rect -7 39 -6 41
rect -10 21 -6 39
rect -10 19 -9 21
rect -7 19 -6 21
rect -10 12 -6 19
rect -10 8 314 12
<< alu2 >>
rect -12 81 314 82
rect -12 79 -9 81
rect -7 79 314 81
rect -12 78 314 79
rect -12 61 314 62
rect -12 59 -9 61
rect -7 59 314 61
rect -12 58 314 59
rect -12 41 314 42
rect -12 39 -9 41
rect -7 39 314 41
rect -12 38 314 39
rect -12 21 314 22
rect -12 19 -9 21
rect -7 19 9 21
rect 11 19 29 21
rect 31 19 49 21
rect 51 19 69 21
rect 71 19 89 21
rect 91 19 109 21
rect 111 19 129 21
rect 131 19 149 21
rect 151 19 169 21
rect 171 19 189 21
rect 191 19 209 21
rect 211 19 229 21
rect 231 19 249 21
rect 251 19 269 21
rect 271 19 289 21
rect 291 19 309 21
rect 311 19 314 21
rect -12 18 314 19
<< alu3 >>
rect 8 91 12 94
rect 8 89 9 91
rect 11 89 12 91
rect 8 71 12 89
rect 8 69 9 71
rect 11 69 12 71
rect 8 51 12 69
rect 8 49 9 51
rect 11 49 12 51
rect 8 31 12 49
rect 8 29 9 31
rect 11 29 12 31
rect 8 21 12 29
rect 8 19 9 21
rect 11 19 12 21
rect 8 11 12 19
rect 8 9 9 11
rect 11 9 12 11
rect 8 6 12 9
rect 28 21 32 92
rect 28 19 29 21
rect 31 19 32 21
rect 28 8 32 19
rect 48 21 52 92
rect 48 19 49 21
rect 51 19 52 21
rect 48 8 52 19
rect 68 21 72 92
rect 68 19 69 21
rect 71 19 72 21
rect 68 8 72 19
rect 88 21 92 92
rect 88 19 89 21
rect 91 19 92 21
rect 88 8 92 19
rect 108 21 112 92
rect 108 19 109 21
rect 111 19 112 21
rect 108 8 112 19
rect 128 21 132 92
rect 128 19 129 21
rect 131 19 132 21
rect 128 8 132 19
rect 148 21 152 92
rect 148 19 149 21
rect 151 19 152 21
rect 148 8 152 19
rect 168 21 172 92
rect 168 19 169 21
rect 171 19 172 21
rect 168 8 172 19
rect 188 21 192 92
rect 188 19 189 21
rect 191 19 192 21
rect 188 8 192 19
rect 208 21 212 92
rect 208 19 209 21
rect 211 19 212 21
rect 208 8 212 19
rect 228 21 232 92
rect 228 19 229 21
rect 231 19 232 21
rect 228 8 232 19
rect 248 21 252 92
rect 248 19 249 21
rect 251 19 252 21
rect 248 8 252 19
rect 268 21 272 92
rect 268 19 269 21
rect 271 19 272 21
rect 268 8 272 19
rect 288 21 292 92
rect 288 19 289 21
rect 291 19 292 21
rect 288 8 292 19
rect 308 21 312 92
rect 308 19 309 21
rect 311 19 312 21
rect 308 8 312 19
<< alu4 >>
rect -10 91 314 92
rect -10 89 9 91
rect 11 89 314 91
rect -10 88 314 89
rect -10 71 314 72
rect -10 69 9 71
rect 11 69 314 71
rect -10 68 314 69
rect -10 51 314 52
rect -10 49 9 51
rect 11 49 314 51
rect -10 48 314 49
rect -10 31 314 32
rect -10 29 -1 31
rect 1 29 9 31
rect 11 29 19 31
rect 21 29 39 31
rect 41 29 59 31
rect 61 29 79 31
rect 81 29 99 31
rect 101 29 119 31
rect 121 29 139 31
rect 141 29 159 31
rect 161 29 179 31
rect 181 29 199 31
rect 201 29 219 31
rect 221 29 239 31
rect 241 29 259 31
rect 261 29 279 31
rect 281 29 299 31
rect 301 29 314 31
rect -10 28 314 29
rect -10 11 314 12
rect -10 9 9 11
rect 11 9 314 11
rect -10 8 314 9
<< alu5 >>
rect -2 31 2 92
rect -2 29 -1 31
rect 1 29 2 31
rect -2 8 2 29
rect 18 31 22 92
rect 18 29 19 31
rect 21 29 22 31
rect 18 8 22 29
rect 38 31 42 92
rect 38 29 39 31
rect 41 29 42 31
rect 38 8 42 29
rect 58 31 62 92
rect 58 29 59 31
rect 61 29 62 31
rect 58 8 62 29
rect 78 31 82 92
rect 78 29 79 31
rect 81 29 82 31
rect 78 8 82 29
rect 98 31 102 92
rect 98 29 99 31
rect 101 29 102 31
rect 98 8 102 29
rect 118 31 122 92
rect 118 29 119 31
rect 121 29 122 31
rect 118 8 122 29
rect 138 31 142 92
rect 138 29 139 31
rect 141 29 142 31
rect 138 8 142 29
rect 158 31 162 92
rect 158 29 159 31
rect 161 29 162 31
rect 158 8 162 29
rect 178 31 182 92
rect 178 29 179 31
rect 181 29 182 31
rect 178 8 182 29
rect 198 31 202 92
rect 198 29 199 31
rect 201 29 202 31
rect 198 8 202 29
rect 218 31 222 92
rect 218 29 219 31
rect 221 29 222 31
rect 218 8 222 29
rect 238 31 242 92
rect 238 29 239 31
rect 241 29 242 31
rect 238 8 242 29
rect 258 31 262 92
rect 258 29 259 31
rect 261 29 262 31
rect 258 8 262 29
rect 278 31 282 92
rect 278 29 279 31
rect 281 29 282 31
rect 278 8 282 29
rect 298 31 302 92
rect 298 29 299 31
rect 301 29 302 31
rect 298 8 302 29
<< via1 >>
rect -9 79 -7 81
rect -9 59 -7 61
rect -9 39 -7 41
rect -9 19 -7 21
<< via2 >>
rect 9 19 11 21
rect 29 19 31 21
rect 49 19 51 21
rect 69 19 71 21
rect 89 19 91 21
rect 109 19 111 21
rect 129 19 131 21
rect 149 19 151 21
rect 169 19 171 21
rect 189 19 191 21
rect 209 19 211 21
rect 229 19 231 21
rect 249 19 251 21
rect 269 19 271 21
rect 289 19 291 21
rect 309 19 311 21
<< via3 >>
rect 9 89 11 91
rect 9 69 11 71
rect 9 49 11 51
rect 9 29 11 31
rect 9 9 11 11
<< via4 >>
rect -1 29 1 31
rect 19 29 21 31
rect 39 29 41 31
rect 59 29 61 31
rect 79 29 81 31
rect 99 29 101 31
rect 119 29 121 31
rect 139 29 141 31
rect 159 29 161 31
rect 179 29 181 31
rect 199 29 201 31
rect 219 29 221 31
rect 239 29 241 31
rect 259 29 261 31
rect 279 29 281 31
rect 299 29 301 31
<< end >>
