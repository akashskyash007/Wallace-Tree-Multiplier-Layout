magic
tech scmos
timestamp 1199470294
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 45 83 47 88
rect 53 83 55 88
rect 21 77 23 82
rect 33 71 35 76
rect 21 42 23 57
rect 33 52 35 57
rect 33 50 41 52
rect 33 48 37 50
rect 39 48 41 50
rect 33 46 41 48
rect 21 40 31 42
rect 21 38 27 40
rect 29 38 31 40
rect 11 36 31 38
rect 11 33 13 36
rect 35 29 37 46
rect 45 43 47 57
rect 53 52 55 57
rect 53 50 63 52
rect 57 48 59 50
rect 61 48 63 50
rect 57 46 63 48
rect 45 41 53 43
rect 45 39 49 41
rect 51 39 53 41
rect 45 37 53 39
rect 47 29 49 37
rect 57 29 59 46
rect 11 18 13 23
rect 35 12 37 17
rect 47 12 49 17
rect 57 12 59 17
<< ndif >>
rect 3 31 11 33
rect 3 29 5 31
rect 7 29 11 31
rect 3 23 11 29
rect 13 31 21 33
rect 13 29 17 31
rect 19 29 21 31
rect 13 27 21 29
rect 27 27 35 29
rect 13 23 18 27
rect 27 25 29 27
rect 31 25 35 27
rect 27 23 35 25
rect 30 17 35 23
rect 37 21 47 29
rect 37 19 41 21
rect 43 19 47 21
rect 37 17 47 19
rect 49 17 57 29
rect 59 23 64 29
rect 59 21 67 23
rect 59 19 63 21
rect 65 19 67 21
rect 59 17 67 19
rect 51 10 55 17
rect 51 8 57 10
rect 51 6 53 8
rect 55 6 57 8
rect 51 4 57 6
<< pdif >>
rect 16 71 21 77
rect 13 69 21 71
rect 13 67 15 69
rect 17 67 21 69
rect 13 61 21 67
rect 13 59 15 61
rect 17 59 21 61
rect 13 57 21 59
rect 23 71 31 77
rect 40 71 45 83
rect 23 69 27 71
rect 29 69 33 71
rect 23 57 33 69
rect 35 69 45 71
rect 35 67 39 69
rect 41 67 45 69
rect 35 61 45 67
rect 35 59 39 61
rect 41 59 45 61
rect 35 57 45 59
rect 47 57 53 83
rect 55 81 63 83
rect 55 79 59 81
rect 61 79 63 81
rect 55 57 63 79
<< alu1 >>
rect -2 95 72 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 72 95
rect -2 88 72 93
rect 26 71 30 88
rect 58 81 62 88
rect 58 79 59 81
rect 61 79 62 81
rect 58 77 62 79
rect 14 69 18 71
rect 14 67 15 69
rect 17 67 18 69
rect 26 69 27 71
rect 29 69 30 71
rect 26 67 30 69
rect 38 69 42 71
rect 38 67 39 69
rect 41 67 42 69
rect 47 68 62 73
rect 14 63 18 67
rect 8 61 22 63
rect 38 61 42 67
rect 8 59 15 61
rect 17 59 22 61
rect 8 57 22 59
rect 18 36 22 57
rect 28 59 39 61
rect 41 59 42 61
rect 28 57 42 59
rect 28 42 32 57
rect 36 50 42 53
rect 36 48 37 50
rect 39 48 42 50
rect 36 46 42 48
rect 26 40 32 42
rect 26 38 27 40
rect 29 38 32 40
rect 26 36 32 38
rect 4 31 8 33
rect 4 29 5 31
rect 7 29 8 31
rect 4 12 8 29
rect 16 31 22 36
rect 16 29 17 31
rect 19 29 22 31
rect 16 27 22 29
rect 28 27 32 36
rect 38 32 42 46
rect 48 42 52 63
rect 58 50 62 68
rect 58 48 59 50
rect 61 48 62 50
rect 58 46 62 48
rect 48 41 63 42
rect 48 39 49 41
rect 51 39 63 41
rect 48 37 63 39
rect 38 27 53 32
rect 28 25 29 27
rect 31 25 32 27
rect 28 23 32 25
rect 39 21 67 22
rect 39 19 41 21
rect 43 19 63 21
rect 65 19 67 21
rect 39 18 67 19
rect -2 8 72 12
rect -2 7 53 8
rect -2 5 9 7
rect 11 5 19 7
rect 21 6 53 7
rect 55 6 72 8
rect 21 5 72 6
rect -2 0 72 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 11 23 13 33
rect 35 17 37 29
rect 47 17 49 29
rect 57 17 59 29
<< pmos >>
rect 21 57 23 77
rect 33 57 35 71
rect 45 57 47 83
rect 53 57 55 83
<< polyct1 >>
rect 37 48 39 50
rect 27 38 29 40
rect 59 48 61 50
rect 49 39 51 41
<< ndifct1 >>
rect 5 29 7 31
rect 17 29 19 31
rect 29 25 31 27
rect 41 19 43 21
rect 63 19 65 21
rect 53 6 55 8
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 15 67 17 69
rect 15 59 17 61
rect 27 69 29 71
rect 39 67 41 69
rect 39 59 41 61
rect 59 79 61 81
<< labels >>
rlabel ndifct1 42 20 42 20 6 n2
rlabel ndifct1 30 26 30 26 6 zn
rlabel polyct1 28 39 28 39 6 zn
rlabel pdifct1 40 60 40 60 6 zn
rlabel pdifct1 40 68 40 68 6 zn
rlabel ndifct1 64 20 64 20 6 n2
rlabel alu1 10 60 10 60 6 z
rlabel alu1 20 45 20 45 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 40 40 40 6 b
rlabel alu1 50 30 50 30 6 b
rlabel alu1 50 50 50 50 6 a2
rlabel alu1 50 70 50 70 6 a1
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 40 60 40 6 a2
rlabel alu1 60 60 60 60 6 a1
<< end >>
