magic
tech scmos
timestamp 1199203066
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 30 68 32 73
rect 37 68 39 73
rect 10 61 12 65
rect 20 61 22 65
rect 10 47 12 52
rect 9 45 15 47
rect 9 43 11 45
rect 13 43 15 45
rect 9 41 15 43
rect 9 23 11 41
rect 20 32 22 52
rect 30 38 32 52
rect 37 49 39 52
rect 37 47 46 49
rect 37 45 42 47
rect 44 45 46 47
rect 37 43 46 45
rect 16 30 22 32
rect 16 28 18 30
rect 20 28 22 30
rect 16 26 22 28
rect 26 36 33 38
rect 26 34 29 36
rect 31 34 33 36
rect 26 32 33 34
rect 16 23 18 26
rect 26 23 28 32
rect 37 29 39 43
rect 37 15 39 19
rect 9 8 11 13
rect 16 8 18 13
rect 26 8 28 13
<< ndif >>
rect 30 23 37 29
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 13 9 17
rect 11 13 16 23
rect 18 20 26 23
rect 18 18 21 20
rect 23 18 26 20
rect 18 13 26 18
rect 28 19 37 23
rect 39 25 44 29
rect 39 23 46 25
rect 39 21 42 23
rect 44 21 46 23
rect 39 19 46 21
rect 28 13 35 19
rect 30 11 36 13
rect 30 9 32 11
rect 34 9 36 11
rect 30 7 36 9
<< pdif >>
rect 2 71 8 73
rect 2 69 4 71
rect 6 69 8 71
rect 2 61 8 69
rect 22 71 28 73
rect 22 69 24 71
rect 26 69 28 71
rect 22 68 28 69
rect 22 67 30 68
rect 24 61 30 67
rect 2 52 10 61
rect 12 59 20 61
rect 12 57 15 59
rect 17 57 20 59
rect 12 52 20 57
rect 22 52 30 61
rect 32 52 37 68
rect 39 64 44 68
rect 39 62 46 64
rect 39 60 42 62
rect 44 60 46 62
rect 39 58 46 60
rect 39 52 44 58
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 71 50 79
rect -2 69 4 71
rect 6 69 24 71
rect 26 69 50 71
rect -2 68 50 69
rect 2 62 46 63
rect 2 60 42 62
rect 44 60 46 62
rect 2 59 46 60
rect 2 57 15 59
rect 17 57 22 59
rect 2 21 6 57
rect 26 47 30 55
rect 34 49 46 55
rect 10 45 30 47
rect 10 43 11 45
rect 13 43 30 45
rect 42 47 46 49
rect 44 45 46 47
rect 10 41 22 43
rect 42 41 46 45
rect 26 36 38 39
rect 26 34 29 36
rect 31 34 38 36
rect 26 33 38 34
rect 10 30 22 31
rect 10 28 18 30
rect 20 28 22 30
rect 10 25 22 28
rect 34 25 38 33
rect 2 19 4 21
rect 2 17 6 19
rect 10 17 14 25
rect -2 11 50 12
rect -2 9 32 11
rect 34 9 50 11
rect -2 1 50 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 9 13 11 23
rect 16 13 18 23
rect 26 13 28 23
rect 37 19 39 29
<< pmos >>
rect 10 52 12 61
rect 20 52 22 61
rect 30 52 32 68
rect 37 52 39 68
<< polyct1 >>
rect 11 43 13 45
rect 42 45 44 47
rect 18 28 20 30
rect 29 34 31 36
<< ndifct0 >>
rect 21 18 23 20
rect 42 21 44 23
<< ndifct1 >>
rect 4 19 6 21
rect 32 9 34 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct1 >>
rect 4 69 6 71
rect 24 69 26 71
rect 15 57 17 59
rect 42 60 44 62
<< alu0 >>
rect 13 56 19 57
rect 41 43 42 49
rect 6 17 7 23
rect 41 23 45 25
rect 41 21 42 23
rect 44 21 45 23
rect 19 20 45 21
rect 19 18 21 20
rect 23 18 45 20
rect 19 17 45 18
<< labels >>
rlabel alu0 32 19 32 19 6 n1
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 24 12 24 6 b
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 44 20 44 6 c
rlabel polyct1 12 44 12 44 6 c
rlabel alu1 20 60 20 60 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 36 28 36 6 a1
rlabel alu1 28 52 28 52 6 c
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 36 32 36 32 6 a1
rlabel alu1 36 52 36 52 6 a2
rlabel alu1 44 48 44 48 6 a2
<< end >>
