magic
tech scmos
timestamp 1199201807
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 12 66 14 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 12 28 14 39
rect 19 36 21 39
rect 29 36 31 39
rect 39 36 41 39
rect 19 34 25 36
rect 19 32 21 34
rect 23 32 25 34
rect 19 30 25 32
rect 29 34 35 36
rect 29 32 31 34
rect 33 32 35 34
rect 29 30 35 32
rect 39 34 47 36
rect 39 32 43 34
rect 45 32 47 34
rect 39 30 47 32
rect 9 26 15 28
rect 9 24 11 26
rect 13 24 15 26
rect 9 22 15 24
rect 10 19 12 22
rect 20 19 22 30
rect 32 22 34 30
rect 39 22 41 30
rect 10 8 12 13
rect 20 8 22 13
rect 32 8 34 13
rect 39 8 41 13
<< ndif >>
rect 24 19 32 22
rect 2 13 10 19
rect 12 17 20 19
rect 12 15 15 17
rect 17 15 20 17
rect 12 13 20 15
rect 22 13 32 19
rect 34 13 39 22
rect 41 19 46 22
rect 41 17 48 19
rect 41 15 44 17
rect 46 15 48 17
rect 41 13 48 15
rect 2 7 8 13
rect 2 5 4 7
rect 6 5 8 7
rect 2 3 8 5
rect 24 7 30 13
rect 24 5 26 7
rect 28 5 30 7
rect 24 3 30 5
<< pdif >>
rect 7 60 12 66
rect 5 58 12 60
rect 5 56 7 58
rect 9 56 12 58
rect 5 50 12 56
rect 5 48 7 50
rect 9 48 12 50
rect 5 46 12 48
rect 7 39 12 46
rect 14 39 19 66
rect 21 57 29 66
rect 21 55 24 57
rect 26 55 29 57
rect 21 39 29 55
rect 31 64 39 66
rect 31 62 34 64
rect 36 62 39 64
rect 31 39 39 62
rect 41 59 46 66
rect 41 57 48 59
rect 41 55 44 57
rect 46 55 48 57
rect 41 53 48 55
rect 41 39 46 53
<< alu1 >>
rect -2 64 58 72
rect 2 58 11 59
rect 2 56 7 58
rect 9 56 11 58
rect 2 55 11 56
rect 2 18 6 55
rect 18 45 30 51
rect 34 45 46 51
rect 10 26 14 43
rect 18 37 24 45
rect 20 34 24 37
rect 20 32 21 34
rect 23 32 24 34
rect 20 30 24 32
rect 29 34 38 35
rect 29 32 31 34
rect 33 32 38 34
rect 29 31 38 32
rect 33 26 38 31
rect 42 34 46 45
rect 42 32 43 34
rect 45 32 46 34
rect 42 30 46 32
rect 10 24 11 26
rect 13 24 23 26
rect 10 22 23 24
rect 33 22 47 26
rect 2 17 48 18
rect 2 15 15 17
rect 17 15 44 17
rect 46 15 48 17
rect 2 14 48 15
rect -2 7 58 8
rect -2 5 4 7
rect 6 5 26 7
rect 28 5 49 7
rect 51 5 58 7
rect -2 0 58 5
<< ptie >>
rect 47 7 53 9
rect 47 5 49 7
rect 51 5 53 7
rect 47 3 53 5
<< nmos >>
rect 10 13 12 19
rect 20 13 22 19
rect 32 13 34 22
rect 39 13 41 22
<< pmos >>
rect 12 39 14 66
rect 19 39 21 66
rect 29 39 31 66
rect 39 39 41 66
<< polyct1 >>
rect 21 32 23 34
rect 31 32 33 34
rect 43 32 45 34
rect 11 24 13 26
<< ndifct1 >>
rect 15 15 17 17
rect 44 15 46 17
rect 4 5 6 7
rect 26 5 28 7
<< ptiect1 >>
rect 49 5 51 7
<< pdifct0 >>
rect 7 48 9 50
rect 24 55 26 57
rect 34 62 36 64
rect 44 55 46 57
<< pdifct1 >>
rect 7 56 9 58
<< alu0 >>
rect 32 62 34 64
rect 36 62 38 64
rect 32 61 38 62
rect 22 57 48 58
rect 22 55 24 57
rect 26 55 44 57
rect 46 55 48 57
rect 22 54 48 55
rect 6 50 11 51
rect 6 48 7 50
rect 9 48 11 50
rect 6 47 11 48
<< labels >>
rlabel alu0 35 56 35 56 6 n1
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 24 20 24 6 c
rlabel alu1 12 36 12 36 6 c
rlabel alu1 20 44 20 44 6 b
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 16 36 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 28 48 28 48 6 b
rlabel alu1 36 48 36 48 6 a2
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 16 44 16 6 z
rlabel alu1 44 24 44 24 6 a1
rlabel alu1 44 44 44 44 6 a2
<< end >>
