magic
tech scmos
timestamp 1199202296
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 58 41 62
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 33 41 35
rect 9 26 11 33
rect 19 26 21 33
rect 27 31 29 33
rect 31 31 37 33
rect 39 31 41 33
rect 27 29 41 31
rect 29 26 31 29
rect 39 26 41 29
rect 9 12 11 17
rect 19 2 21 6
rect 29 2 31 6
rect 39 2 41 6
<< ndif >>
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 14 6 19 17
rect 21 17 29 26
rect 21 15 24 17
rect 26 15 29 17
rect 21 10 29 15
rect 21 8 24 10
rect 26 8 29 10
rect 21 6 29 8
rect 31 24 39 26
rect 31 22 34 24
rect 36 22 39 24
rect 31 17 39 22
rect 31 15 34 17
rect 36 15 39 17
rect 31 6 39 15
rect 41 17 49 26
rect 41 15 45 17
rect 47 15 49 17
rect 41 10 49 15
rect 41 8 45 10
rect 47 8 49 10
rect 41 6 49 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 56 29 62
rect 21 54 24 56
rect 26 54 29 56
rect 21 38 29 54
rect 31 58 36 66
rect 31 49 39 58
rect 31 47 34 49
rect 36 47 39 49
rect 31 42 39 47
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 56 48 58
rect 41 54 44 56
rect 46 54 48 56
rect 41 49 48 54
rect 41 47 44 49
rect 46 47 48 49
rect 41 38 48 47
<< alu1 >>
rect -2 67 58 72
rect -2 65 49 67
rect 51 65 58 67
rect -2 64 58 65
rect 10 40 14 43
rect 33 49 38 51
rect 33 47 34 49
rect 36 47 38 49
rect 33 42 38 47
rect 16 40 34 42
rect 36 40 38 42
rect 10 38 38 40
rect 10 26 14 38
rect 42 34 46 43
rect 25 33 46 34
rect 25 31 29 33
rect 31 31 37 33
rect 39 31 46 33
rect 25 30 46 31
rect 10 24 39 26
rect 10 22 14 24
rect 16 22 34 24
rect 36 22 39 24
rect 10 21 18 22
rect 33 17 39 22
rect 33 15 34 17
rect 36 15 39 17
rect 33 13 39 15
rect -2 7 58 8
rect -2 5 5 7
rect 7 5 58 7
rect -2 0 58 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 47 67 53 69
rect 47 65 49 67
rect 51 65 53 67
rect 47 63 53 65
<< nmos >>
rect 9 17 11 26
rect 19 6 21 26
rect 29 6 31 26
rect 39 6 41 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 58
<< polyct1 >>
rect 29 31 31 33
rect 37 31 39 33
<< ndifct0 >>
rect 4 19 6 21
rect 24 15 26 17
rect 24 8 26 10
rect 45 15 47 17
rect 45 8 47 10
<< ndifct1 >>
rect 14 22 16 24
rect 34 22 36 24
rect 34 15 36 17
<< ntiect1 >>
rect 49 65 51 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 47 16 49
rect 24 62 26 64
rect 24 54 26 56
rect 44 54 46 56
rect 44 47 46 49
<< pdifct1 >>
rect 14 40 16 42
rect 34 47 36 49
rect 34 40 36 42
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 23 62 24 64
rect 26 62 27 64
rect 23 56 27 62
rect 23 54 24 56
rect 26 54 27 56
rect 23 52 27 54
rect 42 56 48 64
rect 42 54 44 56
rect 46 54 48 56
rect 13 49 17 51
rect 13 47 14 49
rect 16 47 17 49
rect 13 43 17 47
rect 14 42 17 43
rect 42 49 48 54
rect 42 47 44 49
rect 46 47 48 49
rect 42 46 48 47
rect 3 21 7 23
rect 3 19 4 21
rect 6 19 7 21
rect 3 8 7 19
rect 22 17 28 18
rect 22 15 24 17
rect 26 15 28 17
rect 22 10 28 15
rect 43 17 49 18
rect 43 15 45 17
rect 47 15 49 17
rect 22 8 24 10
rect 26 8 28 10
rect 43 10 49 15
rect 43 8 45 10
rect 47 8 49 10
<< labels >>
rlabel alu1 12 32 12 32 6 z
rlabel alu1 20 24 20 24 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 28 32 28 32 6 a
rlabel alu1 36 32 36 32 6 a
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 40 44 40 6 a
<< end >>
