magic
tech scmos
timestamp 1199202438
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 42 68 71 70
rect 9 56 11 61
rect 35 60 37 65
rect 42 60 44 68
rect 52 60 54 64
rect 59 60 61 64
rect 69 60 71 68
rect 19 50 21 55
rect 35 51 37 54
rect 31 49 37 51
rect 31 47 33 49
rect 35 47 37 49
rect 31 45 37 47
rect 9 35 11 38
rect 19 35 21 38
rect 9 33 31 35
rect 10 16 12 33
rect 24 31 27 33
rect 29 31 31 33
rect 24 29 31 31
rect 24 26 26 29
rect 35 20 37 45
rect 42 35 44 54
rect 52 45 54 48
rect 48 43 54 45
rect 59 43 61 48
rect 48 41 50 43
rect 52 41 54 43
rect 48 39 54 41
rect 58 41 64 43
rect 58 39 60 41
rect 62 39 64 41
rect 58 37 64 39
rect 42 33 54 35
rect 41 27 47 29
rect 41 25 43 27
rect 45 25 47 27
rect 41 23 47 25
rect 42 20 44 23
rect 52 20 54 33
rect 59 20 61 37
rect 69 33 71 48
rect 65 31 71 33
rect 65 29 67 31
rect 69 29 71 31
rect 65 27 71 29
rect 69 24 71 27
rect 24 15 26 20
rect 35 9 37 14
rect 42 9 44 14
rect 52 9 54 14
rect 59 9 61 14
rect 69 13 71 18
rect 10 2 12 7
<< ndif >>
rect 2 16 8 18
rect 17 24 24 26
rect 17 22 19 24
rect 21 22 24 24
rect 17 20 24 22
rect 26 24 33 26
rect 26 22 29 24
rect 31 22 33 24
rect 26 20 33 22
rect 63 20 69 24
rect 2 14 4 16
rect 6 14 10 16
rect 2 12 10 14
rect 5 7 10 12
rect 12 11 19 16
rect 28 14 35 20
rect 37 14 42 20
rect 44 18 52 20
rect 44 16 47 18
rect 49 16 52 18
rect 44 14 52 16
rect 54 14 59 20
rect 61 18 69 20
rect 71 22 78 24
rect 71 20 74 22
rect 76 20 78 22
rect 71 18 78 20
rect 61 14 67 18
rect 12 9 15 11
rect 17 9 19 11
rect 63 11 67 14
rect 12 7 19 9
rect 63 7 69 11
rect 63 5 65 7
rect 67 5 69 7
rect 63 3 69 5
<< pdif >>
rect 28 58 35 60
rect 28 56 30 58
rect 32 56 35 58
rect 4 51 9 56
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 50 17 56
rect 28 54 35 56
rect 37 54 42 60
rect 44 58 52 60
rect 44 56 47 58
rect 49 56 52 58
rect 44 54 52 56
rect 11 48 19 50
rect 11 46 14 48
rect 16 46 19 48
rect 11 38 19 46
rect 21 48 28 50
rect 21 46 24 48
rect 26 46 28 48
rect 21 44 28 46
rect 21 38 26 44
rect 47 48 52 54
rect 54 48 59 60
rect 61 58 69 60
rect 61 56 64 58
rect 66 56 69 58
rect 61 48 69 56
rect 71 54 76 60
rect 71 52 78 54
rect 71 50 74 52
rect 76 50 78 52
rect 71 48 78 50
<< alu1 >>
rect -2 67 82 72
rect -2 65 5 67
rect 7 65 13 67
rect 15 65 82 67
rect -2 64 82 65
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 2 40 4 42
rect 6 40 7 42
rect 2 38 7 40
rect 2 27 6 38
rect 2 21 14 27
rect 2 16 8 21
rect 2 14 4 16
rect 6 14 8 16
rect 2 13 8 14
rect 58 41 63 43
rect 58 39 60 41
rect 62 39 63 41
rect 58 37 63 39
rect 58 26 62 37
rect 49 22 62 26
rect 66 31 70 33
rect 66 29 67 31
rect 69 29 70 31
rect 66 18 70 29
rect 57 14 70 18
rect -2 7 82 8
rect -2 5 25 7
rect 27 5 65 7
rect 67 5 82 7
rect -2 0 82 5
<< ptie >>
rect 23 7 29 9
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< ntie >>
rect 3 67 17 69
rect 3 65 5 67
rect 7 65 13 67
rect 15 65 17 67
rect 3 63 17 65
<< nmos >>
rect 24 20 26 26
rect 10 7 12 16
rect 35 14 37 20
rect 42 14 44 20
rect 52 14 54 20
rect 59 14 61 20
rect 69 18 71 24
<< pmos >>
rect 9 38 11 56
rect 35 54 37 60
rect 42 54 44 60
rect 19 38 21 50
rect 52 48 54 60
rect 59 48 61 60
rect 69 48 71 60
<< polyct0 >>
rect 33 47 35 49
rect 27 31 29 33
rect 50 41 52 43
rect 43 25 45 27
<< polyct1 >>
rect 60 39 62 41
rect 67 29 69 31
<< ndifct0 >>
rect 19 22 21 24
rect 29 22 31 24
rect 47 16 49 18
rect 74 20 76 22
rect 15 9 17 11
<< ndifct1 >>
rect 4 14 6 16
rect 65 5 67 7
<< ntiect1 >>
rect 5 65 7 67
rect 13 65 15 67
<< ptiect1 >>
rect 25 5 27 7
<< pdifct0 >>
rect 30 56 32 58
rect 47 56 49 58
rect 14 46 16 48
rect 24 46 26 48
rect 64 56 66 58
rect 74 50 76 52
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
<< alu0 >>
rect 12 48 18 64
rect 29 58 33 64
rect 29 56 30 58
rect 32 56 33 58
rect 29 54 33 56
rect 41 58 51 59
rect 41 56 47 58
rect 49 56 51 58
rect 41 55 51 56
rect 63 58 67 64
rect 63 56 64 58
rect 66 56 67 58
rect 12 46 14 48
rect 16 46 18 48
rect 12 45 18 46
rect 23 49 37 50
rect 23 48 33 49
rect 23 46 24 48
rect 26 47 33 48
rect 35 47 37 49
rect 26 46 37 47
rect 23 42 27 46
rect 41 42 45 55
rect 63 54 67 56
rect 73 52 77 54
rect 73 50 74 52
rect 76 50 77 52
rect 18 38 27 42
rect 35 38 45 42
rect 49 46 78 50
rect 49 43 53 46
rect 49 41 50 43
rect 52 41 53 43
rect 18 24 22 38
rect 35 34 39 38
rect 49 34 53 41
rect 25 33 39 34
rect 25 31 27 33
rect 29 31 39 33
rect 25 30 39 31
rect 18 22 19 24
rect 21 22 22 24
rect 18 20 22 22
rect 28 24 32 26
rect 28 22 29 24
rect 31 22 32 24
rect 14 11 18 13
rect 14 9 15 11
rect 17 9 18 11
rect 14 8 18 9
rect 28 8 32 22
rect 35 19 39 30
rect 42 30 53 34
rect 42 27 46 30
rect 42 25 43 27
rect 45 25 46 27
rect 42 23 46 25
rect 35 18 51 19
rect 74 24 78 46
rect 73 22 78 24
rect 73 20 74 22
rect 76 20 78 22
rect 73 18 78 20
rect 35 16 47 18
rect 49 16 51 18
rect 35 15 51 16
<< labels >>
rlabel alu0 32 32 32 32 6 n1
rlabel alu0 25 44 25 44 6 n2
rlabel alu0 20 31 20 31 6 n2
rlabel alu0 30 48 30 48 6 n2
rlabel alu0 43 17 43 17 6 n1
rlabel alu0 44 28 44 28 6 en
rlabel alu0 51 40 51 40 6 en
rlabel alu0 46 57 46 57 6 n1
rlabel alu0 76 34 76 34 6 en
rlabel alu0 75 50 75 50 6 en
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 52 24 52 24 6 d
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 60 16 60 16 6 e
rlabel alu1 68 24 68 24 6 e
rlabel alu1 60 36 60 36 6 d
<< end >>
