magic
tech scmos
timestamp 1199469175
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -5 48 95 105
<< pwell >>
rect -5 -5 95 48
<< poly >>
rect 11 93 13 98
rect 41 93 43 98
rect 53 93 55 98
rect 65 93 67 98
rect 77 93 79 98
rect 11 52 13 55
rect 11 50 32 52
rect 25 48 28 50
rect 30 48 32 50
rect 25 46 32 48
rect 25 36 27 46
rect 41 43 43 55
rect 53 52 55 55
rect 65 52 67 55
rect 53 49 57 52
rect 65 50 73 52
rect 65 49 69 50
rect 55 43 57 49
rect 67 48 69 49
rect 71 48 73 50
rect 67 46 73 48
rect 41 41 51 43
rect 45 39 47 41
rect 49 39 51 41
rect 45 37 51 39
rect 55 41 63 43
rect 55 39 59 41
rect 61 39 63 41
rect 55 37 63 39
rect 47 34 49 37
rect 55 34 57 37
rect 67 34 69 46
rect 77 43 79 55
rect 77 41 83 43
rect 77 40 79 41
rect 75 39 79 40
rect 81 39 83 41
rect 75 37 83 39
rect 75 34 77 37
rect 25 12 27 17
rect 47 12 49 17
rect 55 12 57 17
rect 67 12 69 17
rect 75 12 77 17
<< ndif >>
rect 17 34 25 36
rect 17 32 19 34
rect 21 32 25 34
rect 17 26 25 32
rect 17 24 19 26
rect 21 24 25 26
rect 17 22 25 24
rect 20 17 25 22
rect 27 34 41 36
rect 27 31 47 34
rect 27 29 31 31
rect 33 29 47 31
rect 27 21 47 29
rect 27 19 31 21
rect 33 19 47 21
rect 27 17 47 19
rect 49 17 55 34
rect 57 21 67 34
rect 57 19 61 21
rect 63 19 67 21
rect 57 17 67 19
rect 69 17 75 34
rect 77 21 86 34
rect 77 19 81 21
rect 83 19 86 21
rect 77 17 86 19
<< pdif >>
rect 3 91 11 93
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 55 11 69
rect 13 71 18 93
rect 36 83 41 93
rect 33 81 41 83
rect 33 79 35 81
rect 37 79 41 81
rect 33 77 41 79
rect 13 69 21 71
rect 13 67 17 69
rect 19 67 21 69
rect 13 61 21 67
rect 13 59 17 61
rect 19 59 21 61
rect 13 57 21 59
rect 13 55 18 57
rect 36 55 41 77
rect 43 71 53 93
rect 43 69 47 71
rect 49 69 53 71
rect 43 55 53 69
rect 55 81 65 93
rect 55 79 59 81
rect 61 79 65 81
rect 55 55 65 79
rect 67 91 77 93
rect 67 89 71 91
rect 73 89 77 91
rect 67 55 77 89
rect 79 82 84 93
rect 79 80 87 82
rect 79 78 83 80
rect 85 78 87 80
rect 79 72 87 78
rect 79 70 83 72
rect 85 70 87 72
rect 79 68 87 70
rect 79 55 84 68
<< alu1 >>
rect -2 95 92 100
rect -2 93 26 95
rect 28 93 92 95
rect -2 91 92 93
rect -2 89 5 91
rect 7 89 71 91
rect 73 89 92 91
rect -2 88 92 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 71 8 79
rect 33 81 86 82
rect 33 79 35 81
rect 37 79 59 81
rect 61 80 86 81
rect 61 79 83 80
rect 33 78 83 79
rect 85 78 86 80
rect 4 69 5 71
rect 7 69 8 71
rect 4 67 8 69
rect 16 69 22 73
rect 16 67 17 69
rect 19 67 22 69
rect 16 62 22 67
rect 7 61 22 62
rect 7 59 17 61
rect 19 59 22 61
rect 7 58 22 59
rect 18 34 22 58
rect 38 71 51 72
rect 38 69 47 71
rect 49 69 51 71
rect 38 68 51 69
rect 38 51 42 68
rect 58 62 62 73
rect 47 58 62 62
rect 26 50 42 51
rect 26 48 28 50
rect 30 48 42 50
rect 26 47 42 48
rect 18 32 19 34
rect 21 32 22 34
rect 18 26 22 32
rect 18 24 19 26
rect 21 24 22 26
rect 18 17 22 24
rect 30 31 34 33
rect 30 29 31 31
rect 33 29 34 31
rect 30 21 34 29
rect 30 19 31 21
rect 33 19 34 21
rect 30 12 34 19
rect 38 22 42 47
rect 48 43 52 53
rect 46 41 52 43
rect 46 39 47 41
rect 49 39 52 41
rect 46 37 52 39
rect 58 41 62 58
rect 58 39 59 41
rect 61 39 62 41
rect 58 37 62 39
rect 68 62 72 73
rect 82 72 86 78
rect 82 70 83 72
rect 85 70 86 72
rect 82 68 86 70
rect 68 58 83 62
rect 68 50 72 58
rect 68 48 69 50
rect 71 48 72 50
rect 68 37 72 48
rect 78 41 82 53
rect 78 39 79 41
rect 81 39 82 41
rect 48 32 52 37
rect 78 32 82 39
rect 48 27 63 32
rect 67 27 82 32
rect 38 21 65 22
rect 38 19 61 21
rect 63 19 65 21
rect 38 18 65 19
rect 80 21 84 23
rect 80 19 81 21
rect 83 19 84 21
rect 80 12 84 19
rect -2 7 92 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 92 7
rect -2 0 92 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 24 95 30 97
rect 24 93 26 95
rect 28 93 30 95
rect 24 91 30 93
<< nmos >>
rect 25 17 27 36
rect 47 17 49 34
rect 55 17 57 34
rect 67 17 69 34
rect 75 17 77 34
<< pmos >>
rect 11 55 13 93
rect 41 55 43 93
rect 53 55 55 93
rect 65 55 67 93
rect 77 55 79 93
<< polyct1 >>
rect 28 48 30 50
rect 69 48 71 50
rect 47 39 49 41
rect 59 39 61 41
rect 79 39 81 41
<< ndifct1 >>
rect 19 32 21 34
rect 19 24 21 26
rect 31 29 33 31
rect 31 19 33 21
rect 61 19 63 21
rect 81 19 83 21
<< ntiect1 >>
rect 26 93 28 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 5 69 7 71
rect 35 79 37 81
rect 17 67 19 69
rect 17 59 19 61
rect 47 69 49 71
rect 59 79 61 81
rect 71 89 73 91
rect 83 78 85 80
rect 83 70 85 72
<< labels >>
rlabel polyct1 29 49 29 49 6 zn
rlabel pdifct1 36 80 36 80 6 n3
rlabel ndifct1 62 20 62 20 6 zn
rlabel pdifct1 48 70 48 70 6 zn
rlabel pdifct1 60 80 60 80 6 n3
rlabel pdifct1 84 71 84 71 6 n3
rlabel pdifct1 84 79 84 79 6 n3
rlabel alu1 10 60 10 60 6 z
rlabel alu1 20 45 20 45 6 z
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 60 30 60 30 6 b1
rlabel alu1 50 40 50 40 6 b1
rlabel alu1 60 55 60 55 6 b2
rlabel alu1 50 60 50 60 6 b2
rlabel alu1 45 94 45 94 6 vdd
rlabel alu1 70 30 70 30 6 a1
rlabel polyct1 80 40 80 40 6 a1
rlabel alu1 70 55 70 55 6 a2
rlabel alu1 80 60 80 60 6 a2
<< end >>
