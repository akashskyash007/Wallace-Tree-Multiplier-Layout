magic
tech scmos
timestamp 1199203641
<< ab >>
rect 0 0 104 80
<< nwell >>
rect -5 36 109 88
<< pwell >>
rect -5 -8 109 36
<< poly >>
rect 63 70 65 74
rect 73 70 75 74
rect 83 70 85 74
rect 93 70 95 74
rect 9 65 21 67
rect 9 62 11 65
rect 19 62 21 65
rect 29 65 50 67
rect 29 62 31 65
rect 39 62 41 65
rect 48 63 50 65
rect 48 61 54 63
rect 48 59 50 61
rect 52 59 54 61
rect 48 57 54 59
rect 63 47 65 50
rect 73 47 75 50
rect 83 47 85 50
rect 93 47 95 50
rect 55 45 79 47
rect 9 38 11 42
rect 19 39 21 42
rect 18 37 24 39
rect 29 38 31 42
rect 18 35 20 37
rect 22 35 24 37
rect 39 35 41 42
rect 11 30 13 34
rect 18 33 24 35
rect 18 30 20 33
rect 28 30 30 34
rect 35 33 41 35
rect 35 30 37 33
rect 55 30 57 45
rect 73 43 75 45
rect 77 43 79 45
rect 73 41 79 43
rect 83 45 95 47
rect 83 43 91 45
rect 93 43 95 45
rect 83 41 95 43
rect 63 37 69 39
rect 63 35 65 37
rect 67 35 69 37
rect 63 33 69 35
rect 65 30 67 33
rect 75 30 77 41
rect 85 30 87 41
rect 11 8 13 17
rect 18 14 20 17
rect 28 14 30 17
rect 18 12 30 14
rect 35 8 37 17
rect 55 15 57 20
rect 85 15 87 20
rect 11 6 37 8
rect 65 6 67 10
rect 75 6 77 10
<< ndif >>
rect 3 21 11 30
rect 3 19 6 21
rect 8 19 11 21
rect 3 17 11 19
rect 13 17 18 30
rect 20 28 28 30
rect 20 26 23 28
rect 25 26 28 28
rect 20 21 28 26
rect 20 19 23 21
rect 25 19 28 21
rect 20 17 28 19
rect 30 17 35 30
rect 37 21 55 30
rect 37 19 40 21
rect 42 20 55 21
rect 57 28 65 30
rect 57 26 60 28
rect 62 26 65 28
rect 57 20 65 26
rect 42 19 53 20
rect 37 17 53 19
rect 60 10 65 20
rect 67 28 75 30
rect 67 26 70 28
rect 72 26 75 28
rect 67 21 75 26
rect 67 19 70 21
rect 72 19 75 21
rect 67 10 75 19
rect 77 28 85 30
rect 77 26 80 28
rect 82 26 85 28
rect 77 20 85 26
rect 87 20 96 30
rect 77 10 82 20
rect 89 19 96 20
rect 89 17 91 19
rect 93 17 96 19
rect 89 15 96 17
<< pdif >>
rect 56 68 63 70
rect 56 66 58 68
rect 60 66 63 68
rect 4 55 9 62
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 60 19 62
rect 11 58 14 60
rect 16 58 19 60
rect 11 53 19 58
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 53 29 62
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 46 39 62
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 55 46 62
rect 41 53 48 55
rect 41 51 44 53
rect 46 51 48 53
rect 41 49 48 51
rect 56 50 63 66
rect 65 54 73 70
rect 65 52 68 54
rect 70 52 73 54
rect 65 50 73 52
rect 75 68 83 70
rect 75 66 78 68
rect 80 66 83 68
rect 75 50 83 66
rect 85 61 93 70
rect 85 59 88 61
rect 90 59 93 61
rect 85 50 93 59
rect 95 68 102 70
rect 95 66 98 68
rect 100 66 102 68
rect 95 50 102 66
rect 41 42 46 49
<< alu1 >>
rect -2 81 106 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 106 81
rect -2 68 106 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 22 53 48 54
rect 22 51 24 53
rect 26 51 44 53
rect 46 51 48 53
rect 22 50 48 51
rect 22 46 27 50
rect 2 44 4 46
rect 6 44 24 46
rect 26 44 27 46
rect 2 42 27 44
rect 82 46 86 55
rect 73 45 86 46
rect 73 43 75 45
rect 77 43 86 45
rect 73 42 86 43
rect 90 45 94 47
rect 90 43 91 45
rect 93 43 94 45
rect 2 30 6 42
rect 90 38 94 43
rect 2 28 50 30
rect 2 26 23 28
rect 25 26 50 28
rect 22 21 26 26
rect 22 19 23 21
rect 25 19 26 21
rect 22 17 26 19
rect 46 22 50 26
rect 63 37 94 38
rect 63 35 65 37
rect 67 35 94 37
rect 63 34 94 35
rect 69 28 74 30
rect 69 26 70 28
rect 72 26 74 28
rect 69 22 74 26
rect 46 21 74 22
rect 46 19 70 21
rect 72 19 74 21
rect 46 18 74 19
rect -2 1 106 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 106 1
rect -2 -2 106 -1
<< ptie >>
rect 0 1 104 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 104 1
rect 0 -3 104 -1
<< ntie >>
rect 0 81 104 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 104 81
rect 0 77 104 79
<< nmos >>
rect 11 17 13 30
rect 18 17 20 30
rect 28 17 30 30
rect 35 17 37 30
rect 55 20 57 30
rect 65 10 67 30
rect 75 10 77 30
rect 85 20 87 30
<< pmos >>
rect 9 42 11 62
rect 19 42 21 62
rect 29 42 31 62
rect 39 42 41 62
rect 63 50 65 70
rect 73 50 75 70
rect 83 50 85 70
rect 93 50 95 70
<< polyct0 >>
rect 50 59 52 61
rect 20 35 22 37
<< polyct1 >>
rect 75 43 77 45
rect 91 43 93 45
rect 65 35 67 37
<< ndifct0 >>
rect 6 19 8 21
rect 40 19 42 21
rect 60 26 62 28
rect 80 26 82 28
rect 91 17 93 19
<< ndifct1 >>
rect 23 26 25 28
rect 23 19 25 21
rect 70 26 72 28
rect 70 19 72 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
<< pdifct0 >>
rect 58 66 60 68
rect 14 58 16 60
rect 14 51 16 53
rect 34 44 36 46
rect 68 52 70 54
rect 78 66 80 68
rect 88 59 90 61
rect 98 66 100 68
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 51 26 53
rect 24 44 26 46
rect 44 51 46 53
<< alu0 >>
rect 56 66 58 68
rect 60 66 62 68
rect 56 65 62 66
rect 76 66 78 68
rect 80 66 82 68
rect 76 65 82 66
rect 96 66 98 68
rect 100 66 102 68
rect 96 65 102 66
rect 12 61 102 62
rect 12 60 50 61
rect 12 58 14 60
rect 16 59 50 60
rect 52 59 88 61
rect 90 59 102 61
rect 16 58 102 59
rect 12 53 18 58
rect 66 54 72 55
rect 12 51 14 53
rect 16 51 18 53
rect 12 50 18 51
rect 54 52 68 54
rect 70 52 72 54
rect 54 50 72 52
rect 32 46 38 47
rect 32 44 34 46
rect 36 44 38 46
rect 32 42 38 44
rect 54 42 58 50
rect 32 38 58 42
rect 18 37 38 38
rect 18 35 20 37
rect 22 35 38 37
rect 18 34 38 35
rect 4 21 10 22
rect 4 19 6 21
rect 8 19 10 21
rect 4 12 10 19
rect 39 21 43 23
rect 39 19 40 21
rect 42 19 43 21
rect 39 12 43 19
rect 54 29 58 38
rect 54 28 64 29
rect 54 26 60 28
rect 62 26 64 28
rect 54 25 64 26
rect 98 29 102 58
rect 78 28 102 29
rect 78 26 80 28
rect 82 26 102 28
rect 78 25 102 26
rect 90 19 94 21
rect 90 17 91 19
rect 93 17 94 19
rect 90 12 94 17
<< labels >>
rlabel alu0 15 56 15 56 6 an
rlabel alu0 28 36 28 36 6 bn
rlabel alu0 59 27 59 27 6 bn
rlabel alu0 45 40 45 40 6 bn
rlabel alu0 63 52 63 52 6 bn
rlabel alu0 90 27 90 27 6 an
rlabel alu0 57 60 57 60 6 an
rlabel alu1 20 28 20 28 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 4 44 4 44 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 28 28 28 28 6 z
rlabel alu1 44 28 44 28 6 z
rlabel alu1 36 28 36 28 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 52 6 52 6 6 vss
rlabel alu1 60 20 60 20 6 z
rlabel alu1 68 20 68 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 76 36 76 36 6 a
rlabel alu1 68 36 68 36 6 a
rlabel polyct1 76 44 76 44 6 b
rlabel alu1 52 74 52 74 6 vdd
rlabel alu1 84 36 84 36 6 a
rlabel polyct1 92 44 92 44 6 a
rlabel alu1 84 52 84 52 6 b
<< end >>
