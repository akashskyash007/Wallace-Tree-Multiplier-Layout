magic
tech scmos
timestamp 1199203379
<< ab >>
rect 0 0 48 72
<< nwell >>
rect -5 32 53 77
<< pwell >>
rect -5 -5 53 32
<< alu1 >>
rect -2 67 50 72
rect -2 65 8 67
rect 10 65 15 67
rect 17 65 23 67
rect 25 65 31 67
rect 33 65 38 67
rect 40 65 50 67
rect -2 64 50 65
rect -2 7 50 8
rect -2 5 8 7
rect 10 5 15 7
rect 17 5 23 7
rect 25 5 31 7
rect 33 5 38 7
rect 40 5 50 7
rect -2 0 50 5
<< ptie >>
rect 6 7 42 26
rect 6 5 8 7
rect 10 5 15 7
rect 17 5 23 7
rect 25 5 31 7
rect 33 5 38 7
rect 40 5 42 7
rect 6 3 42 5
<< ntie >>
rect 6 67 42 69
rect 6 65 8 67
rect 10 65 15 67
rect 17 65 23 67
rect 25 65 31 67
rect 33 65 38 67
rect 40 65 42 67
rect 6 38 42 65
<< ntiect1 >>
rect 8 65 10 67
rect 15 65 17 67
rect 23 65 25 67
rect 31 65 33 67
rect 38 65 40 67
<< ptiect1 >>
rect 8 5 10 7
rect 15 5 17 7
rect 23 5 25 7
rect 31 5 33 7
rect 38 5 40 7
<< labels >>
rlabel alu1 24 4 24 4 6 vss
rlabel alu1 24 68 24 68 6 vdd
<< end >>
