magic
tech scmos
timestamp 1199203263
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 9 66 11 70
rect 29 68 55 70
rect 22 60 24 65
rect 29 60 31 68
rect 36 60 38 64
rect 46 57 48 62
rect 53 57 55 68
rect 60 57 62 61
rect 9 35 11 38
rect 22 35 24 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 9 26 11 29
rect 20 18 22 29
rect 29 27 31 38
rect 36 35 38 38
rect 46 35 48 38
rect 36 33 48 35
rect 53 33 55 38
rect 60 35 62 38
rect 60 33 67 35
rect 44 27 48 33
rect 60 31 63 33
rect 65 31 67 33
rect 60 29 67 31
rect 29 25 39 27
rect 29 23 35 25
rect 37 23 39 25
rect 29 21 39 23
rect 44 25 50 27
rect 44 23 46 25
rect 48 23 50 25
rect 44 21 50 23
rect 30 18 32 21
rect 44 18 46 21
rect 9 7 11 12
rect 20 5 22 10
rect 30 5 32 10
rect 44 5 46 10
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 12 9 15
rect 11 18 18 26
rect 11 15 20 18
rect 11 13 15 15
rect 17 13 20 15
rect 11 12 20 13
rect 13 10 20 12
rect 22 16 30 18
rect 22 14 25 16
rect 27 14 30 16
rect 22 10 30 14
rect 32 10 44 18
rect 46 16 53 18
rect 46 14 49 16
rect 51 14 53 16
rect 46 12 53 14
rect 46 10 51 12
rect 34 7 42 10
rect 34 5 37 7
rect 39 5 42 7
rect 34 3 42 5
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 20 66
rect 11 62 16 64
rect 18 62 20 64
rect 11 60 20 62
rect 11 57 22 60
rect 11 55 16 57
rect 18 55 22 57
rect 11 38 22 55
rect 24 38 29 60
rect 31 38 36 60
rect 38 57 43 60
rect 38 55 46 57
rect 38 53 41 55
rect 43 53 46 55
rect 38 48 46 53
rect 38 46 41 48
rect 43 46 46 48
rect 38 38 46 46
rect 48 38 53 57
rect 55 38 60 57
rect 62 55 70 57
rect 62 53 65 55
rect 67 53 70 55
rect 62 48 70 53
rect 62 46 65 48
rect 67 46 70 48
rect 62 38 70 46
<< alu1 >>
rect -2 67 74 72
rect -2 65 65 67
rect 67 65 74 67
rect -2 64 74 65
rect 2 49 14 51
rect 2 47 4 49
rect 6 47 14 49
rect 2 45 14 47
rect 2 42 6 45
rect 2 40 4 42
rect 2 26 6 40
rect 26 38 63 42
rect 26 35 30 38
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 17 7 22
rect 20 33 30 35
rect 57 34 63 38
rect 20 31 21 33
rect 23 31 30 33
rect 20 29 30 31
rect 34 30 47 34
rect 57 33 67 34
rect 57 31 63 33
rect 65 31 67 33
rect 57 30 67 31
rect 34 25 38 30
rect 34 23 35 25
rect 37 23 38 25
rect 34 21 38 23
rect 44 25 63 26
rect 44 23 46 25
rect 48 23 63 25
rect 44 22 63 23
rect 2 15 4 17
rect 6 15 7 17
rect 2 13 7 15
rect 57 14 63 22
rect -2 7 74 8
rect -2 5 37 7
rect 39 5 65 7
rect 67 5 74 7
rect -2 0 74 5
<< ptie >>
rect 63 7 69 24
rect 63 5 65 7
rect 67 5 69 7
rect 63 3 69 5
<< ntie >>
rect 63 67 69 69
rect 63 65 65 67
rect 67 65 69 67
rect 63 63 69 65
<< nmos >>
rect 9 12 11 26
rect 20 10 22 18
rect 30 10 32 18
rect 44 10 46 18
<< pmos >>
rect 9 38 11 66
rect 22 38 24 60
rect 29 38 31 60
rect 36 38 38 60
rect 46 38 48 57
rect 53 38 55 57
rect 60 38 62 57
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 21 31 23 33
rect 63 31 65 33
rect 35 23 37 25
rect 46 23 48 25
<< ndifct0 >>
rect 15 13 17 15
rect 25 14 27 16
rect 49 14 51 16
<< ndifct1 >>
rect 4 22 6 24
rect 4 15 6 17
rect 37 5 39 7
<< ntiect1 >>
rect 65 65 67 67
<< ptiect1 >>
rect 65 5 67 7
<< pdifct0 >>
rect 16 62 18 64
rect 16 55 18 57
rect 41 53 43 55
rect 41 46 43 48
rect 65 53 67 55
rect 65 46 67 48
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
<< alu0 >>
rect 14 62 16 64
rect 18 62 20 64
rect 14 57 20 62
rect 14 55 16 57
rect 18 55 20 57
rect 14 54 20 55
rect 39 55 45 56
rect 39 53 41 55
rect 43 53 45 55
rect 39 49 45 53
rect 18 48 45 49
rect 18 46 41 48
rect 43 46 45 48
rect 18 45 45 46
rect 63 55 69 64
rect 63 53 65 55
rect 67 53 69 55
rect 63 48 69 53
rect 63 46 65 48
rect 67 46 69 48
rect 63 45 69 46
rect 6 38 7 45
rect 18 42 22 45
rect 10 38 22 42
rect 10 33 14 38
rect 10 31 11 33
rect 13 31 14 33
rect 10 25 14 31
rect 10 21 27 25
rect 23 17 27 21
rect 23 16 53 17
rect 13 15 19 16
rect 13 13 15 15
rect 17 13 19 15
rect 23 14 25 16
rect 27 14 49 16
rect 51 14 53 16
rect 23 13 53 14
rect 13 8 19 13
<< labels >>
rlabel alu0 12 31 12 31 6 zn
rlabel alu0 42 50 42 50 6 zn
rlabel alu0 31 47 31 47 6 zn
rlabel alu0 38 15 38 15 6 zn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 32 28 32 6 a
rlabel alu1 36 4 36 4 6 vss
rlabel polyct1 36 24 36 24 6 b
rlabel alu1 44 32 44 32 6 b
rlabel alu1 52 24 52 24 6 c
rlabel alu1 44 40 44 40 6 a
rlabel alu1 52 40 52 40 6 a
rlabel alu1 36 40 36 40 6 a
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 20 60 20 6 c
rlabel alu1 60 36 60 36 6 a
<< end >>
