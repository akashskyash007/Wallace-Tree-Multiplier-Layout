magic
tech scmos
timestamp 1199202903
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 12 66 14 70
rect 19 66 21 70
rect 12 35 14 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 32 21 38
rect 19 30 25 32
rect 10 20 12 29
rect 19 28 21 30
rect 23 28 25 30
rect 19 26 25 28
rect 21 23 23 26
rect 10 7 12 12
rect 21 11 23 15
<< ndif >>
rect 16 20 21 23
rect 2 12 10 20
rect 12 16 21 20
rect 12 14 15 16
rect 17 15 21 16
rect 23 19 30 23
rect 23 17 26 19
rect 28 17 30 19
rect 23 15 30 17
rect 17 14 19 15
rect 12 12 19 14
rect 2 7 8 12
rect 2 5 4 7
rect 6 5 8 7
rect 2 3 8 5
<< pdif >>
rect 7 59 12 66
rect 5 57 12 59
rect 5 55 7 57
rect 9 55 12 57
rect 5 50 12 55
rect 5 48 7 50
rect 9 48 12 50
rect 5 46 12 48
rect 7 38 12 46
rect 14 38 19 66
rect 21 64 30 66
rect 21 62 26 64
rect 28 62 30 64
rect 21 57 30 62
rect 21 55 26 57
rect 28 55 30 57
rect 21 38 30 55
<< alu1 >>
rect -2 64 34 72
rect 5 57 11 58
rect 5 55 7 57
rect 9 55 11 57
rect 5 51 11 55
rect 2 50 11 51
rect 2 48 7 50
rect 9 48 11 50
rect 2 47 11 48
rect 2 19 6 47
rect 18 39 22 43
rect 10 35 22 39
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 26 31 30 35
rect 10 29 14 31
rect 18 30 30 31
rect 18 28 21 30
rect 23 28 30 30
rect 18 27 30 28
rect 18 21 22 27
rect 2 17 14 19
rect 2 16 19 17
rect 2 14 15 16
rect 17 14 19 16
rect 2 13 19 14
rect -2 7 34 8
rect -2 5 4 7
rect 6 5 25 7
rect 27 5 34 7
rect -2 0 34 5
<< ptie >>
rect 23 7 29 9
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< nmos >>
rect 10 12 12 20
rect 21 15 23 23
<< pmos >>
rect 12 38 14 66
rect 19 38 21 66
<< polyct1 >>
rect 11 31 13 33
rect 21 28 23 30
<< ndifct0 >>
rect 26 17 28 19
<< ndifct1 >>
rect 15 14 17 16
rect 4 5 6 7
<< ptiect1 >>
rect 25 5 27 7
<< pdifct0 >>
rect 26 62 28 64
rect 26 55 28 57
<< pdifct1 >>
rect 7 55 9 57
rect 7 48 9 50
<< alu0 >>
rect 25 62 26 64
rect 28 62 29 64
rect 25 57 29 62
rect 25 55 26 57
rect 28 55 29 57
rect 25 53 29 55
rect 25 19 29 21
rect 25 17 26 19
rect 28 17 29 19
rect 25 8 29 17
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 24 20 24 6 a
rlabel alu1 20 40 20 40 6 b
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 32 28 32 6 a
<< end >>
