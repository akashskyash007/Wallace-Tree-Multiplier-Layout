magic
tech scmos
timestamp 1199201748
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 20 62 22 67
rect 30 62 32 67
rect 42 62 44 67
rect 52 62 54 67
rect 9 56 11 61
rect 9 35 11 44
rect 20 35 22 52
rect 30 49 32 52
rect 30 47 38 49
rect 30 45 34 47
rect 36 45 38 47
rect 30 43 38 45
rect 42 43 44 52
rect 9 33 16 35
rect 9 31 12 33
rect 14 31 16 33
rect 9 29 16 31
rect 20 33 28 35
rect 20 31 24 33
rect 26 31 28 33
rect 20 29 28 31
rect 9 24 11 29
rect 25 26 27 29
rect 32 26 34 43
rect 42 41 48 43
rect 42 39 44 41
rect 46 39 48 41
rect 39 37 48 39
rect 39 26 41 37
rect 52 35 54 52
rect 52 33 58 35
rect 52 31 54 33
rect 56 31 58 33
rect 46 29 58 31
rect 46 26 48 29
rect 9 13 11 18
rect 25 9 27 14
rect 32 9 34 14
rect 39 9 41 14
rect 46 9 48 14
<< ndif >>
rect 13 24 25 26
rect 2 22 9 24
rect 2 20 4 22
rect 6 20 9 22
rect 2 18 9 20
rect 11 18 25 24
rect 13 14 25 18
rect 27 14 32 26
rect 34 14 39 26
rect 41 14 46 26
rect 48 20 53 26
rect 48 18 55 20
rect 48 16 51 18
rect 53 16 55 18
rect 48 14 55 16
rect 13 7 23 14
rect 13 5 17 7
rect 19 5 23 7
rect 13 3 23 5
<< pdif >>
rect 34 67 40 69
rect 34 65 36 67
rect 38 65 40 67
rect 34 62 40 65
rect 13 58 20 62
rect 13 56 15 58
rect 17 56 20 58
rect 4 50 9 56
rect 2 48 9 50
rect 2 46 4 48
rect 6 46 9 48
rect 2 44 9 46
rect 11 52 20 56
rect 22 58 30 62
rect 22 56 25 58
rect 27 56 30 58
rect 22 52 30 56
rect 32 52 42 62
rect 44 58 52 62
rect 44 56 47 58
rect 49 56 52 58
rect 44 52 52 56
rect 54 60 61 62
rect 54 58 57 60
rect 59 58 61 60
rect 54 52 61 58
rect 11 44 18 52
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 36 67
rect 38 65 66 67
rect -2 64 66 65
rect 2 48 7 59
rect 2 46 4 48
rect 6 46 7 48
rect 2 44 7 46
rect 33 47 47 50
rect 2 22 6 44
rect 33 45 34 47
rect 36 46 47 47
rect 36 45 37 46
rect 33 42 37 45
rect 58 42 62 51
rect 25 38 37 42
rect 41 41 62 42
rect 41 39 44 41
rect 46 39 62 41
rect 41 38 62 39
rect 22 33 31 34
rect 22 31 24 33
rect 26 31 31 33
rect 22 30 31 31
rect 41 33 62 34
rect 41 31 54 33
rect 56 31 62 33
rect 41 30 62 31
rect 2 20 4 22
rect 2 19 6 20
rect 2 13 14 19
rect 26 26 31 30
rect 26 22 39 26
rect 58 13 62 30
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 17 7
rect 19 5 57 7
rect 59 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 55 7 61 9
rect 55 5 57 7
rect 59 5 61 7
rect 55 3 61 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 18 11 24
rect 25 14 27 26
rect 32 14 34 26
rect 39 14 41 26
rect 46 14 48 26
<< pmos >>
rect 9 44 11 56
rect 20 52 22 62
rect 30 52 32 62
rect 42 52 44 62
rect 52 52 54 62
<< polyct0 >>
rect 12 31 14 33
<< polyct1 >>
rect 34 45 36 47
rect 24 31 26 33
rect 44 39 46 41
rect 54 31 56 33
<< ndifct0 >>
rect 51 16 53 18
<< ndifct1 >>
rect 4 20 6 22
rect 17 5 19 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
rect 57 5 59 7
<< pdifct0 >>
rect 15 56 17 58
rect 25 56 27 58
rect 47 56 49 58
rect 57 58 59 60
<< pdifct1 >>
rect 36 65 38 67
rect 4 46 6 48
<< alu0 >>
rect 14 58 18 64
rect 56 60 60 64
rect 14 56 15 58
rect 17 56 18 58
rect 14 54 18 56
rect 23 58 51 59
rect 23 56 25 58
rect 27 56 47 58
rect 49 56 51 58
rect 56 58 57 60
rect 59 58 60 60
rect 56 56 60 58
rect 23 55 51 56
rect 23 50 27 55
rect 14 46 27 50
rect 14 34 18 46
rect 10 33 18 34
rect 10 31 12 33
rect 14 31 18 33
rect 10 30 18 31
rect 14 27 18 30
rect 6 19 7 24
rect 14 23 22 27
rect 18 17 22 23
rect 50 18 54 20
rect 50 17 51 18
rect 18 16 51 17
rect 53 16 54 18
rect 18 13 54 16
<< labels >>
rlabel alu0 16 36 16 36 6 zn
rlabel alu0 52 16 52 16 6 zn
rlabel alu0 37 57 37 57 6 zn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 32 44 32 6 d
rlabel alu1 44 40 44 40 6 c
rlabel alu1 36 48 36 48 6 b
rlabel alu1 44 48 44 48 6 b
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 60 20 60 20 6 d
rlabel alu1 52 32 52 32 6 d
rlabel alu1 52 40 52 40 6 c
rlabel alu1 60 48 60 48 6 c
<< end >>
