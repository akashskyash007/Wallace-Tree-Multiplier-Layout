magic
tech scmos
timestamp 1199203184
<< ab >>
rect 0 0 136 72
<< nwell >>
rect -5 32 141 77
<< pwell >>
rect -5 -5 141 32
<< poly >>
rect 31 66 33 70
rect 39 66 41 70
rect 47 66 49 70
rect 57 66 59 70
rect 65 66 67 70
rect 73 66 75 70
rect 83 66 85 70
rect 91 66 93 70
rect 99 66 101 70
rect 109 66 111 70
rect 116 66 118 70
rect 123 66 125 70
rect 9 57 11 61
rect 19 59 21 64
rect 9 35 11 38
rect 19 35 21 38
rect 31 35 33 38
rect 39 35 41 38
rect 47 35 49 38
rect 57 35 59 38
rect 65 35 67 38
rect 73 35 75 38
rect 83 35 85 38
rect 91 35 93 38
rect 99 35 101 38
rect 109 35 111 38
rect 9 33 21 35
rect 9 31 14 33
rect 16 31 21 33
rect 9 29 21 31
rect 26 33 33 35
rect 26 31 28 33
rect 30 31 33 33
rect 26 29 33 31
rect 37 33 43 35
rect 47 33 59 35
rect 63 33 69 35
rect 37 31 39 33
rect 41 31 43 33
rect 37 29 43 31
rect 49 31 51 33
rect 53 31 55 33
rect 49 29 55 31
rect 63 31 65 33
rect 67 31 69 33
rect 63 29 69 31
rect 73 33 85 35
rect 89 33 95 35
rect 73 31 75 33
rect 77 31 79 33
rect 73 29 79 31
rect 89 31 91 33
rect 93 31 95 33
rect 89 29 95 31
rect 99 33 111 35
rect 99 32 105 33
rect 99 30 101 32
rect 103 30 105 32
rect 9 26 11 29
rect 19 26 21 29
rect 29 25 33 29
rect 51 26 53 29
rect 29 23 43 25
rect 29 20 31 23
rect 41 20 43 23
rect 9 3 11 8
rect 19 3 21 8
rect 29 3 31 8
rect 67 24 69 29
rect 89 24 91 29
rect 67 22 91 24
rect 67 19 69 22
rect 77 19 79 22
rect 89 19 91 22
rect 99 28 105 30
rect 116 29 118 38
rect 123 35 125 38
rect 123 33 134 35
rect 123 31 130 33
rect 132 31 134 33
rect 123 29 134 31
rect 99 19 101 28
rect 113 27 119 29
rect 113 25 115 27
rect 117 25 119 27
rect 113 23 119 25
rect 125 19 127 29
rect 41 2 43 6
rect 51 2 53 6
rect 67 4 69 9
rect 77 4 79 9
rect 89 2 91 7
rect 99 2 101 7
rect 125 8 127 13
<< ndif >>
rect 4 19 9 26
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 8 9 13
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 8 19 22
rect 21 20 26 26
rect 46 20 51 26
rect 21 17 29 20
rect 21 15 24 17
rect 26 15 29 17
rect 21 8 29 15
rect 31 10 41 20
rect 31 8 35 10
rect 37 8 41 10
rect 33 6 41 8
rect 43 17 51 20
rect 43 15 46 17
rect 48 15 51 17
rect 43 6 51 15
rect 53 19 65 26
rect 53 10 67 19
rect 53 8 59 10
rect 61 9 67 10
rect 69 17 77 19
rect 69 15 72 17
rect 74 15 77 17
rect 69 9 77 15
rect 79 9 89 19
rect 61 8 65 9
rect 53 6 65 8
rect 81 7 89 9
rect 91 17 99 19
rect 91 15 94 17
rect 96 15 99 17
rect 91 7 99 15
rect 101 7 109 19
rect 118 17 125 19
rect 118 15 120 17
rect 122 15 125 17
rect 118 13 125 15
rect 127 17 134 19
rect 127 15 130 17
rect 132 15 134 17
rect 127 13 134 15
rect 81 5 83 7
rect 85 5 87 7
rect 81 3 87 5
rect 103 5 105 7
rect 107 5 109 7
rect 103 3 109 5
<< pdif >>
rect 23 64 31 66
rect 23 62 25 64
rect 27 62 31 64
rect 23 59 31 62
rect 14 57 19 59
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 38 9 53
rect 11 55 19 57
rect 11 53 14 55
rect 16 53 19 55
rect 11 48 19 53
rect 11 46 14 48
rect 16 46 19 48
rect 11 38 19 46
rect 21 38 31 59
rect 33 38 39 66
rect 41 38 47 66
rect 49 57 57 66
rect 49 55 52 57
rect 54 55 57 57
rect 49 38 57 55
rect 59 38 65 66
rect 67 38 73 66
rect 75 64 83 66
rect 75 62 78 64
rect 80 62 83 64
rect 75 38 83 62
rect 85 38 91 66
rect 93 38 99 66
rect 101 57 109 66
rect 101 55 104 57
rect 106 55 109 57
rect 101 38 109 55
rect 111 38 116 66
rect 118 38 123 66
rect 125 64 134 66
rect 125 62 130 64
rect 132 62 134 64
rect 125 57 134 62
rect 125 55 130 57
rect 132 55 134 57
rect 125 38 134 55
<< alu1 >>
rect -2 67 138 72
rect -2 65 5 67
rect 7 65 138 67
rect -2 64 138 65
rect 16 57 108 58
rect 16 55 52 57
rect 54 55 104 57
rect 106 55 108 57
rect 16 54 108 55
rect 2 25 6 47
rect 25 46 134 50
rect 17 35 23 42
rect 10 33 23 35
rect 10 31 14 33
rect 16 31 23 33
rect 10 29 23 31
rect 41 38 69 42
rect 41 35 45 38
rect 34 33 45 35
rect 34 31 39 33
rect 41 31 45 33
rect 34 30 45 31
rect 49 33 55 34
rect 49 31 51 33
rect 53 31 55 33
rect 2 24 18 25
rect 2 22 14 24
rect 16 22 18 24
rect 2 21 18 22
rect 34 21 38 30
rect 49 26 55 31
rect 63 33 69 38
rect 63 31 65 33
rect 67 31 69 33
rect 63 30 69 31
rect 73 33 79 46
rect 73 31 75 33
rect 77 31 79 33
rect 73 30 79 31
rect 89 38 119 42
rect 89 33 95 38
rect 89 31 91 33
rect 93 31 95 33
rect 89 30 95 31
rect 102 32 106 34
rect 103 30 106 32
rect 102 26 106 30
rect 49 22 106 26
rect 113 27 119 38
rect 129 33 134 46
rect 129 31 130 33
rect 132 31 134 33
rect 129 29 134 31
rect 113 25 115 27
rect 117 25 119 27
rect 113 22 119 25
rect -2 7 138 8
rect -2 5 83 7
rect 85 5 105 7
rect 107 5 115 7
rect 117 5 138 7
rect -2 0 138 5
<< ptie >>
rect 113 7 119 9
rect 113 5 115 7
rect 117 5 119 7
rect 113 3 119 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 8 11 26
rect 19 8 21 26
rect 29 8 31 20
rect 41 6 43 20
rect 51 6 53 26
rect 67 9 69 19
rect 77 9 79 19
rect 89 7 91 19
rect 99 7 101 19
rect 125 13 127 19
<< pmos >>
rect 9 38 11 57
rect 19 38 21 59
rect 31 38 33 66
rect 39 38 41 66
rect 47 38 49 66
rect 57 38 59 66
rect 65 38 67 66
rect 73 38 75 66
rect 83 38 85 66
rect 91 38 93 66
rect 99 38 101 66
rect 109 38 111 66
rect 116 38 118 66
rect 123 38 125 66
<< polyct0 >>
rect 28 31 30 33
rect 101 30 102 32
<< polyct1 >>
rect 14 31 16 33
rect 39 31 41 33
rect 51 31 53 33
rect 65 31 67 33
rect 75 31 77 33
rect 91 31 93 33
rect 102 30 103 32
rect 130 31 132 33
rect 115 25 117 27
<< ndifct0 >>
rect 4 15 6 17
rect 24 15 26 17
rect 35 8 37 10
rect 46 15 48 17
rect 59 8 61 10
rect 72 15 74 17
rect 94 15 96 17
rect 120 15 122 17
rect 130 15 132 17
<< ndifct1 >>
rect 14 22 16 24
rect 83 5 85 7
rect 105 5 107 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 115 5 117 7
<< pdifct0 >>
rect 25 62 27 64
rect 4 53 6 55
rect 14 53 16 55
rect 14 46 16 48
rect 78 62 80 64
rect 130 62 132 64
rect 130 55 132 57
<< pdifct1 >>
rect 52 55 54 57
rect 104 55 106 57
<< alu0 >>
rect 2 55 8 64
rect 23 62 25 64
rect 27 62 29 64
rect 23 61 29 62
rect 76 62 78 64
rect 80 62 82 64
rect 76 61 82 62
rect 128 62 130 64
rect 132 62 134 64
rect 2 53 4 55
rect 6 53 8 55
rect 2 52 8 53
rect 13 55 16 58
rect 13 53 14 55
rect 128 57 134 62
rect 128 55 130 57
rect 132 55 134 57
rect 128 54 134 55
rect 16 53 18 54
rect 13 49 18 53
rect 2 48 18 49
rect 2 47 14 48
rect 6 46 14 47
rect 16 46 18 48
rect 6 45 18 46
rect 27 33 31 46
rect 27 31 28 33
rect 30 31 31 33
rect 27 29 31 31
rect 100 32 102 34
rect 100 30 101 32
rect 100 26 102 30
rect 2 17 124 18
rect 2 15 4 17
rect 6 15 24 17
rect 26 15 46 17
rect 48 15 72 17
rect 74 15 94 17
rect 96 15 120 17
rect 122 15 124 17
rect 2 14 124 15
rect 129 17 133 19
rect 129 15 130 17
rect 132 15 133 17
rect 33 10 39 11
rect 33 8 35 10
rect 37 8 39 10
rect 57 10 63 11
rect 57 8 59 10
rect 61 8 63 10
rect 129 8 133 15
<< labels >>
rlabel alu0 63 16 63 16 6 n3
rlabel alu1 12 32 12 32 6 b
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 36 20 36 6 b
rlabel alu1 20 56 20 56 6 z
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 44 40 44 40 6 a2
rlabel alu1 28 48 28 48 6 a1
rlabel alu1 36 48 36 48 6 a1
rlabel alu1 44 48 44 48 6 a1
rlabel alu1 36 56 36 56 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 68 4 68 4 6 vss
rlabel alu1 60 24 60 24 6 a3
rlabel alu1 68 24 68 24 6 a3
rlabel alu1 76 24 76 24 6 a3
rlabel alu1 52 28 52 28 6 a3
rlabel alu1 52 40 52 40 6 a2
rlabel alu1 76 40 76 40 6 a1
rlabel alu1 60 40 60 40 6 a2
rlabel alu1 52 48 52 48 6 a1
rlabel alu1 60 48 60 48 6 a1
rlabel alu1 68 48 68 48 6 a1
rlabel alu1 60 56 60 56 6 z
rlabel alu1 68 56 68 56 6 z
rlabel alu1 76 56 76 56 6 z
rlabel alu1 52 56 52 56 6 z
rlabel alu1 68 68 68 68 6 vdd
rlabel alu1 84 24 84 24 6 a3
rlabel alu1 100 24 100 24 6 a3
rlabel alu1 92 24 92 24 6 a3
rlabel alu1 100 40 100 40 6 a2
rlabel alu1 108 40 108 40 6 a2
rlabel alu1 92 36 92 36 6 a2
rlabel alu1 84 48 84 48 6 a1
rlabel alu1 100 48 100 48 6 a1
rlabel alu1 108 48 108 48 6 a1
rlabel alu1 92 48 92 48 6 a1
rlabel alu1 100 56 100 56 6 z
rlabel alu1 92 56 92 56 6 z
rlabel alu1 84 56 84 56 6 z
rlabel alu1 116 32 116 32 6 a2
rlabel alu1 132 36 132 36 6 a1
rlabel alu1 116 48 116 48 6 a1
rlabel alu1 124 48 124 48 6 a1
<< end >>
