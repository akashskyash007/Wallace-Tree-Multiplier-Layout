magic
tech scmos
timestamp 1199203404
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 28 66 30 71
rect 38 70 40 74
rect 45 70 47 74
rect 55 70 57 74
rect 65 70 67 74
rect 9 58 11 63
rect 9 39 11 42
rect 28 39 30 50
rect 38 44 40 50
rect 9 37 30 39
rect 34 42 40 44
rect 34 40 36 42
rect 38 40 40 42
rect 34 38 40 40
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 25 30 27 37
rect 35 30 37 38
rect 45 30 47 50
rect 55 47 57 50
rect 55 45 61 47
rect 55 43 57 45
rect 59 43 61 45
rect 55 41 61 43
rect 55 30 57 41
rect 65 39 67 50
rect 65 37 71 39
rect 65 35 67 37
rect 69 35 71 37
rect 62 33 71 35
rect 62 30 64 33
rect 9 26 15 28
rect 9 24 11 26
rect 13 24 15 26
rect 9 22 15 24
rect 13 11 15 22
rect 25 15 27 20
rect 35 15 37 20
rect 45 11 47 20
rect 55 15 57 20
rect 62 15 64 20
rect 13 9 47 11
<< ndif >>
rect 17 20 25 30
rect 27 26 35 30
rect 27 24 30 26
rect 32 24 35 26
rect 27 20 35 24
rect 37 28 45 30
rect 37 26 40 28
rect 42 26 45 28
rect 37 20 45 26
rect 47 28 55 30
rect 47 26 50 28
rect 52 26 55 28
rect 47 20 55 26
rect 57 20 62 30
rect 64 20 73 30
rect 17 19 23 20
rect 17 17 19 19
rect 21 17 23 19
rect 17 15 23 17
rect 66 19 73 20
rect 66 17 68 19
rect 70 17 73 19
rect 66 15 73 17
<< pdif >>
rect 33 66 38 70
rect 23 63 28 66
rect 21 61 28 63
rect 21 59 23 61
rect 25 59 28 61
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 48 9 54
rect 2 46 4 48
rect 6 46 9 48
rect 2 42 9 46
rect 11 48 16 58
rect 21 57 28 59
rect 23 50 28 57
rect 30 54 38 66
rect 30 52 33 54
rect 35 52 38 54
rect 30 50 38 52
rect 40 50 45 70
rect 47 68 55 70
rect 47 66 50 68
rect 52 66 55 68
rect 47 50 55 66
rect 57 61 65 70
rect 57 59 60 61
rect 62 59 65 61
rect 57 50 65 59
rect 67 68 74 70
rect 67 66 70 68
rect 72 66 74 68
rect 67 61 74 66
rect 67 59 70 61
rect 72 59 74 61
rect 67 50 74 59
rect 11 46 18 48
rect 11 44 14 46
rect 16 44 18 46
rect 11 42 18 44
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 26 54 38 55
rect 26 52 33 54
rect 35 52 38 54
rect 26 49 38 52
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 2 17 6 33
rect 26 31 30 49
rect 50 49 62 55
rect 56 45 62 49
rect 56 43 57 45
rect 59 43 62 45
rect 56 41 62 43
rect 66 37 70 39
rect 66 35 67 37
rect 69 35 70 37
rect 66 31 70 35
rect 58 25 70 31
rect -2 1 82 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 25 20 27 30
rect 35 20 37 30
rect 45 20 47 30
rect 55 20 57 30
rect 62 20 64 30
<< pmos >>
rect 9 42 11 58
rect 28 50 30 66
rect 38 50 40 70
rect 45 50 47 70
rect 55 50 57 70
rect 65 50 67 70
<< polyct0 >>
rect 36 40 38 42
rect 11 24 13 26
<< polyct1 >>
rect 11 35 13 37
rect 57 43 59 45
rect 67 35 69 37
<< ndifct0 >>
rect 30 24 32 26
rect 40 26 42 28
rect 50 26 52 28
rect 19 17 21 19
rect 68 17 70 19
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 23 59 25 61
rect 4 54 6 56
rect 4 46 6 48
rect 50 66 52 68
rect 60 59 62 61
rect 70 66 72 68
rect 70 59 72 61
rect 14 44 16 46
<< pdifct1 >>
rect 33 52 35 54
<< alu0 >>
rect 3 56 7 68
rect 48 66 50 68
rect 52 66 54 68
rect 48 65 54 66
rect 68 66 70 68
rect 72 66 74 68
rect 21 61 64 62
rect 21 59 23 61
rect 25 59 60 61
rect 62 59 64 61
rect 21 58 64 59
rect 68 61 74 66
rect 68 59 70 61
rect 72 59 74 61
rect 68 58 74 59
rect 3 54 4 56
rect 6 54 7 56
rect 3 48 7 54
rect 3 46 4 48
rect 6 46 7 48
rect 3 44 7 46
rect 12 46 22 47
rect 12 44 14 46
rect 16 44 22 46
rect 12 43 22 44
rect 18 27 22 43
rect 42 43 46 58
rect 34 42 51 43
rect 34 40 36 42
rect 38 40 51 42
rect 34 39 51 40
rect 30 31 41 35
rect 37 29 41 31
rect 47 29 51 39
rect 37 28 44 29
rect 9 26 34 27
rect 9 24 11 26
rect 13 24 30 26
rect 32 24 34 26
rect 37 26 40 28
rect 42 26 44 28
rect 37 25 44 26
rect 47 28 54 29
rect 47 26 50 28
rect 52 26 54 28
rect 47 25 54 26
rect 9 23 34 24
rect 17 19 23 20
rect 17 17 19 19
rect 21 17 23 19
rect 17 12 23 17
rect 67 19 71 21
rect 67 17 68 19
rect 70 17 71 19
rect 67 12 71 17
<< labels >>
rlabel alu0 21 25 21 25 6 bn
rlabel alu0 17 45 17 45 6 bn
rlabel alu0 49 34 49 34 6 an
rlabel alu0 42 41 42 41 6 an
rlabel alu0 42 60 42 60 6 an
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 28 4 28 6 b
rlabel alu1 28 44 28 44 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 52 52 52 52 6 a2
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 28 60 28 6 a1
rlabel alu1 68 32 68 32 6 a1
rlabel alu1 60 48 60 48 6 a2
<< end >>
