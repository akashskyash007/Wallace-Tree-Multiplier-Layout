magic
tech scmos
timestamp 1199203289
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 60 11 65
rect 22 55 24 60
rect 29 55 31 60
rect 36 55 38 60
rect 9 31 11 48
rect 22 42 24 45
rect 17 40 24 42
rect 17 38 19 40
rect 21 38 24 40
rect 17 36 24 38
rect 9 29 15 31
rect 9 27 11 29
rect 13 27 15 29
rect 9 25 15 27
rect 9 21 11 25
rect 19 21 21 36
rect 29 35 31 45
rect 36 42 38 45
rect 36 40 43 42
rect 29 33 35 35
rect 29 31 31 33
rect 33 31 35 33
rect 29 29 35 31
rect 29 21 31 29
rect 41 27 43 40
rect 41 25 47 27
rect 41 23 43 25
rect 45 23 47 25
rect 41 21 47 23
rect 41 18 43 21
rect 9 10 11 15
rect 19 11 21 15
rect 29 11 31 15
rect 41 7 43 12
<< ndif >>
rect 2 19 9 21
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 19 19 21
rect 11 17 14 19
rect 16 17 19 19
rect 11 15 19 17
rect 21 19 29 21
rect 21 17 24 19
rect 26 17 29 19
rect 21 15 29 17
rect 31 18 39 21
rect 31 15 41 18
rect 33 12 41 15
rect 43 16 50 18
rect 43 14 46 16
rect 48 14 50 16
rect 43 12 50 14
rect 33 7 39 12
rect 33 5 35 7
rect 37 5 39 7
rect 33 3 39 5
<< pdif >>
rect 13 67 20 69
rect 13 65 15 67
rect 17 65 20 67
rect 13 60 20 65
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 54 9 56
rect 4 48 9 54
rect 11 55 20 60
rect 11 48 22 55
rect 13 45 22 48
rect 24 45 29 55
rect 31 45 36 55
rect 38 51 43 55
rect 38 49 45 51
rect 38 47 41 49
rect 43 47 45 49
rect 38 45 45 47
<< alu1 >>
rect -2 67 58 72
rect -2 65 15 67
rect 17 65 26 67
rect 28 65 45 67
rect 47 65 58 67
rect -2 64 58 65
rect 2 58 15 59
rect 2 56 4 58
rect 6 56 15 58
rect 2 54 15 56
rect 2 19 6 54
rect 17 40 31 42
rect 17 38 19 40
rect 21 38 31 40
rect 17 30 23 38
rect 41 34 47 42
rect 29 33 47 34
rect 29 31 31 33
rect 33 31 47 33
rect 29 30 47 31
rect 2 17 4 19
rect 2 13 6 17
rect 33 25 47 26
rect 33 23 43 25
rect 45 23 47 25
rect 33 22 47 23
rect -2 7 58 8
rect -2 5 15 7
rect 17 5 25 7
rect 27 5 35 7
rect 37 5 58 7
rect -2 0 58 5
<< ptie >>
rect 13 7 29 9
rect 13 5 15 7
rect 17 5 25 7
rect 27 5 29 7
rect 13 3 29 5
<< ntie >>
rect 24 67 49 69
rect 24 65 26 67
rect 28 65 45 67
rect 47 65 49 67
rect 24 63 49 65
<< nmos >>
rect 9 15 11 21
rect 19 15 21 21
rect 29 15 31 21
rect 41 12 43 18
<< pmos >>
rect 9 48 11 60
rect 22 45 24 55
rect 29 45 31 55
rect 36 45 38 55
<< polyct0 >>
rect 11 27 13 29
<< polyct1 >>
rect 19 38 21 40
rect 31 31 33 33
rect 43 23 45 25
<< ndifct0 >>
rect 14 17 16 19
rect 24 17 26 19
rect 46 14 48 16
<< ndifct1 >>
rect 4 17 6 19
rect 35 5 37 7
<< ntiect1 >>
rect 26 65 28 67
rect 45 65 47 67
<< ptiect1 >>
rect 15 5 17 7
rect 25 5 27 7
<< pdifct0 >>
rect 41 47 43 49
<< pdifct1 >>
rect 15 65 17 67
rect 4 56 6 58
<< alu0 >>
rect 10 49 45 50
rect 10 47 41 49
rect 43 47 45 49
rect 10 46 45 47
rect 10 29 14 46
rect 10 27 11 29
rect 13 27 14 29
rect 10 23 27 27
rect 6 15 7 21
rect 12 19 18 20
rect 12 17 14 19
rect 16 17 18 19
rect 12 8 18 17
rect 23 19 27 23
rect 23 17 24 19
rect 26 17 27 19
rect 23 16 50 17
rect 23 14 46 16
rect 48 14 50 16
rect 23 13 50 14
<< labels >>
rlabel alu0 12 36 12 36 6 zn
rlabel alu0 25 20 25 20 6 zn
rlabel alu0 36 15 36 15 6 zn
rlabel alu0 27 48 27 48 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 36 20 36 6 a
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 24 36 24 6 c
rlabel alu1 36 32 36 32 6 b
rlabel alu1 28 40 28 40 6 a
rlabel alu1 28 68 28 68 6 vdd
rlabel polyct1 44 24 44 24 6 c
rlabel alu1 44 36 44 36 6 b
<< end >>
