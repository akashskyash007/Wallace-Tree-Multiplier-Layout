magic
tech scmos
timestamp 1199202314
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 9 59 11 63
rect 19 57 21 61
rect 9 35 11 38
rect 19 35 21 38
rect 9 33 21 35
rect 9 31 16 33
rect 18 31 21 33
rect 9 29 21 31
rect 9 26 11 29
rect 19 26 21 29
rect 9 2 11 6
rect 19 2 21 6
<< ndif >>
rect 2 17 9 26
rect 2 15 4 17
rect 6 15 9 17
rect 2 10 9 15
rect 2 8 4 10
rect 6 8 9 10
rect 2 6 9 8
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 11 15 14 17
rect 16 15 19 17
rect 11 6 19 15
rect 21 17 28 26
rect 21 15 24 17
rect 26 15 28 17
rect 21 10 28 15
rect 21 8 24 10
rect 26 8 28 10
rect 21 6 28 8
<< pdif >>
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 16 59
rect 11 55 19 57
rect 11 53 14 55
rect 16 53 19 55
rect 11 48 19 53
rect 11 46 14 48
rect 16 46 19 48
rect 11 38 19 46
rect 21 55 28 57
rect 21 53 24 55
rect 26 53 28 55
rect 21 48 28 53
rect 21 46 24 48
rect 26 46 28 48
rect 21 38 28 46
<< alu1 >>
rect -2 67 34 72
rect -2 65 22 67
rect 24 65 34 67
rect -2 64 34 65
rect 12 55 18 56
rect 12 53 14 55
rect 16 53 18 55
rect 12 51 18 53
rect 2 48 18 51
rect 2 46 14 48
rect 16 46 18 48
rect 2 25 6 46
rect 17 35 23 42
rect 10 33 23 35
rect 10 31 16 33
rect 18 31 23 33
rect 10 29 23 31
rect 2 24 18 25
rect 2 22 14 24
rect 16 22 18 24
rect 2 21 18 22
rect 13 17 18 21
rect 13 15 14 17
rect 16 15 18 17
rect 13 13 18 15
rect -2 0 34 8
<< ntie >>
rect 17 67 29 69
rect 17 65 22 67
rect 24 65 29 67
rect 17 63 29 65
<< nmos >>
rect 9 6 11 26
rect 19 6 21 26
<< pmos >>
rect 9 38 11 59
rect 19 38 21 57
<< polyct1 >>
rect 16 31 18 33
<< ndifct0 >>
rect 4 15 6 17
rect 4 8 6 10
rect 24 15 26 17
rect 24 8 26 10
<< ndifct1 >>
rect 14 22 16 24
rect 14 15 16 17
<< ntiect1 >>
rect 22 65 24 67
<< pdifct0 >>
rect 4 55 6 57
rect 24 53 26 55
rect 24 46 26 48
<< pdifct1 >>
rect 14 53 16 55
rect 14 46 16 48
<< alu0 >>
rect 2 57 8 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 6 45 18 46
rect 22 55 28 64
rect 22 53 24 55
rect 26 53 28 55
rect 22 48 28 53
rect 22 46 24 48
rect 26 46 28 48
rect 22 45 28 46
rect 2 17 8 18
rect 2 15 4 17
rect 6 15 8 17
rect 2 10 8 15
rect 22 17 28 18
rect 22 15 24 17
rect 26 15 28 17
rect 2 8 4 10
rect 6 8 8 10
rect 22 10 28 15
rect 22 8 24 10
rect 26 8 28 10
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 32 12 32 6 a
rlabel alu1 12 48 12 48 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 16 68 16 68 6 vdd
<< end >>
