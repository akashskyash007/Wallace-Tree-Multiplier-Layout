magic
tech scmos
timestamp 1199203692
<< ab >>
rect 0 0 168 72
<< nwell >>
rect -5 32 173 77
<< pwell >>
rect -5 -5 173 32
<< poly >>
rect 11 66 13 70
rect 19 66 21 70
rect 27 66 29 70
rect 37 66 39 70
rect 44 66 46 70
rect 54 66 56 70
rect 75 66 77 70
rect 104 66 106 70
rect 114 66 116 70
rect 121 66 123 70
rect 131 66 133 70
rect 139 66 141 70
rect 147 66 149 70
rect 86 42 92 44
rect 86 40 88 42
rect 90 40 92 42
rect 86 38 92 40
rect 159 43 165 45
rect 159 41 161 43
rect 163 41 165 43
rect 159 39 165 41
rect 11 35 13 38
rect 19 35 21 38
rect 27 35 29 38
rect 37 35 39 38
rect 44 35 46 38
rect 54 35 56 38
rect 75 35 77 38
rect 86 35 88 38
rect 2 33 13 35
rect 2 31 4 33
rect 6 31 13 33
rect 2 29 13 31
rect 17 33 23 35
rect 17 31 19 33
rect 21 31 23 33
rect 17 29 23 31
rect 27 33 40 35
rect 27 31 36 33
rect 38 31 40 33
rect 44 32 48 35
rect 54 32 58 35
rect 27 29 40 31
rect 11 26 13 29
rect 19 26 21 29
rect 27 26 29 29
rect 37 26 39 29
rect 46 28 48 32
rect 46 26 52 28
rect 46 24 48 26
rect 50 24 52 26
rect 46 22 52 24
rect 46 19 48 22
rect 56 19 58 32
rect 62 33 77 35
rect 62 31 64 33
rect 66 31 77 33
rect 62 29 77 31
rect 83 33 88 35
rect 104 34 106 38
rect 68 26 70 29
rect 11 7 13 12
rect 19 7 21 12
rect 27 7 29 12
rect 37 7 39 12
rect 83 18 85 33
rect 92 32 106 34
rect 92 30 94 32
rect 96 30 106 32
rect 92 28 106 30
rect 104 25 106 28
rect 114 25 116 38
rect 121 35 123 38
rect 131 35 133 38
rect 139 35 141 38
rect 147 35 149 38
rect 159 35 161 39
rect 121 33 133 35
rect 121 31 123 33
rect 125 31 133 33
rect 121 29 133 31
rect 137 33 143 35
rect 137 31 139 33
rect 141 31 143 33
rect 137 29 143 31
rect 147 33 161 35
rect 121 25 123 29
rect 131 25 133 29
rect 139 25 141 29
rect 147 25 149 33
rect 79 16 85 18
rect 79 14 81 16
rect 83 14 85 16
rect 79 12 85 14
rect 68 8 70 12
rect 160 17 166 19
rect 160 15 162 17
rect 164 15 166 17
rect 160 13 166 15
rect 104 8 106 12
rect 46 2 48 7
rect 56 4 58 7
rect 114 4 116 12
rect 121 8 123 12
rect 131 8 133 12
rect 139 8 141 12
rect 147 8 149 12
rect 160 4 162 13
rect 56 2 162 4
<< ndif >>
rect 3 12 11 26
rect 13 12 19 26
rect 21 12 27 26
rect 29 24 37 26
rect 29 22 32 24
rect 34 22 37 24
rect 29 12 37 22
rect 39 19 44 26
rect 60 19 68 26
rect 39 12 46 19
rect 3 7 9 12
rect 41 7 46 12
rect 48 16 56 19
rect 48 14 51 16
rect 53 14 56 16
rect 48 7 56 14
rect 58 18 68 19
rect 58 16 62 18
rect 64 16 68 18
rect 58 12 68 16
rect 70 18 75 26
rect 70 16 77 18
rect 70 14 73 16
rect 75 14 77 16
rect 70 12 77 14
rect 58 11 66 12
rect 58 9 62 11
rect 64 9 66 11
rect 58 7 66 9
rect 97 16 104 25
rect 97 14 99 16
rect 101 14 104 16
rect 97 12 104 14
rect 106 23 114 25
rect 106 21 109 23
rect 111 21 114 23
rect 106 16 114 21
rect 106 14 109 16
rect 111 14 114 16
rect 106 12 114 14
rect 116 12 121 25
rect 123 17 131 25
rect 123 15 126 17
rect 128 15 131 17
rect 123 12 131 15
rect 133 12 139 25
rect 141 12 147 25
rect 149 23 158 25
rect 149 21 154 23
rect 156 21 158 23
rect 149 16 158 21
rect 149 14 154 16
rect 156 14 158 16
rect 149 12 158 14
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< pdif >>
rect 3 64 11 66
rect 3 62 6 64
rect 8 62 11 64
rect 3 38 11 62
rect 13 38 19 66
rect 21 38 27 66
rect 29 49 37 66
rect 29 47 32 49
rect 34 47 37 49
rect 29 38 37 47
rect 39 38 44 66
rect 46 57 54 66
rect 46 55 49 57
rect 51 55 54 57
rect 46 38 54 55
rect 56 64 75 66
rect 56 62 60 64
rect 62 62 70 64
rect 72 62 75 64
rect 56 38 75 62
rect 77 44 82 66
rect 97 64 104 66
rect 97 62 99 64
rect 101 62 104 64
rect 77 42 84 44
rect 77 40 80 42
rect 82 40 84 42
rect 77 38 84 40
rect 97 38 104 62
rect 106 42 114 66
rect 106 40 109 42
rect 111 40 114 42
rect 106 38 114 40
rect 116 38 121 66
rect 123 49 131 66
rect 123 47 126 49
rect 128 47 131 49
rect 123 38 131 47
rect 133 38 139 66
rect 141 38 147 66
rect 149 59 155 66
rect 149 57 157 59
rect 149 55 152 57
rect 154 55 157 57
rect 149 38 157 55
<< alu1 >>
rect -2 67 170 72
rect -2 65 88 67
rect 90 65 161 67
rect 163 65 170 67
rect -2 64 170 65
rect 10 49 141 50
rect 10 47 32 49
rect 34 47 126 49
rect 128 47 141 49
rect 10 46 141 47
rect 10 25 14 46
rect 25 38 73 42
rect 25 35 30 38
rect 18 33 30 35
rect 137 42 141 46
rect 137 38 150 42
rect 18 31 19 33
rect 21 31 30 33
rect 18 29 30 31
rect 34 33 68 34
rect 34 31 36 33
rect 38 31 64 33
rect 66 31 68 33
rect 34 30 68 31
rect 73 32 97 34
rect 73 30 94 32
rect 96 30 97 32
rect 93 28 97 30
rect 10 24 36 25
rect 10 22 32 24
rect 34 22 36 24
rect 10 21 36 22
rect 146 18 150 38
rect 154 29 166 35
rect 124 17 150 18
rect 124 15 126 17
rect 128 15 150 17
rect 124 14 150 15
rect 161 17 166 29
rect 161 15 162 17
rect 164 15 166 17
rect 161 13 166 15
rect -2 7 170 8
rect -2 5 5 7
rect 7 5 170 7
rect -2 0 170 5
<< ptie >>
rect 87 10 93 24
rect 87 8 89 10
rect 91 8 93 10
rect 87 6 93 8
<< ntie >>
rect 86 67 92 69
rect 86 65 88 67
rect 90 65 92 67
rect 159 67 165 69
rect 86 48 92 65
rect 159 65 161 67
rect 163 65 165 67
rect 159 63 165 65
<< nmos >>
rect 11 12 13 26
rect 19 12 21 26
rect 27 12 29 26
rect 37 12 39 26
rect 46 7 48 19
rect 56 7 58 19
rect 68 12 70 26
rect 104 12 106 25
rect 114 12 116 25
rect 121 12 123 25
rect 131 12 133 25
rect 139 12 141 25
rect 147 12 149 25
<< pmos >>
rect 11 38 13 66
rect 19 38 21 66
rect 27 38 29 66
rect 37 38 39 66
rect 44 38 46 66
rect 54 38 56 66
rect 75 38 77 66
rect 104 38 106 66
rect 114 38 116 66
rect 121 38 123 66
rect 131 38 133 66
rect 139 38 141 66
rect 147 38 149 66
<< polyct0 >>
rect 88 40 90 42
rect 161 41 163 43
rect 4 31 6 33
rect 48 24 50 26
rect 123 31 125 33
rect 139 31 141 33
rect 81 14 83 16
<< polyct1 >>
rect 19 31 21 33
rect 36 31 38 33
rect 64 31 66 33
rect 94 30 96 32
rect 162 15 164 17
<< ndifct0 >>
rect 51 14 53 16
rect 62 16 64 18
rect 73 14 75 16
rect 62 9 64 11
rect 99 14 101 16
rect 109 21 111 23
rect 109 14 111 16
rect 154 21 156 23
rect 154 14 156 16
<< ndifct1 >>
rect 32 22 34 24
rect 126 15 128 17
rect 5 5 7 7
<< ntiect1 >>
rect 88 65 90 67
rect 161 65 163 67
<< ptiect0 >>
rect 89 8 91 10
<< pdifct0 >>
rect 6 62 8 64
rect 49 55 51 57
rect 60 62 62 64
rect 70 62 72 64
rect 99 62 101 64
rect 80 40 82 42
rect 109 40 111 42
rect 152 55 154 57
<< pdifct1 >>
rect 32 47 34 49
rect 126 47 128 49
<< alu0 >>
rect 4 62 6 64
rect 8 62 10 64
rect 4 61 10 62
rect 58 62 60 64
rect 62 62 70 64
rect 72 62 74 64
rect 58 61 74 62
rect 97 62 99 64
rect 101 62 103 64
rect 97 61 103 62
rect 3 57 148 58
rect 3 55 49 57
rect 51 55 148 57
rect 3 54 148 55
rect 3 33 7 54
rect 144 50 148 54
rect 151 57 155 64
rect 151 55 152 57
rect 154 55 155 57
rect 151 53 155 55
rect 3 31 4 33
rect 6 31 7 33
rect 3 17 7 31
rect 144 46 164 50
rect 78 42 104 43
rect 73 38 75 42
rect 78 40 80 42
rect 82 40 88 42
rect 90 40 104 42
rect 78 39 104 40
rect 71 34 75 38
rect 100 34 104 39
rect 107 42 113 43
rect 160 43 164 46
rect 107 40 109 42
rect 111 40 134 42
rect 107 38 134 40
rect 160 41 161 43
rect 163 41 164 43
rect 160 39 164 41
rect 130 34 134 38
rect 71 30 73 34
rect 100 33 127 34
rect 100 31 123 33
rect 125 31 127 33
rect 100 30 127 31
rect 130 33 143 34
rect 130 31 139 33
rect 141 31 143 33
rect 130 30 143 31
rect 46 26 52 27
rect 130 26 134 30
rect 46 24 48 26
rect 50 25 89 26
rect 107 25 134 26
rect 50 24 134 25
rect 46 23 134 24
rect 46 22 109 23
rect 85 21 109 22
rect 111 22 134 23
rect 111 21 113 22
rect 60 18 66 19
rect 3 16 55 17
rect 3 14 51 16
rect 53 14 55 16
rect 3 13 55 14
rect 60 16 62 18
rect 64 16 66 18
rect 60 11 66 16
rect 71 16 85 17
rect 71 14 73 16
rect 75 14 81 16
rect 83 14 85 16
rect 71 13 85 14
rect 97 16 103 17
rect 97 14 99 16
rect 101 14 103 16
rect 60 9 62 11
rect 64 9 66 11
rect 60 8 66 9
rect 88 10 92 12
rect 88 8 89 10
rect 91 8 92 10
rect 97 8 103 14
rect 107 16 113 21
rect 107 14 109 16
rect 111 14 113 16
rect 153 23 157 25
rect 153 21 154 23
rect 156 21 157 23
rect 153 16 157 21
rect 153 14 154 16
rect 156 14 157 16
rect 107 13 113 14
rect 153 8 157 14
<< labels >>
rlabel alu0 5 35 5 35 6 an
rlabel alu0 29 15 29 15 6 an
rlabel alu0 78 15 78 15 6 cn
rlabel alu0 110 19 110 19 6 bn
rlabel alu0 67 24 67 24 6 bn
rlabel alu0 91 41 91 41 6 cn
rlabel alu0 113 32 113 32 6 cn
rlabel alu0 136 32 136 32 6 bn
rlabel alu0 120 40 120 40 6 bn
rlabel alu0 162 44 162 44 6 an
rlabel alu0 75 56 75 56 6 an
rlabel alu1 12 32 12 32 6 z
rlabel polyct1 20 32 20 32 6 b
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 44 32 44 32 6 c
rlabel alu1 52 32 52 32 6 c
rlabel alu1 60 32 60 32 6 c
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 52 40 52 40 6 b
rlabel alu1 60 40 60 40 6 b
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 84 4 84 4 6 vss
rlabel alu1 76 32 76 32 6 b
rlabel alu1 84 32 84 32 6 b
rlabel alu1 92 32 92 32 6 b
rlabel alu1 68 40 68 40 6 b
rlabel alu1 68 48 68 48 6 z
rlabel alu1 76 48 76 48 6 z
rlabel alu1 84 48 84 48 6 z
rlabel alu1 92 48 92 48 6 z
rlabel alu1 84 68 84 68 6 vdd
rlabel alu1 132 16 132 16 6 z
rlabel alu1 100 48 100 48 6 z
rlabel alu1 108 48 108 48 6 z
rlabel alu1 116 48 116 48 6 z
rlabel alu1 124 48 124 48 6 z
rlabel alu1 132 48 132 48 6 z
rlabel alu1 140 16 140 16 6 z
rlabel alu1 164 24 164 24 6 a
rlabel alu1 148 28 148 28 6 z
rlabel alu1 156 32 156 32 6 a
rlabel alu1 140 40 140 40 6 z
<< end >>
