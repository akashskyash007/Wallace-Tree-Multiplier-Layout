magic
tech scmos
timestamp 1199202224
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 70 11 74
rect 32 67 34 72
rect 39 67 41 72
rect 57 70 59 74
rect 67 70 69 74
rect 77 70 79 74
rect 22 58 24 63
rect 9 32 11 45
rect 22 42 24 45
rect 15 40 24 42
rect 15 38 17 40
rect 19 38 21 40
rect 32 39 34 42
rect 39 39 41 42
rect 57 39 59 42
rect 67 39 69 42
rect 77 39 79 42
rect 15 36 21 38
rect 9 30 15 32
rect 9 28 11 30
rect 13 28 15 30
rect 9 26 15 28
rect 9 23 11 26
rect 19 23 21 36
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 39 37 61 39
rect 39 35 50 37
rect 52 35 57 37
rect 59 35 61 37
rect 39 33 61 35
rect 65 37 71 39
rect 65 35 67 37
rect 69 35 71 37
rect 65 33 71 35
rect 75 37 81 39
rect 75 35 77 37
rect 79 35 81 37
rect 75 33 81 35
rect 29 30 31 33
rect 39 30 41 33
rect 59 30 61 33
rect 66 30 68 33
rect 9 6 11 10
rect 19 8 21 13
rect 29 11 31 16
rect 39 11 41 16
rect 77 24 79 33
rect 59 6 61 10
rect 66 6 68 10
rect 77 6 79 10
<< ndif >>
rect 24 23 29 30
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 17 19 23
rect 11 15 14 17
rect 16 15 19 17
rect 11 13 19 15
rect 21 20 29 23
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 16 39 26
rect 41 28 48 30
rect 41 26 44 28
rect 46 26 48 28
rect 41 21 48 26
rect 54 23 59 30
rect 41 19 44 21
rect 46 19 48 21
rect 41 16 48 19
rect 52 21 59 23
rect 52 19 54 21
rect 56 19 59 21
rect 52 17 59 19
rect 21 13 26 16
rect 11 10 16 13
rect 54 10 59 17
rect 61 10 66 30
rect 68 24 75 30
rect 68 14 77 24
rect 68 12 71 14
rect 73 12 77 14
rect 68 10 77 12
rect 79 21 86 24
rect 79 19 82 21
rect 84 19 86 21
rect 79 17 86 19
rect 79 10 84 17
<< pdif >>
rect 4 58 9 70
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 11 68 20 70
rect 11 66 15 68
rect 17 66 20 68
rect 43 68 57 70
rect 43 67 50 68
rect 11 58 20 66
rect 27 58 32 67
rect 11 45 22 58
rect 24 49 32 58
rect 24 47 27 49
rect 29 47 32 49
rect 24 45 32 47
rect 27 42 32 45
rect 34 42 39 67
rect 41 66 50 67
rect 52 66 57 68
rect 41 61 57 66
rect 41 59 50 61
rect 52 59 57 61
rect 41 42 57 59
rect 59 60 67 70
rect 59 58 62 60
rect 64 58 67 60
rect 59 53 67 58
rect 59 51 62 53
rect 64 51 67 53
rect 59 42 67 51
rect 69 68 77 70
rect 69 66 72 68
rect 74 66 77 68
rect 69 61 77 66
rect 69 59 72 61
rect 74 59 77 61
rect 69 42 77 59
rect 79 55 84 70
rect 79 53 86 55
rect 79 51 82 53
rect 84 51 86 53
rect 79 46 86 51
rect 79 44 82 46
rect 84 44 86 46
rect 79 42 86 44
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 2 58 15 62
rect 2 56 7 58
rect 2 54 4 56
rect 6 54 7 56
rect 2 49 7 54
rect 2 47 4 49
rect 6 47 7 49
rect 2 45 7 47
rect 2 23 6 45
rect 33 42 71 46
rect 33 39 38 42
rect 30 37 38 39
rect 30 35 31 37
rect 33 35 38 37
rect 30 33 38 35
rect 48 37 63 38
rect 48 35 50 37
rect 52 35 57 37
rect 59 35 63 37
rect 48 34 63 35
rect 2 21 7 23
rect 50 25 54 34
rect 81 53 87 55
rect 81 51 82 53
rect 84 51 87 53
rect 81 46 87 51
rect 81 44 82 46
rect 84 44 87 46
rect 81 42 87 44
rect 83 22 87 42
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect 65 21 87 22
rect 65 19 82 21
rect 84 19 87 21
rect 65 18 87 19
rect -2 1 98 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 9 10 11 23
rect 19 13 21 23
rect 29 16 31 30
rect 39 16 41 30
rect 59 10 61 30
rect 66 10 68 30
rect 77 10 79 24
<< pmos >>
rect 9 45 11 70
rect 22 45 24 58
rect 32 42 34 67
rect 39 42 41 67
rect 57 42 59 70
rect 67 42 69 70
rect 77 42 79 70
<< polyct0 >>
rect 17 38 19 40
rect 11 28 13 30
rect 67 35 69 37
rect 77 35 79 37
<< polyct1 >>
rect 31 35 33 37
rect 50 35 52 37
rect 57 35 59 37
<< ndifct0 >>
rect 14 15 16 17
rect 24 18 26 20
rect 34 26 36 28
rect 44 26 46 28
rect 44 19 46 21
rect 54 19 56 21
rect 71 12 73 14
<< ndifct1 >>
rect 4 19 6 21
rect 82 19 84 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 15 66 17 68
rect 27 47 29 49
rect 50 66 52 68
rect 50 59 52 61
rect 62 58 64 60
rect 62 51 64 53
rect 72 66 74 68
rect 72 59 74 61
<< pdifct1 >>
rect 4 54 6 56
rect 4 47 6 49
rect 82 51 84 53
rect 82 44 84 46
<< alu0 >>
rect 13 66 15 68
rect 17 66 19 68
rect 13 65 19 66
rect 48 66 50 68
rect 52 66 54 68
rect 48 61 54 66
rect 70 66 72 68
rect 74 66 76 68
rect 48 59 50 61
rect 52 59 54 61
rect 48 58 54 59
rect 61 60 65 62
rect 61 58 62 60
rect 64 58 65 60
rect 70 61 76 66
rect 70 59 72 61
rect 74 59 76 61
rect 70 58 76 59
rect 18 54 42 58
rect 61 54 65 58
rect 16 50 22 54
rect 38 53 78 54
rect 38 51 62 53
rect 64 51 78 53
rect 16 40 20 50
rect 26 49 30 51
rect 38 50 78 51
rect 26 47 27 49
rect 29 47 30 49
rect 26 46 30 47
rect 16 38 17 40
rect 19 38 20 40
rect 16 36 20 38
rect 23 42 30 46
rect 23 31 27 42
rect 66 37 70 42
rect 66 35 67 37
rect 69 35 70 37
rect 9 30 27 31
rect 9 28 11 30
rect 13 29 27 30
rect 13 28 38 29
rect 9 27 34 28
rect 23 26 34 27
rect 36 26 38 28
rect 23 25 38 26
rect 43 28 47 30
rect 43 26 44 28
rect 46 26 47 28
rect 43 21 47 26
rect 66 33 70 35
rect 74 39 78 50
rect 74 37 80 39
rect 74 35 77 37
rect 79 35 80 37
rect 74 33 80 35
rect 74 30 78 33
rect 58 26 78 30
rect 58 22 62 26
rect 22 20 44 21
rect 13 17 17 19
rect 22 18 24 20
rect 26 19 44 20
rect 46 19 47 21
rect 26 18 47 19
rect 52 21 62 22
rect 52 19 54 21
rect 56 19 62 21
rect 52 18 62 19
rect 22 17 47 18
rect 13 15 14 17
rect 16 15 17 17
rect 13 12 17 15
rect 69 14 75 15
rect 69 12 71 14
rect 73 12 75 14
<< labels >>
rlabel alu0 18 45 18 45 6 con
rlabel alu0 45 23 45 23 6 n2
rlabel alu0 34 19 34 19 6 n2
rlabel alu0 30 27 30 27 6 son
rlabel alu0 18 29 18 29 6 son
rlabel alu0 28 46 28 46 6 son
rlabel alu0 57 20 57 20 6 con
rlabel alu0 63 56 63 56 6 con
rlabel alu0 76 40 76 40 6 con
rlabel alu0 58 52 58 52 6 con
rlabel alu1 4 36 4 36 6 so
rlabel alu1 12 60 12 60 6 so
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 68 20 68 20 6 co
rlabel alu1 52 32 52 32 6 a
rlabel alu1 60 36 60 36 6 a
rlabel alu1 68 44 68 44 6 b
rlabel alu1 60 44 60 44 6 b
rlabel alu1 52 44 52 44 6 b
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 84 20 84 20 6 co
rlabel alu1 76 20 76 20 6 co
rlabel alu1 84 48 84 48 6 co
<< end >>
