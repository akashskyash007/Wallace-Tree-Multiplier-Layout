magic
tech scmos
timestamp 1199201816
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 64 11 69
rect 21 64 23 69
rect 61 66 63 71
rect 39 58 41 63
rect 49 58 51 63
rect 9 49 11 52
rect 9 47 15 49
rect 9 45 11 47
rect 13 45 15 47
rect 9 43 15 45
rect 9 22 11 43
rect 21 39 23 52
rect 61 47 63 50
rect 60 45 66 47
rect 60 43 62 45
rect 64 43 66 45
rect 39 39 41 42
rect 17 37 23 39
rect 17 35 19 37
rect 21 35 23 37
rect 17 33 23 35
rect 33 37 41 39
rect 33 35 35 37
rect 37 35 41 37
rect 49 39 51 42
rect 60 41 66 43
rect 49 37 55 39
rect 49 35 51 37
rect 53 35 55 37
rect 33 33 45 35
rect 49 33 55 35
rect 21 30 23 33
rect 43 30 45 33
rect 53 30 55 33
rect 60 30 62 41
rect 21 19 23 24
rect 9 11 11 16
rect 43 19 45 24
rect 53 18 55 23
rect 60 18 62 23
<< ndif >>
rect 13 24 21 30
rect 23 28 30 30
rect 23 26 26 28
rect 28 26 30 28
rect 23 24 30 26
rect 34 24 43 30
rect 45 28 53 30
rect 45 26 48 28
rect 50 26 53 28
rect 45 24 53 26
rect 13 22 19 24
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 19 22
rect 13 11 19 16
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
rect 34 11 41 24
rect 48 23 53 24
rect 55 23 60 30
rect 62 27 69 30
rect 62 25 65 27
rect 67 25 69 27
rect 62 23 69 25
rect 34 9 37 11
rect 39 9 41 11
rect 34 7 41 9
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 64 19 69
rect 53 64 61 66
rect 4 58 9 64
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 52 9 54
rect 11 52 21 64
rect 23 58 28 64
rect 53 62 55 64
rect 57 62 61 64
rect 53 58 61 62
rect 23 56 30 58
rect 23 54 26 56
rect 28 54 30 56
rect 23 52 30 54
rect 34 48 39 58
rect 32 46 39 48
rect 32 44 34 46
rect 36 44 39 46
rect 32 42 39 44
rect 41 54 49 58
rect 41 52 44 54
rect 46 52 49 54
rect 41 42 49 52
rect 51 50 61 58
rect 63 63 68 66
rect 63 61 70 63
rect 63 59 66 61
rect 68 59 70 61
rect 63 54 70 59
rect 63 52 66 54
rect 68 52 70 54
rect 63 50 70 52
rect 51 42 58 50
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 71 74 79
rect -2 69 15 71
rect 17 69 74 71
rect -2 68 74 69
rect 10 57 22 63
rect 10 47 14 57
rect 10 45 11 47
rect 13 45 14 47
rect 10 43 14 45
rect 18 39 22 47
rect 10 37 22 39
rect 10 35 19 37
rect 21 35 22 37
rect 10 33 22 35
rect 33 47 38 55
rect 33 46 46 47
rect 33 44 34 46
rect 36 44 46 46
rect 33 41 46 44
rect 57 45 70 47
rect 57 43 62 45
rect 64 43 70 45
rect 57 42 70 43
rect 10 25 14 33
rect 42 29 46 41
rect 42 28 52 29
rect 42 26 48 28
rect 50 26 52 28
rect 42 25 52 26
rect 66 33 70 42
rect -2 11 74 12
rect -2 9 15 11
rect 17 9 37 11
rect 39 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 21 24 23 30
rect 43 24 45 30
rect 9 16 11 22
rect 53 23 55 30
rect 60 23 62 30
<< pmos >>
rect 9 52 11 64
rect 21 52 23 64
rect 39 42 41 58
rect 49 42 51 58
rect 61 50 63 66
<< polyct0 >>
rect 35 35 37 37
rect 51 35 53 37
<< polyct1 >>
rect 11 45 13 47
rect 62 43 64 45
rect 19 35 21 37
<< ndifct0 >>
rect 26 26 28 28
rect 4 18 6 20
rect 65 25 67 27
<< ndifct1 >>
rect 48 26 50 28
rect 15 9 17 11
rect 37 9 39 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 54 6 56
rect 55 62 57 64
rect 26 54 28 56
rect 44 52 46 54
rect 66 59 68 61
rect 66 52 68 54
<< pdifct1 >>
rect 15 69 17 71
rect 34 44 36 46
<< alu0 >>
rect 54 64 58 68
rect 2 56 7 58
rect 2 54 4 56
rect 6 54 7 56
rect 2 52 7 54
rect 54 62 55 64
rect 57 62 58 64
rect 54 60 58 62
rect 64 61 70 62
rect 64 59 66 61
rect 68 59 70 61
rect 2 21 6 52
rect 25 56 29 58
rect 25 54 26 56
rect 28 54 29 56
rect 64 55 70 59
rect 25 38 29 54
rect 42 54 70 55
rect 42 52 44 54
rect 46 52 66 54
rect 68 52 70 54
rect 42 51 70 52
rect 25 37 39 38
rect 25 35 35 37
rect 37 35 39 37
rect 25 34 39 35
rect 25 28 29 34
rect 25 26 26 28
rect 28 26 29 28
rect 25 24 29 26
rect 49 37 60 38
rect 49 35 51 37
rect 53 35 60 37
rect 49 34 60 35
rect 56 21 60 34
rect 2 20 60 21
rect 2 18 4 20
rect 6 18 60 20
rect 2 17 60 18
rect 64 27 68 29
rect 64 25 65 27
rect 67 25 68 27
rect 64 12 68 25
<< labels >>
rlabel alu0 4 55 4 55 6 a2n
rlabel alu0 27 41 27 41 6 bn
rlabel alu0 32 36 32 36 6 bn
rlabel alu0 31 19 31 19 6 a2n
rlabel alu0 54 36 54 36 6 a2n
rlabel alu0 56 53 56 53 6 n1
rlabel alu0 67 56 67 56 6 n1
rlabel alu1 12 32 12 32 6 b
rlabel alu1 12 56 12 56 6 a2
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 60 20 60 6 a2
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 44 36 44 36 6 z
rlabel alu1 36 44 36 44 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 44 60 44 6 a1
rlabel alu1 68 40 68 40 6 a1
<< end >>
