magic
tech scmos
timestamp 1199980634
<< ab >>
rect 0 0 32 88
<< nwell >>
rect -8 40 40 97
<< pwell >>
rect -8 -9 40 40
<< poly >>
rect 5 80 14 86
rect 18 84 27 86
rect 18 82 23 84
rect 25 82 27 84
rect 18 80 27 82
rect 9 77 11 80
rect 21 77 23 80
rect 9 48 11 51
rect 21 48 23 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 42 30 48
rect 2 36 17 38
rect 2 34 7 36
rect 9 34 17 36
rect 2 32 17 34
rect 21 32 30 38
rect 9 29 11 32
rect 21 29 23 32
rect 9 8 11 11
rect 21 8 23 11
rect 5 2 14 8
rect 18 6 27 8
rect 18 4 23 6
rect 25 4 27 6
rect 18 2 27 4
<< ndif >>
rect 2 15 9 29
rect 2 13 4 15
rect 6 13 9 15
rect 2 11 9 13
rect 11 25 21 29
rect 11 23 15 25
rect 17 23 21 25
rect 11 17 21 23
rect 11 15 15 17
rect 17 15 21 17
rect 11 11 21 15
rect 23 11 30 29
<< pdif >>
rect 2 74 9 77
rect 2 72 4 74
rect 6 72 9 74
rect 2 67 9 72
rect 2 65 4 67
rect 6 65 9 67
rect 2 51 9 65
rect 11 65 21 77
rect 11 63 15 65
rect 17 63 21 65
rect 11 57 21 63
rect 11 55 15 57
rect 17 55 21 57
rect 11 51 21 55
rect 23 51 30 77
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 83 6 85
rect -2 81 6 83
rect 30 83 31 85
rect 33 83 34 85
rect 30 81 34 83
rect 2 76 6 81
rect 2 74 7 76
rect 2 72 4 74
rect 6 72 7 74
rect 2 67 7 72
rect 2 65 4 67
rect 6 65 7 67
rect 2 63 7 65
rect 14 65 18 67
rect 14 63 15 65
rect 17 63 18 65
rect 14 57 18 63
rect 14 55 15 57
rect 17 55 18 57
rect 6 46 10 48
rect 6 44 7 46
rect 9 44 10 46
rect 6 36 10 44
rect 6 34 7 36
rect 9 34 10 36
rect 6 21 10 34
rect 14 25 18 55
rect 14 23 15 25
rect 17 23 18 25
rect 14 17 18 23
rect 3 15 7 17
rect 3 13 4 15
rect 6 13 7 15
rect 14 15 15 17
rect 17 15 18 17
rect 14 13 18 15
rect 3 7 7 13
rect -2 5 7 7
rect -2 3 -1 5
rect 1 3 7 5
rect 30 5 34 7
rect 30 3 31 5
rect 33 3 34 5
rect -2 -2 2 3
rect 30 -2 34 3
<< alu2 >>
rect -2 85 34 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 80 34 83
rect -2 5 34 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 34 5
rect -2 -2 34 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
<< polyct0 >>
rect 23 82 25 84
rect 23 4 25 6
<< polyct1 >>
rect 7 44 9 46
rect 7 34 9 36
<< ndifct1 >>
rect 4 13 6 15
rect 15 23 17 25
rect 15 15 17 17
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
<< pdifct1 >>
rect 4 72 6 74
rect 4 65 6 67
rect 15 63 17 65
rect 15 55 17 57
<< alu0 >>
rect 21 84 30 85
rect 21 82 23 84
rect 25 82 30 84
rect 21 81 30 82
rect 21 6 30 7
rect 21 4 23 6
rect 25 4 30 6
rect 21 3 30 4
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect -1 3 1 5
rect 31 3 33 5
<< labels >>
rlabel alu1 8 32 8 32 6 a
rlabel alu1 16 40 16 40 6 z
rlabel alu2 16 4 16 4 6 vss
rlabel alu2 16 84 16 84 6 vdd
<< end >>
