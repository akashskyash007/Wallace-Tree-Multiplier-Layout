magic
tech scmos
timestamp 1199203106
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 12 66 14 70
rect 22 66 24 70
rect 29 66 31 70
rect 12 46 14 52
rect 9 44 15 46
rect 9 42 11 44
rect 13 42 15 44
rect 9 40 15 42
rect 9 18 11 40
rect 22 36 24 39
rect 17 34 24 36
rect 17 32 19 34
rect 21 32 24 34
rect 17 30 24 32
rect 29 35 31 39
rect 29 33 38 35
rect 29 31 34 33
rect 36 31 38 33
rect 19 18 21 30
rect 29 29 38 31
rect 29 18 31 29
rect 9 2 11 6
rect 19 2 21 6
rect 29 2 31 6
<< ndif >>
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 4 6 9 12
rect 11 16 19 18
rect 11 14 14 16
rect 16 14 19 16
rect 11 6 19 14
rect 21 10 29 18
rect 21 8 24 10
rect 26 8 29 10
rect 21 6 29 8
rect 31 16 38 18
rect 31 14 34 16
rect 36 14 38 16
rect 31 12 38 14
rect 31 6 36 12
<< pdif >>
rect 4 64 12 66
rect 4 62 7 64
rect 9 62 12 64
rect 4 52 12 62
rect 14 57 22 66
rect 14 55 17 57
rect 19 55 22 57
rect 14 52 22 55
rect 17 39 22 52
rect 24 39 29 66
rect 31 64 38 66
rect 31 62 34 64
rect 36 62 38 64
rect 31 57 38 62
rect 31 55 34 57
rect 36 55 38 57
rect 31 39 38 55
<< alu1 >>
rect -2 64 42 72
rect 2 57 23 58
rect 2 55 17 57
rect 19 55 23 57
rect 2 54 23 55
rect 2 18 6 54
rect 10 44 14 46
rect 10 42 11 44
rect 13 42 14 44
rect 25 43 31 50
rect 10 26 14 42
rect 18 38 31 43
rect 25 33 38 34
rect 25 31 34 33
rect 36 31 38 33
rect 25 30 38 31
rect 10 22 23 26
rect 34 21 38 30
rect 2 16 8 18
rect 2 14 4 16
rect 6 14 8 16
rect 2 13 8 14
rect -2 0 42 8
<< nmos >>
rect 9 6 11 18
rect 19 6 21 18
rect 29 6 31 18
<< pmos >>
rect 12 52 14 66
rect 22 39 24 66
rect 29 39 31 66
<< polyct0 >>
rect 19 32 21 34
<< polyct1 >>
rect 11 42 13 44
rect 34 31 36 33
<< ndifct0 >>
rect 14 14 16 16
rect 24 8 26 10
rect 34 14 36 16
<< ndifct1 >>
rect 4 14 6 16
<< pdifct0 >>
rect 7 62 9 64
rect 34 62 36 64
rect 34 55 36 57
<< pdifct1 >>
rect 17 55 19 57
<< alu0 >>
rect 5 62 7 64
rect 9 62 11 64
rect 5 61 11 62
rect 32 62 34 64
rect 36 62 38 64
rect 32 57 38 62
rect 32 55 34 57
rect 36 55 38 57
rect 32 54 38 55
rect 18 34 22 38
rect 18 32 19 34
rect 21 32 22 34
rect 18 30 22 32
rect 12 16 38 18
rect 12 14 14 16
rect 16 14 34 16
rect 36 14 38 16
rect 12 13 18 14
rect 32 13 38 14
rect 22 10 28 11
rect 22 8 24 10
rect 26 8 28 10
<< labels >>
rlabel alu0 25 16 25 16 6 n1
rlabel ndifct0 35 15 35 15 6 n1
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 36 12 36 6 b
rlabel alu1 12 56 12 56 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 20 24 20 24 6 b
rlabel alu1 28 32 28 32 6 a1
rlabel alu1 20 40 20 40 6 a2
rlabel alu1 28 44 28 44 6 a2
rlabel alu1 20 56 20 56 6 z
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 36 24 36 24 6 a1
<< end >>
