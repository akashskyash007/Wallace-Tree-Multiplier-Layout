magic
tech scmos
timestamp 1199979791
<< ab >>
rect -12 0 308 88
<< alu1 >>
rect -10 65 -6 91
rect -10 63 -9 65
rect -7 63 -6 65
rect -10 49 -6 63
rect -10 47 -9 49
rect -7 47 -6 49
rect -10 33 -6 47
rect -10 31 -9 33
rect -7 31 -6 33
rect -10 17 -6 31
rect -10 15 -9 17
rect -7 15 -6 17
rect -10 1 -6 15
rect -10 -1 -9 1
rect -7 -1 -6 1
rect -10 -3 -6 -1
<< alu2 >>
rect -11 65 307 66
rect -11 63 -9 65
rect -7 63 307 65
rect -11 62 307 63
rect -11 49 307 50
rect -11 47 -9 49
rect -7 47 307 49
rect -11 46 307 47
rect -11 33 307 34
rect -11 31 -9 33
rect -7 31 307 33
rect -11 30 307 31
rect -11 17 307 18
rect -11 15 -9 17
rect -7 15 7 17
rect 9 15 23 17
rect 25 15 39 17
rect 41 15 55 17
rect 57 15 71 17
rect 73 15 87 17
rect 89 15 103 17
rect 105 15 119 17
rect 121 15 135 17
rect 137 15 151 17
rect 153 15 167 17
rect 169 15 183 17
rect 185 15 199 17
rect 201 15 215 17
rect 217 15 231 17
rect 233 15 247 17
rect 249 15 263 17
rect 265 15 279 17
rect 281 15 295 17
rect 297 15 307 17
rect -11 14 307 15
rect -11 1 307 2
rect -11 -1 -9 1
rect -7 -1 307 1
rect -11 -2 307 -1
<< alu3 >>
rect 6 73 10 90
rect 6 71 7 73
rect 9 71 10 73
rect 6 57 10 71
rect 6 55 7 57
rect 9 55 10 57
rect 6 41 10 55
rect 6 39 7 41
rect 9 39 10 41
rect 6 25 10 39
rect 6 23 7 25
rect 9 23 10 25
rect 6 17 10 23
rect 6 15 7 17
rect 9 15 10 17
rect 6 -2 10 15
rect 22 17 26 90
rect 22 15 23 17
rect 25 15 26 17
rect 22 -2 26 15
rect 38 17 42 90
rect 38 15 39 17
rect 41 15 42 17
rect 38 -2 42 15
rect 54 17 58 90
rect 54 15 55 17
rect 57 15 58 17
rect 54 -2 58 15
rect 70 17 74 90
rect 70 15 71 17
rect 73 15 74 17
rect 70 -2 74 15
rect 86 17 90 90
rect 86 15 87 17
rect 89 15 90 17
rect 86 -2 90 15
rect 102 17 106 90
rect 102 15 103 17
rect 105 15 106 17
rect 102 -2 106 15
rect 118 17 122 90
rect 118 15 119 17
rect 121 15 122 17
rect 118 -2 122 15
rect 134 17 138 90
rect 134 15 135 17
rect 137 15 138 17
rect 134 -2 138 15
rect 150 17 154 90
rect 150 15 151 17
rect 153 15 154 17
rect 150 -2 154 15
rect 166 17 170 90
rect 166 15 167 17
rect 169 15 170 17
rect 166 -2 170 15
rect 182 17 186 90
rect 182 15 183 17
rect 185 15 186 17
rect 182 -2 186 15
rect 198 17 202 90
rect 198 15 199 17
rect 201 15 202 17
rect 198 -2 202 15
rect 214 17 218 90
rect 214 15 215 17
rect 217 15 218 17
rect 214 -2 218 15
rect 230 17 234 90
rect 230 15 231 17
rect 233 15 234 17
rect 230 -2 234 15
rect 246 17 250 90
rect 246 15 247 17
rect 249 15 250 17
rect 246 -2 250 15
rect 262 17 266 90
rect 262 15 263 17
rect 265 15 266 17
rect 262 -2 266 15
rect 278 17 282 90
rect 278 15 279 17
rect 281 15 282 17
rect 278 -2 282 15
rect 294 17 298 90
rect 294 15 295 17
rect 297 15 298 17
rect 294 -2 298 15
<< alu4 >>
rect -11 73 307 74
rect -11 71 7 73
rect 9 71 307 73
rect -11 70 307 71
rect -11 57 307 58
rect -11 55 7 57
rect 9 55 307 57
rect -11 54 307 55
rect -11 41 307 42
rect -11 39 7 41
rect 9 39 307 41
rect -11 38 307 39
rect -11 25 307 26
rect -11 23 -1 25
rect 1 23 7 25
rect 9 23 15 25
rect 17 23 31 25
rect 33 23 47 25
rect 49 23 63 25
rect 65 23 79 25
rect 81 23 95 25
rect 97 23 111 25
rect 113 23 127 25
rect 129 23 143 25
rect 145 23 159 25
rect 161 23 175 25
rect 177 23 191 25
rect 193 23 207 25
rect 209 23 223 25
rect 225 23 239 25
rect 241 23 255 25
rect 257 23 271 25
rect 273 23 287 25
rect 289 23 303 25
rect 305 23 307 25
rect -11 22 307 23
<< alu5 >>
rect -2 25 2 90
rect -2 23 -1 25
rect 1 23 2 25
rect -2 -2 2 23
rect 14 25 18 90
rect 14 23 15 25
rect 17 23 18 25
rect 14 -2 18 23
rect 30 25 34 90
rect 30 23 31 25
rect 33 23 34 25
rect 30 -2 34 23
rect 46 25 50 90
rect 46 23 47 25
rect 49 23 50 25
rect 46 -2 50 23
rect 62 25 66 90
rect 62 23 63 25
rect 65 23 66 25
rect 62 -2 66 23
rect 78 25 82 90
rect 78 23 79 25
rect 81 23 82 25
rect 78 -2 82 23
rect 94 25 98 90
rect 94 23 95 25
rect 97 23 98 25
rect 94 -2 98 23
rect 110 25 114 90
rect 110 23 111 25
rect 113 23 114 25
rect 110 -2 114 23
rect 126 25 130 90
rect 126 23 127 25
rect 129 23 130 25
rect 126 -2 130 23
rect 142 25 146 90
rect 142 23 143 25
rect 145 23 146 25
rect 142 -2 146 23
rect 158 25 162 90
rect 158 23 159 25
rect 161 23 162 25
rect 158 -2 162 23
rect 174 25 178 90
rect 174 23 175 25
rect 177 23 178 25
rect 174 -2 178 23
rect 190 25 194 90
rect 190 23 191 25
rect 193 23 194 25
rect 190 -2 194 23
rect 206 25 210 90
rect 206 23 207 25
rect 209 23 210 25
rect 206 -2 210 23
rect 222 25 226 90
rect 222 23 223 25
rect 225 23 226 25
rect 222 -2 226 23
rect 238 25 242 90
rect 238 23 239 25
rect 241 23 242 25
rect 238 -2 242 23
rect 254 25 258 90
rect 254 23 255 25
rect 257 23 258 25
rect 254 -2 258 23
rect 270 25 274 90
rect 270 23 271 25
rect 273 23 274 25
rect 270 -2 274 23
rect 286 25 290 90
rect 286 23 287 25
rect 289 23 290 25
rect 286 -2 290 23
rect 302 25 306 90
rect 302 23 303 25
rect 305 23 306 25
rect 302 -2 306 23
<< via1 >>
rect -9 63 -7 65
rect -9 47 -7 49
rect -9 31 -7 33
rect -9 15 -7 17
rect -9 -1 -7 1
<< via2 >>
rect 7 15 9 17
rect 23 15 25 17
rect 39 15 41 17
rect 55 15 57 17
rect 71 15 73 17
rect 87 15 89 17
rect 103 15 105 17
rect 119 15 121 17
rect 135 15 137 17
rect 151 15 153 17
rect 167 15 169 17
rect 183 15 185 17
rect 199 15 201 17
rect 215 15 217 17
rect 231 15 233 17
rect 247 15 249 17
rect 263 15 265 17
rect 279 15 281 17
rect 295 15 297 17
<< via3 >>
rect 7 71 9 73
rect 7 55 9 57
rect 7 39 9 41
rect 7 23 9 25
<< via4 >>
rect -1 23 1 25
rect 15 23 17 25
rect 31 23 33 25
rect 47 23 49 25
rect 63 23 65 25
rect 79 23 81 25
rect 95 23 97 25
rect 111 23 113 25
rect 127 23 129 25
rect 143 23 145 25
rect 159 23 161 25
rect 175 23 177 25
rect 191 23 193 25
rect 207 23 209 25
rect 223 23 225 25
rect 239 23 241 25
rect 255 23 257 25
rect 271 23 273 25
rect 287 23 289 25
rect 303 23 305 25
<< end >>
