magic
tech scmos
timestamp 1199202265
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 31 39
rect 9 35 19 37
rect 21 35 27 37
rect 29 35 31 37
rect 9 33 31 35
rect 9 30 11 33
rect 19 30 21 33
rect 9 6 11 10
rect 19 6 21 10
<< ndif >>
rect 2 21 9 30
rect 2 19 4 21
rect 6 19 9 21
rect 2 14 9 19
rect 2 12 4 14
rect 6 12 9 14
rect 2 10 9 12
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 10 19 19
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 21 29 26
rect 21 19 24 21
rect 26 19 29 21
rect 21 17 29 19
rect 21 10 27 17
<< pdif >>
rect 4 55 9 69
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 67 19 69
rect 11 65 14 67
rect 16 65 19 67
rect 11 59 19 65
rect 11 57 14 59
rect 16 57 19 59
rect 11 42 19 57
rect 21 53 29 69
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 67 38 69
rect 31 65 34 67
rect 36 65 38 67
rect 31 59 38 65
rect 31 57 34 59
rect 36 57 38 59
rect 31 42 38 57
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 23 53 27 55
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 2 44 4 46
rect 6 44 24 46
rect 26 44 27 46
rect 2 42 27 44
rect 2 30 6 42
rect 34 38 38 47
rect 17 37 38 38
rect 17 35 19 37
rect 21 35 27 37
rect 29 35 38 37
rect 17 34 38 35
rect 2 28 17 30
rect 2 26 14 28
rect 16 26 17 28
rect 13 21 17 26
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect 34 25 38 34
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 10 11 30
rect 19 10 21 30
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
<< polyct1 >>
rect 19 35 21 37
rect 27 35 29 37
<< ndifct0 >>
rect 4 19 6 21
rect 4 12 6 14
rect 24 26 26 28
rect 24 19 26 21
<< ndifct1 >>
rect 14 26 16 28
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 65 16 67
rect 14 57 16 59
rect 34 65 36 67
rect 34 57 36 59
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 51 26 53
rect 24 44 26 46
<< alu0 >>
rect 13 67 17 68
rect 13 65 14 67
rect 16 65 17 67
rect 13 59 17 65
rect 13 57 14 59
rect 16 57 17 59
rect 13 55 17 57
rect 33 67 37 68
rect 33 65 34 67
rect 36 65 37 67
rect 33 59 37 65
rect 33 57 34 59
rect 36 57 37 59
rect 33 55 37 57
rect 2 21 8 22
rect 2 19 4 21
rect 6 19 8 21
rect 2 14 8 19
rect 22 28 28 29
rect 22 26 24 28
rect 26 26 28 28
rect 22 21 28 26
rect 22 19 24 21
rect 26 19 28 21
rect 2 12 4 14
rect 6 12 8 14
rect 22 12 28 19
<< labels >>
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel polyct1 20 36 20 36 6 a
rlabel alu1 20 44 20 44 6 z
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 36 36 36 6 a
<< end >>
