magic
tech scmos
timestamp 1199469914
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -5 48 95 105
<< pwell >>
rect -5 -5 95 48
<< poly >>
rect 13 93 15 98
rect 25 93 27 98
rect 37 93 39 98
rect 49 93 51 98
rect 61 93 63 98
rect 73 93 75 98
rect 13 48 15 60
rect 25 57 27 60
rect 25 55 33 57
rect 25 54 29 55
rect 27 53 29 54
rect 31 53 33 55
rect 27 51 33 53
rect 37 53 39 60
rect 49 53 51 60
rect 61 57 63 60
rect 37 51 51 53
rect 13 46 23 48
rect 17 44 19 46
rect 21 44 23 46
rect 17 42 23 44
rect 21 39 23 42
rect 29 39 31 51
rect 37 49 43 51
rect 45 49 51 51
rect 37 47 51 49
rect 37 39 39 47
rect 49 39 51 47
rect 57 55 63 57
rect 57 53 59 55
rect 61 53 63 55
rect 57 51 63 53
rect 57 39 59 51
rect 73 48 75 60
rect 67 46 75 48
rect 67 45 69 46
rect 65 44 69 45
rect 71 44 75 46
rect 65 42 75 44
rect 65 39 67 42
rect 21 2 23 6
rect 29 2 31 6
rect 37 2 39 6
rect 49 2 51 6
rect 57 2 59 6
rect 65 2 67 6
<< ndif >>
rect 12 11 21 39
rect 12 9 15 11
rect 17 9 21 11
rect 12 6 21 9
rect 23 6 29 39
rect 31 6 37 39
rect 39 21 49 39
rect 39 19 43 21
rect 45 19 49 21
rect 39 6 49 19
rect 51 6 57 39
rect 59 6 65 39
rect 67 21 75 39
rect 67 19 71 21
rect 73 19 75 21
rect 67 11 75 19
rect 67 9 71 11
rect 73 9 75 11
rect 67 6 75 9
<< pdif >>
rect 4 91 13 93
rect 4 89 7 91
rect 9 89 13 91
rect 4 81 13 89
rect 4 79 7 81
rect 9 79 13 81
rect 4 71 13 79
rect 4 69 7 71
rect 9 69 13 71
rect 4 60 13 69
rect 15 81 25 93
rect 15 79 19 81
rect 21 79 25 81
rect 15 71 25 79
rect 15 69 19 71
rect 21 69 25 71
rect 15 60 25 69
rect 27 91 37 93
rect 27 89 31 91
rect 33 89 37 91
rect 27 81 37 89
rect 27 79 31 81
rect 33 79 37 81
rect 27 60 37 79
rect 39 81 49 93
rect 39 79 43 81
rect 45 79 49 81
rect 39 71 49 79
rect 39 69 43 71
rect 45 69 49 71
rect 39 60 49 69
rect 51 91 61 93
rect 51 89 55 91
rect 57 89 61 91
rect 51 81 61 89
rect 51 79 55 81
rect 57 79 61 81
rect 51 60 61 79
rect 63 81 73 93
rect 63 79 67 81
rect 69 79 73 81
rect 63 71 73 79
rect 63 69 67 71
rect 69 69 73 71
rect 63 60 73 69
rect 75 91 84 93
rect 75 89 79 91
rect 81 89 84 91
rect 75 81 84 89
rect 75 79 79 81
rect 81 79 84 81
rect 75 71 84 79
rect 75 69 79 71
rect 81 69 84 71
rect 75 60 84 69
<< alu1 >>
rect -2 91 92 100
rect -2 89 7 91
rect 9 89 31 91
rect 33 89 55 91
rect 57 89 79 91
rect 81 89 92 91
rect -2 88 92 89
rect 6 81 10 88
rect 6 79 7 81
rect 9 79 10 81
rect 6 71 10 79
rect 6 69 7 71
rect 9 69 10 71
rect 6 67 10 69
rect 18 81 22 83
rect 18 79 19 81
rect 21 79 22 81
rect 18 72 22 79
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 77 34 79
rect 42 81 46 83
rect 42 79 43 81
rect 45 79 46 81
rect 42 72 46 79
rect 54 81 58 88
rect 54 79 55 81
rect 57 79 58 81
rect 54 77 58 79
rect 66 81 70 83
rect 66 79 67 81
rect 69 79 70 81
rect 66 72 70 79
rect 78 81 82 88
rect 78 79 79 81
rect 81 79 82 81
rect 18 71 73 72
rect 18 69 19 71
rect 21 69 43 71
rect 45 69 67 71
rect 69 69 73 71
rect 18 68 73 69
rect 78 71 82 79
rect 78 69 79 71
rect 81 69 82 71
rect 18 63 22 68
rect 78 67 82 69
rect 8 57 22 63
rect 27 58 63 62
rect 8 22 12 57
rect 27 55 32 58
rect 27 53 29 55
rect 31 53 32 55
rect 57 55 63 58
rect 57 53 59 55
rect 61 53 63 55
rect 17 46 23 52
rect 17 44 19 46
rect 21 44 23 46
rect 17 32 23 44
rect 27 37 32 53
rect 38 51 52 53
rect 38 49 43 51
rect 45 49 52 51
rect 38 47 52 49
rect 57 48 63 53
rect 48 37 52 47
rect 68 46 73 63
rect 68 44 69 46
rect 71 44 73 46
rect 68 32 73 44
rect 17 28 73 32
rect 8 21 47 22
rect 8 19 43 21
rect 45 19 47 21
rect 8 17 47 19
rect 70 21 74 23
rect 70 19 71 21
rect 73 19 74 21
rect 70 12 74 19
rect -2 11 92 12
rect -2 9 15 11
rect 17 9 71 11
rect 73 9 92 11
rect -2 7 92 9
rect -2 5 83 7
rect 85 5 92 7
rect -2 0 92 5
<< ptie >>
rect 81 7 87 9
rect 81 5 83 7
rect 85 5 87 7
rect 81 3 87 5
<< nmos >>
rect 21 6 23 39
rect 29 6 31 39
rect 37 6 39 39
rect 49 6 51 39
rect 57 6 59 39
rect 65 6 67 39
<< pmos >>
rect 13 60 15 93
rect 25 60 27 93
rect 37 60 39 93
rect 49 60 51 93
rect 61 60 63 93
rect 73 60 75 93
<< polyct1 >>
rect 29 53 31 55
rect 19 44 21 46
rect 43 49 45 51
rect 59 53 61 55
rect 69 44 71 46
<< ndifct1 >>
rect 15 9 17 11
rect 43 19 45 21
rect 71 19 73 21
rect 71 9 73 11
<< ptiect1 >>
rect 83 5 85 7
<< pdifct1 >>
rect 7 89 9 91
rect 7 79 9 81
rect 7 69 9 71
rect 19 79 21 81
rect 19 69 21 71
rect 31 89 33 91
rect 31 79 33 81
rect 43 79 45 81
rect 43 69 45 71
rect 55 89 57 91
rect 55 79 57 81
rect 67 79 69 81
rect 67 69 69 71
rect 79 89 81 91
rect 79 79 81 81
rect 79 69 81 71
<< labels >>
rlabel alu1 10 40 10 40 6 z
rlabel alu1 30 20 30 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 30 30 30 30 6 c
rlabel alu1 20 40 20 40 6 c
rlabel alu1 30 50 30 50 6 b
rlabel pdifct1 20 70 20 70 6 z
rlabel alu1 30 70 30 70 6 z
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 40 20 40 20 6 z
rlabel alu1 40 30 40 30 6 c
rlabel alu1 50 30 50 30 6 c
rlabel alu1 40 50 40 50 6 a
rlabel alu1 50 45 50 45 6 a
rlabel alu1 40 60 40 60 6 b
rlabel alu1 50 60 50 60 6 b
rlabel alu1 40 70 40 70 6 z
rlabel alu1 50 70 50 70 6 z
rlabel alu1 45 94 45 94 6 vdd
rlabel alu1 60 30 60 30 6 c
rlabel polyct1 70 45 70 45 6 c
rlabel alu1 60 55 60 55 6 b
rlabel alu1 60 70 60 70 6 z
rlabel alu1 70 70 70 70 6 z
<< end >>
