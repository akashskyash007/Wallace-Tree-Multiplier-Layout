magic
tech scmos
timestamp 1199543276
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -2 48 62 104
<< pwell >>
rect -2 -4 62 48
<< poly >>
rect 35 95 37 98
rect 47 95 49 98
rect 15 85 17 88
rect 23 85 25 88
rect 15 53 17 55
rect 11 51 17 53
rect 23 53 25 55
rect 23 51 31 53
rect 11 43 13 51
rect 23 49 27 51
rect 29 49 31 51
rect 23 47 31 49
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 35 41 37 55
rect 47 41 49 55
rect 17 39 19 41
rect 21 39 49 41
rect 17 37 23 39
rect 11 25 13 37
rect 23 31 31 33
rect 23 29 27 31
rect 29 29 31 31
rect 23 27 31 29
rect 23 25 25 27
rect 35 25 37 39
rect 47 25 49 39
rect 11 12 13 15
rect 23 12 25 15
rect 35 2 37 5
rect 47 2 49 5
<< ndif >>
rect 3 15 11 25
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 15 23 19
rect 25 15 35 25
rect 3 11 9 15
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 27 11 35 15
rect 27 9 29 11
rect 31 9 35 11
rect 27 5 35 9
rect 37 21 47 25
rect 37 19 41 21
rect 43 19 47 21
rect 37 5 47 19
rect 49 21 57 25
rect 49 19 53 21
rect 55 19 57 21
rect 49 11 57 19
rect 49 9 53 11
rect 55 9 57 11
rect 49 5 57 9
<< pdif >>
rect 27 91 35 95
rect 27 89 29 91
rect 31 89 35 91
rect 27 85 35 89
rect 3 81 15 85
rect 3 79 5 81
rect 7 79 15 81
rect 3 55 15 79
rect 17 55 23 85
rect 25 55 35 85
rect 37 81 47 95
rect 37 79 41 81
rect 43 79 47 81
rect 37 71 47 79
rect 37 69 41 71
rect 43 69 47 71
rect 37 61 47 69
rect 37 59 41 61
rect 43 59 47 61
rect 37 55 47 59
rect 49 91 57 95
rect 49 89 53 91
rect 55 89 57 91
rect 49 81 57 89
rect 49 79 53 81
rect 55 79 57 81
rect 49 71 57 79
rect 49 69 53 71
rect 55 69 57 71
rect 49 61 57 69
rect 49 59 53 61
rect 55 59 57 61
rect 49 55 57 59
<< alu1 >>
rect -2 95 62 100
rect -2 93 5 95
rect 7 93 17 95
rect 19 93 62 95
rect -2 91 62 93
rect -2 89 29 91
rect 31 89 53 91
rect 55 89 62 91
rect -2 88 62 89
rect 4 81 8 82
rect 4 79 5 81
rect 7 79 20 81
rect 4 78 8 79
rect 8 41 12 72
rect 8 39 9 41
rect 11 39 12 41
rect 8 28 12 39
rect 18 42 20 79
rect 28 52 32 82
rect 26 51 32 52
rect 26 49 27 51
rect 29 49 32 51
rect 26 48 32 49
rect 18 41 22 42
rect 18 39 19 41
rect 21 39 22 41
rect 18 38 22 39
rect 18 22 20 38
rect 28 32 32 48
rect 26 31 32 32
rect 26 29 27 31
rect 29 29 32 31
rect 26 28 32 29
rect 16 21 20 22
rect 16 19 17 21
rect 19 19 20 21
rect 16 18 20 19
rect 28 18 32 28
rect 38 81 44 82
rect 38 79 41 81
rect 43 79 44 81
rect 38 78 44 79
rect 52 81 56 88
rect 52 79 53 81
rect 55 79 56 81
rect 38 72 42 78
rect 38 71 44 72
rect 38 69 41 71
rect 43 69 44 71
rect 38 68 44 69
rect 52 71 56 79
rect 52 69 53 71
rect 55 69 56 71
rect 38 62 42 68
rect 38 61 44 62
rect 38 59 41 61
rect 43 59 44 61
rect 38 58 44 59
rect 52 61 56 69
rect 52 59 53 61
rect 55 59 56 61
rect 52 58 56 59
rect 38 22 42 58
rect 38 21 44 22
rect 38 19 41 21
rect 43 19 44 21
rect 38 18 44 19
rect 52 21 56 22
rect 52 19 53 21
rect 55 19 56 21
rect 52 12 56 19
rect -2 11 62 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 53 11
rect 55 9 62 11
rect -2 0 62 9
<< ntie >>
rect 3 95 21 97
rect 3 93 5 95
rect 7 93 17 95
rect 19 93 21 95
rect 3 91 21 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 5 37 25
rect 47 5 49 25
<< pmos >>
rect 15 55 17 85
rect 23 55 25 85
rect 35 55 37 95
rect 47 55 49 95
<< polyct1 >>
rect 27 49 29 51
rect 9 39 11 41
rect 19 39 21 41
rect 27 29 29 31
<< ndifct1 >>
rect 17 19 19 21
rect 5 9 7 11
rect 29 9 31 11
rect 41 19 43 21
rect 53 19 55 21
rect 53 9 55 11
<< ntiect1 >>
rect 5 93 7 95
rect 17 93 19 95
<< pdifct1 >>
rect 29 89 31 91
rect 5 79 7 81
rect 41 79 43 81
rect 41 69 43 71
rect 41 59 43 61
rect 53 89 55 91
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
<< labels >>
rlabel alu1 10 50 10 50 6 i1
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 40 50 40 50 6 q
rlabel alu1 30 50 30 50 6 i0
rlabel alu1 30 94 30 94 6 vdd
<< end >>
