magic
tech scmos
timestamp 1199203611
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 38 63 63 65
rect 28 58 34 60
rect 28 56 30 58
rect 32 56 34 58
rect 18 50 20 55
rect 28 54 34 56
rect 28 50 30 54
rect 38 50 40 63
rect 61 59 63 63
rect 48 50 50 55
rect 18 35 20 38
rect 9 33 20 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 28 30 30 38
rect 38 34 40 38
rect 48 34 50 38
rect 61 35 63 47
rect 47 32 53 34
rect 47 30 49 32
rect 51 30 53 32
rect 12 25 14 29
rect 22 25 24 29
rect 28 28 34 30
rect 32 25 34 28
rect 42 28 53 30
rect 57 33 63 35
rect 57 31 59 33
rect 61 31 63 33
rect 57 29 63 31
rect 42 25 44 28
rect 61 25 63 29
rect 12 14 14 19
rect 22 11 24 19
rect 32 15 34 19
rect 42 15 44 19
rect 61 11 63 19
rect 22 9 63 11
<< ndif >>
rect 4 19 12 25
rect 14 23 22 25
rect 14 21 17 23
rect 19 21 22 23
rect 14 19 22 21
rect 24 23 32 25
rect 24 21 27 23
rect 29 21 32 23
rect 24 19 32 21
rect 34 23 42 25
rect 34 21 37 23
rect 39 21 42 23
rect 34 19 42 21
rect 44 23 61 25
rect 44 21 56 23
rect 58 21 61 23
rect 44 19 61 21
rect 63 23 70 25
rect 63 21 66 23
rect 68 21 70 23
rect 63 19 70 21
rect 4 16 10 19
rect 4 14 6 16
rect 8 14 10 16
rect 4 12 10 14
<< pdif >>
rect 52 59 59 61
rect 52 57 55 59
rect 57 57 61 59
rect 52 50 61 57
rect 8 48 18 50
rect 8 46 11 48
rect 13 46 18 48
rect 8 38 18 46
rect 20 42 28 50
rect 20 40 23 42
rect 25 40 28 42
rect 20 38 28 40
rect 30 42 38 50
rect 30 40 33 42
rect 35 40 38 42
rect 30 38 38 40
rect 40 42 48 50
rect 40 40 43 42
rect 45 40 48 42
rect 40 38 48 40
rect 50 47 61 50
rect 63 53 68 59
rect 63 51 70 53
rect 63 49 66 51
rect 68 49 70 51
rect 63 47 70 49
rect 50 38 59 47
<< alu1 >>
rect -2 67 74 72
rect -2 65 5 67
rect 7 65 13 67
rect 15 65 74 67
rect -2 64 74 65
rect 34 44 38 51
rect 32 42 38 44
rect 32 40 33 42
rect 35 40 38 42
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 2 21 6 29
rect 32 37 38 40
rect 32 34 36 37
rect 25 30 36 34
rect 25 23 31 30
rect 50 37 62 43
rect 25 21 27 23
rect 29 21 31 23
rect 25 20 31 21
rect 58 33 62 37
rect 58 31 59 33
rect 61 31 62 33
rect 58 29 62 31
rect -2 7 74 8
rect -2 5 16 7
rect 18 5 74 7
rect -2 0 74 5
<< ptie >>
rect 14 7 20 9
rect 14 5 16 7
rect 18 5 20 7
rect 14 3 20 5
<< ntie >>
rect 3 67 17 69
rect 3 65 5 67
rect 7 65 13 67
rect 15 65 17 67
rect 3 63 17 65
<< nmos >>
rect 12 19 14 25
rect 22 19 24 25
rect 32 19 34 25
rect 42 19 44 25
rect 61 19 63 25
<< pmos >>
rect 18 38 20 50
rect 28 38 30 50
rect 38 38 40 50
rect 48 38 50 50
rect 61 47 63 59
<< polyct0 >>
rect 30 56 32 58
rect 49 30 51 32
<< polyct1 >>
rect 11 31 13 33
rect 59 31 61 33
<< ndifct0 >>
rect 17 21 19 23
rect 37 21 39 23
rect 56 21 58 23
rect 66 21 68 23
rect 6 14 8 16
<< ndifct1 >>
rect 27 21 29 23
<< ntiect1 >>
rect 5 65 7 67
rect 13 65 15 67
<< ptiect1 >>
rect 16 5 18 7
<< pdifct0 >>
rect 55 57 57 59
rect 11 46 13 48
rect 23 40 25 42
rect 43 40 45 42
rect 66 49 68 51
<< pdifct1 >>
rect 33 40 35 42
<< alu0 >>
rect 10 48 14 64
rect 53 59 59 64
rect 28 58 49 59
rect 28 56 30 58
rect 32 56 49 58
rect 53 57 55 59
rect 57 57 59 59
rect 53 56 59 57
rect 28 55 49 56
rect 45 52 49 55
rect 45 51 70 52
rect 10 46 11 48
rect 13 46 14 48
rect 10 44 14 46
rect 45 49 66 51
rect 68 49 70 51
rect 45 48 70 49
rect 17 42 27 43
rect 17 40 23 42
rect 25 40 27 42
rect 17 39 27 40
rect 17 25 21 39
rect 41 42 46 44
rect 41 40 43 42
rect 45 40 46 42
rect 41 38 46 40
rect 16 23 21 25
rect 16 21 17 23
rect 19 21 21 23
rect 16 19 21 21
rect 41 24 45 38
rect 35 23 45 24
rect 35 21 37 23
rect 39 21 45 23
rect 35 20 45 21
rect 48 32 52 34
rect 48 30 49 32
rect 51 30 52 32
rect 17 17 21 19
rect 48 17 52 30
rect 66 25 70 48
rect 4 16 10 17
rect 4 14 6 16
rect 8 14 10 16
rect 4 8 10 14
rect 17 13 52 17
rect 55 23 59 25
rect 55 21 56 23
rect 58 21 59 23
rect 55 8 59 21
rect 65 23 70 25
rect 65 21 66 23
rect 68 21 70 23
rect 65 19 70 21
<< labels >>
rlabel alu0 19 28 19 28 6 an
rlabel alu0 22 41 22 41 6 an
rlabel alu0 50 23 50 23 6 an
rlabel alu0 40 22 40 22 6 ai
rlabel alu0 43 32 43 32 6 ai
rlabel alu0 38 57 38 57 6 bn
rlabel alu0 68 35 68 35 6 bn
rlabel alu0 57 50 57 50 6 bn
rlabel alu1 4 28 4 28 6 a
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 28 28 28 28 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 52 40 52 40 6 b
rlabel alu1 36 44 36 44 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 36 60 36 6 b
<< end >>
