magic
tech scmos
timestamp 1199203699
<< ab >>
rect 0 0 120 72
<< nwell >>
rect -5 32 125 77
<< pwell >>
rect -5 -5 125 32
<< poly >>
rect 17 63 19 68
rect 29 63 31 68
rect 39 63 41 68
rect 49 63 51 68
rect 77 66 79 70
rect 2 49 8 51
rect 2 47 4 49
rect 6 47 8 49
rect 2 45 8 47
rect 6 41 8 45
rect 89 61 91 66
rect 99 61 101 66
rect 109 61 111 66
rect 77 47 79 50
rect 65 45 79 47
rect 17 41 19 44
rect 6 39 19 41
rect 9 21 11 39
rect 29 34 31 44
rect 39 35 41 44
rect 49 41 51 44
rect 65 43 67 45
rect 69 43 71 45
rect 65 41 71 43
rect 45 39 51 41
rect 45 37 47 39
rect 49 37 51 39
rect 89 37 91 45
rect 45 35 51 37
rect 55 35 91 37
rect 99 36 101 45
rect 17 32 31 34
rect 35 33 41 35
rect 17 30 19 32
rect 21 30 23 32
rect 17 28 23 30
rect 35 31 37 33
rect 39 31 41 33
rect 35 29 41 31
rect 20 21 22 28
rect 39 27 41 29
rect 30 21 32 25
rect 39 24 42 27
rect 40 21 42 24
rect 47 21 49 35
rect 55 33 57 35
rect 59 33 61 35
rect 55 31 61 33
rect 65 29 71 31
rect 65 27 67 29
rect 69 27 71 29
rect 65 25 71 27
rect 69 22 71 25
rect 81 19 83 35
rect 95 34 101 36
rect 109 35 111 45
rect 95 32 97 34
rect 99 32 101 34
rect 95 30 101 32
rect 99 25 101 30
rect 105 33 111 35
rect 105 31 107 33
rect 109 31 111 33
rect 105 29 111 31
rect 91 19 93 24
rect 99 22 103 25
rect 101 19 103 22
rect 108 19 110 29
rect 9 4 11 12
rect 20 8 22 12
rect 30 4 32 12
rect 40 7 42 12
rect 47 7 49 12
rect 9 2 32 4
rect 69 4 71 15
rect 81 8 83 12
rect 91 4 93 12
rect 101 7 103 12
rect 108 7 110 12
rect 69 2 93 4
<< ndif >>
rect 2 19 9 21
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 4 12 9 15
rect 11 16 20 21
rect 11 14 15 16
rect 17 14 20 16
rect 11 12 20 14
rect 22 16 30 21
rect 22 14 25 16
rect 27 14 30 16
rect 22 12 30 14
rect 32 17 40 21
rect 32 15 35 17
rect 37 15 40 17
rect 32 12 40 15
rect 42 12 47 21
rect 49 12 57 21
rect 62 20 69 22
rect 62 18 64 20
rect 66 18 69 20
rect 62 15 69 18
rect 71 19 79 22
rect 71 15 81 19
rect 51 10 57 12
rect 51 8 53 10
rect 55 8 57 10
rect 51 6 57 8
rect 73 12 81 15
rect 83 17 91 19
rect 83 15 86 17
rect 88 15 91 17
rect 83 12 91 15
rect 93 17 101 19
rect 93 15 96 17
rect 98 15 101 17
rect 93 12 101 15
rect 103 12 108 19
rect 110 12 118 19
rect 73 10 75 12
rect 77 10 79 12
rect 73 8 79 10
rect 112 7 118 12
rect 112 5 114 7
rect 116 5 118 7
rect 112 3 118 5
<< pdif >>
rect 21 67 27 69
rect 21 65 23 67
rect 25 65 27 67
rect 21 63 27 65
rect 81 67 87 69
rect 81 66 83 67
rect 12 50 17 63
rect 10 48 17 50
rect 10 46 12 48
rect 14 46 17 48
rect 10 44 17 46
rect 19 44 29 63
rect 31 48 39 63
rect 31 46 34 48
rect 36 46 39 48
rect 31 44 39 46
rect 41 49 49 63
rect 41 47 44 49
rect 46 47 49 49
rect 41 44 49 47
rect 51 59 56 63
rect 72 60 77 66
rect 51 57 58 59
rect 51 55 54 57
rect 56 55 58 57
rect 51 53 58 55
rect 70 58 77 60
rect 70 56 72 58
rect 74 56 77 58
rect 70 54 77 56
rect 51 44 56 53
rect 72 50 77 54
rect 79 65 83 66
rect 85 65 87 67
rect 79 61 87 65
rect 79 50 89 61
rect 81 45 89 50
rect 91 49 99 61
rect 91 47 94 49
rect 96 47 99 49
rect 91 45 99 47
rect 101 50 109 61
rect 101 48 104 50
rect 106 48 109 50
rect 101 45 109 48
rect 111 58 118 61
rect 111 56 114 58
rect 116 56 118 58
rect 111 54 118 56
rect 111 45 116 54
<< alu1 >>
rect -2 67 122 72
rect -2 65 23 67
rect 25 65 62 67
rect 64 65 83 67
rect 85 65 122 67
rect -2 64 122 65
rect 2 54 15 59
rect 2 49 7 54
rect 2 47 4 49
rect 6 47 7 49
rect 2 45 7 47
rect 18 32 22 35
rect 18 30 19 32
rect 21 30 22 32
rect 18 27 22 30
rect 10 21 22 27
rect 66 45 70 51
rect 66 43 67 45
rect 69 43 70 45
rect 66 42 70 43
rect 66 38 79 42
rect 66 29 70 38
rect 102 50 118 51
rect 102 48 104 50
rect 106 48 118 50
rect 102 47 118 48
rect 66 27 67 29
rect 69 27 70 29
rect 66 25 70 27
rect 114 18 118 47
rect 94 17 118 18
rect 94 15 96 17
rect 98 15 118 17
rect 94 14 118 15
rect -2 7 122 8
rect -2 5 63 7
rect 65 5 114 7
rect 116 5 122 7
rect -2 0 122 5
<< ptie >>
rect 61 7 67 9
rect 61 5 63 7
rect 65 5 67 7
rect 61 3 67 5
<< ntie >>
rect 60 67 66 69
rect 60 65 62 67
rect 64 65 66 67
rect 60 63 66 65
<< nmos >>
rect 9 12 11 21
rect 20 12 22 21
rect 30 12 32 21
rect 40 12 42 21
rect 47 12 49 21
rect 69 15 71 22
rect 81 12 83 19
rect 91 12 93 19
rect 101 12 103 19
rect 108 12 110 19
<< pmos >>
rect 17 44 19 63
rect 29 44 31 63
rect 39 44 41 63
rect 49 44 51 63
rect 77 50 79 66
rect 89 45 91 61
rect 99 45 101 61
rect 109 45 111 61
<< polyct0 >>
rect 47 37 49 39
rect 37 31 39 33
rect 57 33 59 35
rect 97 32 99 34
rect 107 31 109 33
<< polyct1 >>
rect 4 47 6 49
rect 67 43 69 45
rect 19 30 21 32
rect 67 27 69 29
<< ndifct0 >>
rect 4 17 6 19
rect 15 14 17 16
rect 25 14 27 16
rect 35 15 37 17
rect 64 18 66 20
rect 53 8 55 10
rect 86 15 88 17
rect 75 10 77 12
<< ndifct1 >>
rect 96 15 98 17
rect 114 5 116 7
<< ntiect1 >>
rect 62 65 64 67
<< ptiect1 >>
rect 63 5 65 7
<< pdifct0 >>
rect 12 46 14 48
rect 34 46 36 48
rect 44 47 46 49
rect 54 55 56 57
rect 72 56 74 58
rect 94 47 96 49
rect 114 56 116 58
<< pdifct1 >>
rect 23 65 25 67
rect 83 65 85 67
rect 104 48 106 50
<< alu0 >>
rect 70 58 118 59
rect 26 57 58 58
rect 26 55 54 57
rect 56 55 58 57
rect 70 56 72 58
rect 74 56 114 58
rect 116 56 118 58
rect 70 55 118 56
rect 26 54 58 55
rect 26 50 30 54
rect 11 48 30 50
rect 11 46 12 48
rect 14 46 30 48
rect 11 39 15 46
rect 3 35 15 39
rect 3 19 7 35
rect 26 34 30 46
rect 33 48 37 50
rect 33 46 34 48
rect 36 46 37 48
rect 42 49 58 50
rect 42 47 44 49
rect 46 47 58 49
rect 42 46 58 47
rect 33 42 37 46
rect 33 39 50 42
rect 33 38 47 39
rect 46 37 47 38
rect 49 37 50 39
rect 26 33 41 34
rect 26 31 37 33
rect 39 31 41 33
rect 26 30 41 31
rect 46 26 50 37
rect 26 22 50 26
rect 54 36 58 46
rect 54 35 61 36
rect 54 33 57 35
rect 59 33 61 35
rect 54 32 61 33
rect 3 17 4 19
rect 6 17 7 19
rect 26 17 30 22
rect 54 18 58 32
rect 84 35 88 55
rect 93 49 97 51
rect 93 47 94 49
rect 96 47 97 49
rect 93 43 97 47
rect 93 39 110 43
rect 76 34 101 35
rect 76 32 97 34
rect 99 32 101 34
rect 76 31 101 32
rect 106 33 110 39
rect 106 31 107 33
rect 109 31 110 33
rect 76 21 80 31
rect 106 27 110 31
rect 3 15 7 17
rect 13 16 19 17
rect 13 14 15 16
rect 17 14 19 16
rect 13 8 19 14
rect 23 16 30 17
rect 23 14 25 16
rect 27 14 30 16
rect 33 17 58 18
rect 62 20 80 21
rect 62 18 64 20
rect 66 18 80 20
rect 62 17 80 18
rect 85 23 110 27
rect 85 17 89 23
rect 33 15 35 17
rect 37 15 58 17
rect 33 14 58 15
rect 85 15 86 17
rect 88 15 89 17
rect 23 13 30 14
rect 85 13 89 15
rect 73 12 79 13
rect 51 10 57 11
rect 51 8 53 10
rect 55 8 57 10
rect 73 10 75 12
rect 77 10 79 12
rect 73 8 79 10
<< labels >>
rlabel ndifct0 26 15 26 15 6 an
rlabel alu0 13 42 13 42 6 bn
rlabel alu0 5 27 5 27 6 bn
rlabel alu0 45 16 45 16 6 iz
rlabel alu0 33 32 33 32 6 bn
rlabel alu0 48 32 48 32 6 an
rlabel alu0 56 32 56 32 6 iz
rlabel alu0 35 44 35 44 6 an
rlabel alu0 50 48 50 48 6 iz
rlabel alu0 42 56 42 56 6 bn
rlabel alu0 71 19 71 19 6 cn
rlabel alu0 87 20 87 20 6 zn
rlabel alu0 108 33 108 33 6 zn
rlabel alu0 88 33 88 33 6 cn
rlabel alu0 95 45 95 45 6 zn
rlabel alu0 94 57 94 57 6 cn
rlabel alu1 12 24 12 24 6 a
rlabel alu1 20 28 20 28 6 a
rlabel alu1 4 52 4 52 6 b
rlabel alu1 12 56 12 56 6 b
rlabel alu1 60 4 60 4 6 vss
rlabel alu1 68 40 68 40 6 c
rlabel alu1 76 40 76 40 6 c
rlabel alu1 60 68 60 68 6 vdd
rlabel alu1 100 16 100 16 6 z
rlabel alu1 108 16 108 16 6 z
rlabel alu1 116 36 116 36 6 z
<< end >>
