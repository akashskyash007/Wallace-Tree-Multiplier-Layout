magic
tech scmos
timestamp 1199469125
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -5 48 75 105
<< pwell >>
rect -5 -5 75 48
<< poly >>
rect 33 89 35 94
rect 45 89 47 94
rect 57 89 59 94
rect 11 83 13 88
rect 11 52 13 63
rect 33 52 35 63
rect 45 52 47 63
rect 57 52 59 63
rect 11 50 22 52
rect 15 48 18 50
rect 20 48 22 50
rect 15 46 22 48
rect 33 50 41 52
rect 33 48 37 50
rect 39 48 41 50
rect 33 46 41 48
rect 45 50 53 52
rect 45 48 49 50
rect 51 48 53 50
rect 45 46 53 48
rect 57 50 63 52
rect 57 48 59 50
rect 61 48 63 50
rect 57 46 63 48
rect 15 37 17 46
rect 33 37 35 46
rect 45 37 47 46
rect 57 42 59 46
rect 53 40 59 42
rect 53 37 55 40
rect 15 22 17 27
rect 33 25 35 30
rect 45 20 47 25
rect 53 20 55 25
<< ndif >>
rect 7 35 15 37
rect 7 33 9 35
rect 11 33 15 35
rect 7 31 15 33
rect 10 27 15 31
rect 17 31 33 37
rect 17 29 21 31
rect 23 30 33 31
rect 35 35 45 37
rect 35 33 39 35
rect 41 33 45 35
rect 35 30 45 33
rect 23 29 31 30
rect 17 27 31 29
rect 40 25 45 30
rect 47 25 53 37
rect 55 31 64 37
rect 55 29 59 31
rect 61 29 64 31
rect 55 25 64 29
<< pdif >>
rect 49 91 55 93
rect 49 89 51 91
rect 53 89 55 91
rect 6 73 11 83
rect 3 71 11 73
rect 3 69 5 71
rect 7 69 11 71
rect 3 67 11 69
rect 6 63 11 67
rect 13 81 21 83
rect 13 79 17 81
rect 19 79 21 81
rect 13 75 21 79
rect 13 63 19 75
rect 28 69 33 89
rect 25 67 33 69
rect 25 65 27 67
rect 29 65 33 67
rect 25 63 33 65
rect 35 81 45 89
rect 35 79 39 81
rect 41 79 45 81
rect 35 63 45 79
rect 47 63 57 89
rect 59 83 64 89
rect 59 81 67 83
rect 59 79 63 81
rect 65 79 67 81
rect 59 77 67 79
rect 59 63 64 77
<< alu1 >>
rect -2 95 72 100
rect -2 93 9 95
rect 11 93 72 95
rect -2 91 72 93
rect -2 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 16 81 20 88
rect 16 79 17 81
rect 19 79 20 81
rect 16 77 20 79
rect 37 81 67 82
rect 37 79 39 81
rect 41 79 63 81
rect 65 79 67 81
rect 37 78 67 79
rect 4 71 22 73
rect 4 69 5 71
rect 7 69 22 71
rect 4 67 22 69
rect 26 67 30 69
rect 8 35 12 67
rect 26 65 27 67
rect 29 65 30 67
rect 26 51 30 65
rect 38 68 53 73
rect 38 52 42 68
rect 58 63 62 73
rect 16 50 30 51
rect 16 48 18 50
rect 20 48 30 50
rect 16 47 30 48
rect 26 42 30 47
rect 36 50 42 52
rect 36 48 37 50
rect 39 48 42 50
rect 36 46 42 48
rect 48 57 62 63
rect 48 50 52 57
rect 48 48 49 50
rect 51 48 52 50
rect 48 46 52 48
rect 57 50 63 52
rect 57 48 59 50
rect 61 48 63 50
rect 57 42 63 48
rect 26 38 42 42
rect 8 33 9 35
rect 11 33 12 35
rect 38 35 42 38
rect 38 33 39 35
rect 41 33 42 35
rect 8 27 12 33
rect 20 31 24 33
rect 38 31 42 33
rect 47 38 63 42
rect 20 29 21 31
rect 23 29 24 31
rect 20 12 24 29
rect 47 18 53 38
rect 58 31 62 33
rect 58 29 59 31
rect 61 29 62 31
rect 58 12 62 29
rect -2 7 72 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 72 7
rect -2 0 72 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 13 97
rect 7 93 9 95
rect 11 93 13 95
rect 7 91 13 93
<< nmos >>
rect 15 27 17 37
rect 33 30 35 37
rect 45 25 47 37
rect 53 25 55 37
<< pmos >>
rect 11 63 13 83
rect 33 63 35 89
rect 45 63 47 89
rect 57 63 59 89
<< polyct1 >>
rect 18 48 20 50
rect 37 48 39 50
rect 49 48 51 50
rect 59 48 61 50
<< ndifct1 >>
rect 9 33 11 35
rect 21 29 23 31
rect 39 33 41 35
rect 59 29 61 31
<< ntiect1 >>
rect 9 93 11 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 51 89 53 91
rect 5 69 7 71
rect 17 79 19 81
rect 27 65 29 67
rect 39 79 41 81
rect 63 79 65 81
<< labels >>
rlabel polyct1 19 49 19 49 6 zn
rlabel ndifct1 40 34 40 34 6 zn
rlabel pdifct1 28 66 28 66 6 zn
rlabel pdifct1 40 80 40 80 6 n2
rlabel pdifct1 64 80 64 80 6 n2
rlabel alu1 10 50 10 50 6 z
rlabel alu1 20 70 20 70 6 z
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 50 30 50 30 6 a1
rlabel alu1 50 70 50 70 6 b
rlabel alu1 50 55 50 55 6 a2
rlabel alu1 40 60 40 60 6 b
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 45 60 45 6 a1
rlabel alu1 60 65 60 65 6 a2
<< end >>
