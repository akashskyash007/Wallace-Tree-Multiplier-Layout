magic
tech scmos
timestamp 1199202103
<< ab >>
rect 0 0 88 80
<< nwell >>
rect -5 36 93 88
<< pwell >>
rect -5 -8 93 36
<< poly >>
rect 9 62 11 67
rect 19 62 21 67
rect 39 63 41 68
rect 46 63 48 68
rect 56 63 58 68
rect 66 63 68 68
rect 76 67 78 72
rect 9 39 11 42
rect 19 39 21 46
rect 39 39 41 47
rect 46 39 48 47
rect 56 39 58 47
rect 66 39 68 47
rect 76 39 78 47
rect 5 37 11 39
rect 5 35 7 37
rect 9 35 11 37
rect 5 33 11 35
rect 17 37 23 39
rect 17 35 19 37
rect 21 35 23 37
rect 17 33 23 35
rect 32 37 42 39
rect 32 35 34 37
rect 36 35 42 37
rect 46 36 49 39
rect 32 33 42 35
rect 9 26 11 33
rect 19 23 21 33
rect 40 30 42 33
rect 47 30 49 36
rect 55 37 61 39
rect 55 35 57 37
rect 59 35 61 37
rect 55 33 61 35
rect 65 37 71 39
rect 65 35 67 37
rect 69 35 71 37
rect 65 33 71 35
rect 76 37 86 39
rect 76 35 82 37
rect 84 35 86 37
rect 76 33 86 35
rect 57 30 59 33
rect 67 30 69 33
rect 77 30 79 33
rect 9 11 11 16
rect 19 11 21 16
rect 40 18 42 23
rect 47 14 49 23
rect 57 18 59 23
rect 67 20 69 23
rect 63 18 69 20
rect 63 14 65 18
rect 47 12 65 14
rect 77 15 79 20
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 4 16 9 20
rect 11 23 16 26
rect 32 23 40 30
rect 42 23 47 30
rect 49 28 57 30
rect 49 26 52 28
rect 54 26 57 28
rect 49 23 57 26
rect 59 27 67 30
rect 59 25 62 27
rect 64 25 67 27
rect 59 23 67 25
rect 69 23 77 30
rect 11 20 19 23
rect 11 18 14 20
rect 16 18 19 20
rect 11 16 19 18
rect 21 20 28 23
rect 21 18 24 20
rect 26 18 28 20
rect 21 16 28 18
rect 32 11 38 23
rect 71 20 77 23
rect 79 28 86 30
rect 79 26 82 28
rect 84 26 86 28
rect 79 24 86 26
rect 79 20 84 24
rect 71 16 75 20
rect 69 14 75 16
rect 69 12 71 14
rect 73 12 75 14
rect 32 9 34 11
rect 36 9 38 11
rect 69 10 75 12
rect 32 7 38 9
<< pdif >>
rect 70 63 76 67
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 53 9 58
rect 2 51 4 53
rect 6 51 9 53
rect 2 49 9 51
rect 4 42 9 49
rect 11 60 19 62
rect 11 58 14 60
rect 16 58 19 60
rect 11 46 19 58
rect 21 60 28 62
rect 21 58 24 60
rect 26 58 28 60
rect 21 53 28 58
rect 21 51 24 53
rect 26 51 28 53
rect 21 49 28 51
rect 32 61 39 63
rect 32 59 34 61
rect 36 59 39 61
rect 21 46 26 49
rect 32 47 39 59
rect 41 47 46 63
rect 48 52 56 63
rect 48 50 51 52
rect 53 50 56 52
rect 48 47 56 50
rect 58 61 66 63
rect 58 59 61 61
rect 63 59 66 61
rect 58 47 66 59
rect 68 61 76 63
rect 68 59 71 61
rect 73 59 76 61
rect 68 47 76 59
rect 78 63 83 67
rect 78 61 85 63
rect 78 59 81 61
rect 83 59 85 61
rect 78 54 85 59
rect 78 52 81 54
rect 83 52 85 54
rect 78 50 85 52
rect 78 47 83 50
rect 11 42 17 46
<< alu1 >>
rect -2 81 90 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 90 81
rect -2 68 90 79
rect 50 52 54 55
rect 50 50 51 52
rect 53 50 54 52
rect 50 47 54 50
rect 2 39 6 47
rect 2 37 14 39
rect 2 35 7 37
rect 9 35 14 37
rect 2 33 14 35
rect 42 43 54 47
rect 42 29 46 43
rect 58 39 62 55
rect 50 37 62 39
rect 50 35 57 37
rect 59 35 62 37
rect 50 33 62 35
rect 74 41 86 47
rect 81 37 86 41
rect 81 35 82 37
rect 84 35 86 37
rect 81 33 86 35
rect 42 28 56 29
rect 42 26 52 28
rect 54 26 56 28
rect 42 25 56 26
rect -2 11 90 12
rect -2 9 34 11
rect 36 9 90 11
rect -2 1 90 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 90 1
rect -2 -2 90 -1
<< ptie >>
rect 0 1 88 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 88 1
rect 0 -3 88 -1
<< ntie >>
rect 0 81 88 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 88 81
rect 0 77 88 79
<< nmos >>
rect 9 16 11 26
rect 40 23 42 30
rect 47 23 49 30
rect 57 23 59 30
rect 67 23 69 30
rect 19 16 21 23
rect 77 20 79 30
<< pmos >>
rect 9 42 11 62
rect 19 46 21 62
rect 39 47 41 63
rect 46 47 48 63
rect 56 47 58 63
rect 66 47 68 63
rect 76 47 78 67
<< polyct0 >>
rect 19 35 21 37
rect 34 35 36 37
rect 67 35 69 37
<< polyct1 >>
rect 7 35 9 37
rect 57 35 59 37
rect 82 35 84 37
<< ndifct0 >>
rect 4 22 6 24
rect 62 25 64 27
rect 14 18 16 20
rect 24 18 26 20
rect 82 26 84 28
rect 71 12 73 14
<< ndifct1 >>
rect 52 26 54 28
rect 34 9 36 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
<< pdifct0 >>
rect 4 58 6 60
rect 4 51 6 53
rect 14 58 16 60
rect 24 58 26 60
rect 24 51 26 53
rect 34 59 36 61
rect 61 59 63 61
rect 71 59 73 61
rect 81 59 83 61
rect 81 52 83 54
<< pdifct1 >>
rect 51 50 53 52
<< alu0 >>
rect 2 60 8 61
rect 2 58 4 60
rect 6 58 8 60
rect 2 54 8 58
rect 12 60 18 68
rect 32 61 38 68
rect 12 58 14 60
rect 16 58 18 60
rect 12 57 18 58
rect 22 60 28 61
rect 22 58 24 60
rect 26 58 28 60
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 42 61 65 62
rect 42 59 61 61
rect 63 59 65 61
rect 42 58 65 59
rect 69 61 75 68
rect 69 59 71 61
rect 73 59 75 61
rect 69 58 75 59
rect 80 61 84 63
rect 80 59 81 61
rect 83 59 84 61
rect 22 54 28 58
rect 42 54 46 58
rect 2 53 17 54
rect 2 51 4 53
rect 6 51 17 53
rect 2 50 17 51
rect 22 53 46 54
rect 22 51 24 53
rect 26 51 46 53
rect 22 50 46 51
rect 13 47 17 50
rect 13 43 22 47
rect 18 38 22 43
rect 18 37 38 38
rect 18 35 19 37
rect 21 35 34 37
rect 36 35 38 37
rect 18 34 38 35
rect 18 29 22 34
rect 3 25 22 29
rect 80 54 84 59
rect 66 52 81 54
rect 83 52 84 54
rect 66 50 84 52
rect 66 37 70 50
rect 66 35 67 37
rect 69 35 76 37
rect 66 33 76 35
rect 72 29 76 33
rect 61 27 65 29
rect 61 25 62 27
rect 64 25 65 27
rect 72 28 86 29
rect 72 26 82 28
rect 84 26 86 28
rect 72 25 86 26
rect 3 24 7 25
rect 3 22 4 24
rect 6 22 7 24
rect 3 20 7 22
rect 61 21 65 25
rect 12 20 18 21
rect 12 18 14 20
rect 16 18 18 20
rect 12 12 18 18
rect 22 20 65 21
rect 22 18 24 20
rect 26 18 65 20
rect 22 17 65 18
rect 70 14 74 16
rect 70 12 71 14
rect 73 12 74 14
<< labels >>
rlabel alu0 5 24 5 24 6 an
rlabel alu0 5 55 5 55 6 an
rlabel alu0 9 52 9 52 6 an
rlabel alu0 28 36 28 36 6 an
rlabel alu0 25 55 25 55 6 n1
rlabel alu0 63 23 63 23 6 n3
rlabel alu0 43 19 43 19 6 n3
rlabel alu0 34 52 34 52 6 n1
rlabel alu0 53 60 53 60 6 n1
rlabel alu0 79 27 79 27 6 bn
rlabel alu0 68 43 68 43 6 bn
rlabel alu0 82 56 82 56 6 bn
rlabel alu1 12 36 12 36 6 a
rlabel alu1 4 40 4 40 6 a
rlabel alu1 44 6 44 6 6 vss
rlabel alu1 44 36 44 36 6 z
rlabel alu1 52 36 52 36 6 c
rlabel alu1 60 44 60 44 6 c
rlabel alu1 52 52 52 52 6 z
rlabel alu1 44 74 44 74 6 vdd
rlabel alu1 76 44 76 44 6 b
rlabel alu1 84 40 84 40 6 b
<< end >>
