magic
tech scmos
timestamp 1199202423
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 61 11 65
rect 9 40 11 43
rect 3 38 11 40
rect 3 36 5 38
rect 7 36 11 38
rect 3 34 11 36
rect 9 30 11 34
rect 9 16 11 21
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 21 9 24
rect 11 21 18 30
rect 13 14 18 21
rect 12 11 18 14
rect 12 9 14 11
rect 16 9 18 11
rect 12 7 18 9
<< pdif >>
rect 2 71 8 73
rect 2 69 4 71
rect 6 69 8 71
rect 2 67 8 69
rect 2 61 7 67
rect 2 43 9 61
rect 11 49 16 61
rect 11 47 18 49
rect 11 45 14 47
rect 16 45 18 47
rect 11 43 18 45
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 71 26 79
rect -2 69 4 71
rect 6 69 26 71
rect -2 68 26 69
rect 2 58 15 62
rect 2 39 6 58
rect 13 47 17 49
rect 13 45 14 47
rect 16 45 17 47
rect 2 38 9 39
rect 2 36 5 38
rect 7 36 9 38
rect 2 35 9 36
rect 13 31 17 45
rect 2 28 17 31
rect 2 26 4 28
rect 6 26 17 28
rect 2 25 17 26
rect 2 17 6 25
rect -2 11 26 12
rect -2 9 14 11
rect 16 9 26 11
rect -2 1 26 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 21 11 30
<< pmos >>
rect 9 43 11 61
<< polyct1 >>
rect 5 36 7 38
<< ndifct1 >>
rect 4 26 6 28
rect 14 9 16 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct1 >>
rect 4 69 6 71
rect 14 45 16 47
<< labels >>
rlabel alu1 4 24 4 24 6 z
rlabel alu1 4 48 4 48 6 a
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 12 60 12 60 6 a
<< end >>
