magic
tech scmos
timestamp 1199470087
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 15 94 17 98
rect 23 94 25 98
rect 35 94 37 98
rect 43 94 45 98
rect 15 43 17 55
rect 23 52 25 55
rect 35 52 37 55
rect 23 50 37 52
rect 27 48 29 50
rect 31 48 33 50
rect 27 46 33 48
rect 15 41 23 43
rect 15 39 19 41
rect 21 39 23 41
rect 15 37 23 39
rect 15 34 17 37
rect 27 34 29 46
rect 43 43 45 55
rect 37 41 45 43
rect 37 39 39 41
rect 41 39 45 41
rect 37 37 45 39
rect 15 8 17 13
rect 27 8 29 13
<< ndif >>
rect 6 21 15 34
rect 6 19 9 21
rect 11 19 15 21
rect 6 13 15 19
rect 17 31 27 34
rect 17 29 21 31
rect 23 29 27 31
rect 17 21 27 29
rect 17 19 21 21
rect 23 19 27 21
rect 17 13 27 19
rect 29 31 38 34
rect 29 29 33 31
rect 35 29 38 31
rect 29 21 38 29
rect 29 19 33 21
rect 35 19 38 21
rect 29 13 38 19
<< pdif >>
rect 6 91 15 94
rect 6 89 9 91
rect 11 89 15 91
rect 6 81 15 89
rect 6 79 9 81
rect 11 79 15 81
rect 6 71 15 79
rect 6 69 9 71
rect 11 69 15 71
rect 6 55 15 69
rect 17 55 23 94
rect 25 71 35 94
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 55 43 94
rect 45 91 54 94
rect 45 89 49 91
rect 51 89 54 91
rect 45 81 54 89
rect 45 79 49 81
rect 51 79 54 81
rect 45 71 54 79
rect 45 69 49 71
rect 51 69 54 71
rect 45 55 54 69
<< alu1 >>
rect -2 91 62 100
rect -2 89 9 91
rect 11 89 49 91
rect 51 89 62 91
rect -2 88 62 89
rect 8 81 12 88
rect 8 79 9 81
rect 11 79 12 81
rect 8 71 12 79
rect 48 81 52 88
rect 48 79 49 81
rect 51 79 52 81
rect 8 69 9 71
rect 11 69 12 71
rect 8 67 12 69
rect 27 71 33 72
rect 27 69 29 71
rect 31 69 33 71
rect 27 63 33 69
rect 48 71 52 79
rect 48 69 49 71
rect 51 69 52 71
rect 48 67 52 69
rect 8 61 33 63
rect 8 59 29 61
rect 31 59 33 61
rect 8 58 33 59
rect 8 33 12 58
rect 38 53 42 63
rect 17 42 22 53
rect 27 50 42 53
rect 27 48 29 50
rect 31 48 42 50
rect 27 47 42 48
rect 17 41 43 42
rect 17 39 19 41
rect 21 39 39 41
rect 41 39 43 41
rect 17 38 43 39
rect 8 31 24 33
rect 8 29 21 31
rect 23 29 24 31
rect 8 27 24 29
rect 8 21 12 23
rect 8 19 9 21
rect 11 19 12 21
rect 8 12 12 19
rect 18 21 24 27
rect 18 19 21 21
rect 23 19 24 21
rect 18 17 24 19
rect 32 31 36 33
rect 32 29 33 31
rect 35 29 36 31
rect 32 21 36 29
rect 32 19 33 21
rect 35 19 36 21
rect 32 12 36 19
rect -2 7 62 12
rect -2 5 49 7
rect 51 5 62 7
rect -2 0 62 5
<< ptie >>
rect 47 7 53 37
rect 47 5 49 7
rect 51 5 53 7
rect 47 3 53 5
<< nmos >>
rect 15 13 17 34
rect 27 13 29 34
<< pmos >>
rect 15 55 17 94
rect 23 55 25 94
rect 35 55 37 94
rect 43 55 45 94
<< polyct1 >>
rect 29 48 31 50
rect 19 39 21 41
rect 39 39 41 41
<< ndifct1 >>
rect 9 19 11 21
rect 21 29 23 31
rect 21 19 23 21
rect 33 29 35 31
rect 33 19 35 21
<< ptiect1 >>
rect 49 5 51 7
<< pdifct1 >>
rect 9 89 11 91
rect 9 79 11 81
rect 9 69 11 71
rect 29 69 31 71
rect 29 59 31 61
rect 49 89 51 91
rect 49 79 51 81
rect 49 69 51 71
<< labels >>
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 25 20 25 6 z
rlabel alu1 20 45 20 45 6 a
rlabel alu1 20 60 20 60 6 z
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 30 40 30 40 6 a
rlabel polyct1 40 40 40 40 6 a
rlabel alu1 30 50 30 50 6 b
rlabel alu1 30 65 30 65 6 z
rlabel alu1 40 55 40 55 6 b
rlabel alu1 30 94 30 94 6 vdd
<< end >>
