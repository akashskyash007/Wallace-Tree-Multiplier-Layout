magic
tech scmos
timestamp 1199202882
<< ab >>
rect 0 0 104 80
<< nwell >>
rect -5 36 109 88
<< pwell >>
rect -5 -8 109 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 78 61 80 66
rect 88 61 90 65
rect 9 33 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 50 39 52 42
rect 60 39 62 42
rect 16 37 28 39
rect 22 35 24 37
rect 26 35 28 37
rect 22 33 28 35
rect 32 37 46 39
rect 32 35 42 37
rect 44 35 46 37
rect 32 33 46 35
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 22 30 24 33
rect 32 30 34 33
rect 9 27 15 29
rect 44 22 46 33
rect 50 37 62 39
rect 67 39 69 42
rect 78 39 80 42
rect 88 39 90 42
rect 67 37 73 39
rect 50 29 56 37
rect 67 35 69 37
rect 71 35 73 37
rect 67 33 73 35
rect 78 37 90 39
rect 78 35 85 37
rect 87 35 90 37
rect 78 33 90 35
rect 78 30 80 33
rect 50 27 52 29
rect 54 27 56 29
rect 50 25 56 27
rect 54 22 56 25
rect 22 6 24 11
rect 32 6 34 11
rect 44 6 46 11
rect 54 6 56 11
rect 78 6 80 11
<< ndif >>
rect 17 24 22 30
rect 13 14 22 24
rect 13 12 16 14
rect 18 12 22 14
rect 13 11 22 12
rect 24 21 32 30
rect 24 19 27 21
rect 29 19 32 21
rect 24 11 32 19
rect 34 22 42 30
rect 71 28 78 30
rect 71 26 73 28
rect 75 26 78 28
rect 34 14 44 22
rect 34 12 38 14
rect 40 12 44 14
rect 34 11 44 12
rect 46 20 54 22
rect 46 18 49 20
rect 51 18 54 20
rect 46 11 54 18
rect 56 15 66 22
rect 71 21 78 26
rect 71 19 73 21
rect 75 19 78 21
rect 71 17 78 19
rect 56 13 61 15
rect 63 13 66 15
rect 56 11 66 13
rect 73 11 78 17
rect 80 23 87 30
rect 80 21 83 23
rect 85 21 87 23
rect 80 15 87 21
rect 80 13 83 15
rect 85 13 87 15
rect 80 11 87 13
rect 13 9 20 11
rect 36 9 42 11
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 42 16 70
rect 18 61 26 70
rect 18 59 21 61
rect 23 59 26 61
rect 18 53 26 59
rect 18 51 21 53
rect 23 51 26 53
rect 18 42 26 51
rect 28 42 33 70
rect 35 68 43 70
rect 35 66 38 68
rect 40 66 43 68
rect 35 61 43 66
rect 35 59 38 61
rect 40 59 43 61
rect 35 42 43 59
rect 45 42 50 70
rect 52 53 60 70
rect 52 51 55 53
rect 57 51 60 53
rect 52 46 60 51
rect 52 44 55 46
rect 57 44 60 46
rect 52 42 60 44
rect 62 42 67 70
rect 69 68 76 70
rect 69 66 72 68
rect 74 66 76 68
rect 69 61 76 66
rect 69 59 72 61
rect 74 59 78 61
rect 69 54 78 59
rect 69 52 72 54
rect 74 52 78 54
rect 69 42 78 52
rect 80 53 88 61
rect 80 51 83 53
rect 85 51 88 53
rect 80 46 88 51
rect 80 44 83 46
rect 85 44 88 46
rect 80 42 88 44
rect 90 59 97 61
rect 90 57 93 59
rect 95 57 97 59
rect 90 42 97 57
<< alu1 >>
rect -2 81 106 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 106 81
rect -2 68 106 79
rect 18 61 24 63
rect 18 59 21 61
rect 23 59 24 61
rect 18 54 24 59
rect 2 53 63 54
rect 2 51 21 53
rect 23 51 55 53
rect 57 51 63 53
rect 2 50 63 51
rect 2 22 6 50
rect 90 38 94 47
rect 22 37 31 38
rect 22 35 24 37
rect 26 35 31 37
rect 22 34 31 35
rect 81 37 94 38
rect 81 35 85 37
rect 87 35 94 37
rect 81 34 94 35
rect 25 30 31 34
rect 25 29 63 30
rect 25 27 52 29
rect 54 27 63 29
rect 25 26 63 27
rect 2 21 55 22
rect 2 19 27 21
rect 29 20 55 21
rect 29 19 49 20
rect 2 18 49 19
rect 51 18 55 20
rect 90 25 94 34
rect -2 1 106 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 106 1
rect -2 -2 106 -1
<< ptie >>
rect 0 1 104 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 104 1
rect 0 -3 104 -1
<< ntie >>
rect 0 81 104 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 104 81
rect 0 77 104 79
<< nmos >>
rect 22 11 24 30
rect 32 11 34 30
rect 44 11 46 22
rect 54 11 56 22
rect 78 11 80 30
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 78 42 80 61
rect 88 42 90 61
<< polyct0 >>
rect 42 35 44 37
rect 11 29 13 31
rect 69 35 71 37
<< polyct1 >>
rect 24 35 26 37
rect 85 35 87 37
rect 52 27 54 29
<< ndifct0 >>
rect 16 12 18 14
rect 73 26 75 28
rect 38 12 40 14
rect 73 19 75 21
rect 61 13 63 15
rect 83 21 85 23
rect 83 13 85 15
<< ndifct1 >>
rect 27 19 29 21
rect 49 18 51 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 38 66 40 68
rect 38 59 40 61
rect 55 44 57 46
rect 72 66 74 68
rect 72 59 74 61
rect 72 52 74 54
rect 83 51 85 53
rect 83 44 85 46
rect 93 57 95 59
<< pdifct1 >>
rect 21 59 23 61
rect 21 51 23 53
rect 55 51 57 53
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 36 66 38 68
rect 40 66 42 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 36 61 42 66
rect 36 59 38 61
rect 40 59 42 61
rect 36 58 42 59
rect 71 66 72 68
rect 74 66 75 68
rect 71 61 75 66
rect 71 59 72 61
rect 74 59 75 61
rect 71 54 75 59
rect 92 59 96 68
rect 92 57 93 59
rect 95 57 96 59
rect 92 55 96 57
rect 71 52 72 54
rect 74 52 75 54
rect 71 50 75 52
rect 82 53 86 55
rect 82 51 83 53
rect 85 51 86 53
rect 54 46 58 50
rect 82 46 86 51
rect 14 42 40 46
rect 54 44 55 46
rect 57 44 58 46
rect 54 42 58 44
rect 72 44 83 46
rect 85 44 86 46
rect 72 42 86 44
rect 14 33 18 42
rect 36 38 40 42
rect 72 38 76 42
rect 36 37 76 38
rect 36 35 42 37
rect 44 35 69 37
rect 71 35 76 37
rect 36 34 76 35
rect 10 31 18 33
rect 10 29 11 31
rect 13 29 18 31
rect 10 27 18 29
rect 72 28 76 34
rect 72 26 73 28
rect 75 26 76 28
rect 72 21 76 26
rect 72 19 73 21
rect 75 19 76 21
rect 47 17 53 18
rect 72 17 76 19
rect 82 23 86 25
rect 82 21 83 23
rect 85 21 86 23
rect 60 15 64 17
rect 14 14 20 15
rect 14 12 16 14
rect 18 12 20 14
rect 36 14 42 15
rect 36 12 38 14
rect 40 12 42 14
rect 60 13 61 15
rect 63 13 64 15
rect 60 12 64 13
rect 82 15 86 21
rect 82 13 83 15
rect 85 13 86 15
rect 82 12 86 13
<< labels >>
rlabel alu0 14 30 14 30 6 an
rlabel alu0 56 36 56 36 6 an
rlabel alu0 74 31 74 31 6 an
rlabel alu0 84 48 84 48 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 44 20 44 20 6 z
rlabel ndifct1 28 20 28 20 6 z
rlabel alu1 28 32 28 32 6 b
rlabel alu1 44 28 44 28 6 b
rlabel alu1 36 28 36 28 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 36 52 36 52 6 z
rlabel alu1 52 6 52 6 6 vss
rlabel alu1 52 20 52 20 6 z
rlabel alu1 52 28 52 28 6 b
rlabel alu1 60 28 60 28 6 b
rlabel alu1 52 52 52 52 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 52 74 52 74 6 vdd
rlabel alu1 84 36 84 36 6 a
rlabel alu1 92 36 92 36 6 a
<< end >>
