magic
tech scmos
timestamp 1199203635
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 40 70 42 74
rect 50 70 52 74
rect 40 53 42 56
rect 50 53 52 56
rect 40 51 63 53
rect 41 49 43 51
rect 45 49 47 51
rect 41 47 47 49
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 29 36 33 39
rect 19 33 25 35
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 36
rect 41 30 43 47
rect 51 37 57 39
rect 51 35 53 37
rect 55 35 57 37
rect 51 33 57 35
rect 51 30 53 33
rect 61 30 63 51
rect 12 6 14 11
rect 19 6 21 11
rect 31 8 33 23
rect 61 18 63 23
rect 41 12 43 16
rect 51 8 53 16
rect 31 6 53 8
<< ndif >>
rect 7 23 12 30
rect 5 21 12 23
rect 5 19 7 21
rect 9 19 12 21
rect 5 17 12 19
rect 7 11 12 17
rect 14 11 19 30
rect 21 23 31 30
rect 33 28 41 30
rect 33 26 36 28
rect 38 26 41 28
rect 33 23 41 26
rect 21 11 29 23
rect 23 9 25 11
rect 27 9 29 11
rect 23 7 29 9
rect 36 16 41 23
rect 43 21 51 30
rect 43 19 46 21
rect 48 19 51 21
rect 43 16 51 19
rect 53 28 61 30
rect 53 26 56 28
rect 58 26 61 28
rect 53 23 61 26
rect 63 27 70 30
rect 63 25 66 27
rect 68 25 70 27
rect 63 23 70 25
rect 53 16 58 23
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 57 9 59
rect 4 42 9 57
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 53 29 70
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 68 40 70
rect 31 66 35 68
rect 37 66 40 68
rect 31 56 40 66
rect 42 61 50 70
rect 42 59 45 61
rect 47 59 50 61
rect 42 56 50 59
rect 52 68 59 70
rect 52 66 55 68
rect 57 66 59 68
rect 52 61 59 66
rect 52 59 55 61
rect 57 59 59 61
rect 52 56 59 59
rect 31 42 38 56
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 53 18 54
rect 2 51 14 53
rect 16 51 18 53
rect 2 50 18 51
rect 2 22 6 50
rect 41 51 55 54
rect 41 49 43 51
rect 45 49 55 51
rect 41 48 55 49
rect 49 42 55 48
rect 66 38 70 47
rect 51 37 70 38
rect 51 35 53 37
rect 55 35 70 37
rect 51 33 70 35
rect 2 21 50 22
rect 2 19 7 21
rect 9 19 46 21
rect 48 19 50 21
rect 2 18 50 19
rect -2 11 74 12
rect -2 9 25 11
rect 27 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 12 11 14 30
rect 19 11 21 30
rect 31 23 33 30
rect 41 16 43 30
rect 51 16 53 30
rect 61 23 63 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 40 56 42 70
rect 50 56 52 70
<< polyct0 >>
rect 11 35 13 37
rect 21 35 23 37
<< polyct1 >>
rect 43 49 45 51
rect 53 35 55 37
<< ndifct0 >>
rect 36 26 38 28
rect 56 26 58 28
rect 66 25 68 27
<< ndifct1 >>
rect 7 19 9 21
rect 25 9 27 11
rect 46 19 48 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 59 6 61
rect 24 51 26 53
rect 24 44 26 46
rect 35 66 37 68
rect 45 59 47 61
rect 55 66 57 68
rect 55 59 57 61
<< pdifct1 >>
rect 14 51 16 53
<< alu0 >>
rect 33 66 35 68
rect 37 66 39 68
rect 33 65 39 66
rect 53 66 55 68
rect 57 66 59 68
rect 2 61 49 62
rect 2 59 4 61
rect 6 59 45 61
rect 47 59 49 61
rect 2 58 49 59
rect 53 61 59 66
rect 53 59 55 61
rect 57 59 59 61
rect 53 58 59 59
rect 23 53 27 55
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 10 44 24 46
rect 26 44 27 46
rect 10 42 27 44
rect 10 37 14 42
rect 31 38 35 58
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 19 37 48 38
rect 19 35 21 37
rect 23 35 48 37
rect 19 34 48 35
rect 10 28 40 30
rect 10 26 36 28
rect 38 26 40 28
rect 34 25 40 26
rect 44 29 48 34
rect 44 28 60 29
rect 44 26 56 28
rect 58 26 60 28
rect 44 25 60 26
rect 65 27 69 29
rect 65 25 66 27
rect 68 25 69 27
rect 65 12 69 25
<< labels >>
rlabel polyct0 12 36 12 36 6 bn
rlabel alu0 25 48 25 48 6 bn
rlabel alu0 33 36 33 36 6 an
rlabel alu0 25 28 25 28 6 bn
rlabel alu0 25 60 25 60 6 an
rlabel alu0 52 27 52 27 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 44 52 44 52 6 a
rlabel alu1 52 48 52 48 6 a
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 36 60 36 6 b
rlabel alu1 68 40 68 40 6 b
<< end >>
