magic
tech scmos
timestamp 1199201646
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 39 11 42
rect 19 39 21 51
rect 29 47 31 51
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 30 11 33
rect 22 30 24 33
rect 29 30 31 41
rect 9 11 11 16
rect 22 12 24 17
rect 29 12 31 17
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 20 9 26
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 17 22 30
rect 24 17 29 30
rect 31 23 36 30
rect 31 21 38 23
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
rect 11 16 20 17
rect 13 11 20 16
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 51 19 59
rect 21 62 29 70
rect 21 60 24 62
rect 26 60 29 62
rect 21 55 29 60
rect 21 53 24 55
rect 26 53 29 55
rect 21 51 29 53
rect 31 68 38 70
rect 31 66 34 68
rect 36 66 38 68
rect 31 61 38 66
rect 31 59 34 61
rect 36 59 38 61
rect 31 51 38 59
rect 11 42 17 51
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 61 7 63
rect 2 59 4 61
rect 6 59 7 61
rect 2 54 7 59
rect 2 52 4 54
rect 6 52 7 54
rect 2 50 7 52
rect 2 28 6 50
rect 34 46 38 55
rect 25 45 38 46
rect 25 43 31 45
rect 33 43 38 45
rect 25 42 38 43
rect 17 37 31 38
rect 17 35 21 37
rect 23 35 31 37
rect 17 34 31 35
rect 2 26 4 28
rect 2 23 6 26
rect 2 20 14 23
rect 2 18 4 20
rect 6 18 14 20
rect 26 25 31 34
rect 2 17 14 18
rect -2 11 42 12
rect -2 9 15 11
rect 17 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 16 11 30
rect 22 17 24 30
rect 29 17 31 30
<< pmos >>
rect 9 42 11 70
rect 19 51 21 70
rect 29 51 31 70
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 31 43 33 45
rect 21 35 23 37
<< ndifct0 >>
rect 34 19 36 21
<< ndifct1 >>
rect 4 26 6 28
rect 4 18 6 20
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 66 16 68
rect 14 59 16 61
rect 24 60 26 62
rect 24 53 26 55
rect 34 66 36 68
rect 34 59 36 61
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 61 18 66
rect 32 66 34 68
rect 36 66 38 68
rect 12 59 14 61
rect 16 59 18 61
rect 12 58 18 59
rect 22 62 28 63
rect 22 60 24 62
rect 26 60 28 62
rect 22 55 28 60
rect 32 61 38 66
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 22 54 24 55
rect 14 53 24 54
rect 26 53 28 55
rect 14 50 28 53
rect 14 46 18 50
rect 10 42 18 46
rect 10 37 14 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 6 23 7 30
rect 10 26 22 30
rect 18 22 22 26
rect 18 21 38 22
rect 18 19 34 21
rect 36 19 38 21
rect 18 18 38 19
<< labels >>
rlabel polyct0 12 36 12 36 6 zn
rlabel alu0 25 56 25 56 6 zn
rlabel alu0 28 20 28 20 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 52 36 52 6 b
<< end >>
