magic
tech scmos
timestamp 1199202894
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 12 63 14 68
rect 19 63 21 68
rect 33 60 35 65
rect 12 42 14 48
rect 9 40 15 42
rect 9 38 11 40
rect 13 38 15 40
rect 9 36 15 38
rect 11 22 13 36
rect 19 31 21 48
rect 33 42 35 48
rect 25 40 35 42
rect 25 38 27 40
rect 29 38 35 40
rect 25 36 35 38
rect 17 29 23 31
rect 33 30 35 36
rect 17 27 19 29
rect 21 27 23 29
rect 17 25 23 27
rect 21 22 23 25
rect 33 19 35 24
rect 11 9 13 14
rect 21 9 23 14
<< ndif >>
rect 25 24 33 30
rect 35 28 42 30
rect 35 26 38 28
rect 40 26 42 28
rect 35 24 42 26
rect 25 22 31 24
rect 3 14 11 22
rect 13 20 21 22
rect 13 18 16 20
rect 18 18 21 20
rect 13 14 21 18
rect 23 19 31 22
rect 23 17 27 19
rect 29 17 31 19
rect 23 14 31 17
rect 3 11 9 14
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
<< pdif >>
rect 5 61 12 63
rect 5 59 7 61
rect 9 59 12 61
rect 5 57 12 59
rect 7 48 12 57
rect 14 48 19 63
rect 21 61 31 63
rect 21 59 27 61
rect 29 60 31 61
rect 29 59 33 60
rect 21 54 33 59
rect 21 52 28 54
rect 30 52 33 54
rect 21 48 33 52
rect 35 54 40 60
rect 35 52 42 54
rect 35 50 38 52
rect 40 50 42 52
rect 35 48 42 50
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 2 61 14 63
rect 2 59 7 61
rect 9 59 14 61
rect 2 57 14 59
rect 2 22 6 57
rect 18 47 22 55
rect 10 43 22 47
rect 10 40 14 43
rect 10 38 11 40
rect 13 38 14 40
rect 26 40 30 47
rect 26 39 27 40
rect 10 33 14 38
rect 18 38 27 39
rect 29 38 30 40
rect 18 33 30 38
rect 2 20 23 22
rect 2 18 16 20
rect 18 18 23 20
rect 2 17 23 18
rect -2 11 50 12
rect -2 9 5 11
rect 7 9 50 11
rect -2 1 50 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 33 24 35 30
rect 11 14 13 22
rect 21 14 23 22
<< pmos >>
rect 12 48 14 63
rect 19 48 21 63
rect 33 48 35 60
<< polyct0 >>
rect 19 27 21 29
<< polyct1 >>
rect 11 38 13 40
rect 27 38 29 40
<< ndifct0 >>
rect 38 26 40 28
rect 27 17 29 19
<< ndifct1 >>
rect 16 18 18 20
rect 5 9 7 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 27 59 29 61
rect 28 52 30 54
rect 38 50 40 52
<< pdifct1 >>
rect 7 59 9 61
<< alu0 >>
rect 26 61 32 68
rect 26 59 27 61
rect 29 59 32 61
rect 26 54 32 59
rect 26 52 28 54
rect 30 52 32 54
rect 26 51 32 52
rect 37 52 41 54
rect 37 50 38 52
rect 40 50 41 52
rect 37 30 41 50
rect 17 29 41 30
rect 17 27 19 29
rect 21 28 41 29
rect 21 27 38 28
rect 17 26 38 27
rect 40 26 41 28
rect 37 24 41 26
rect 26 19 30 21
rect 26 17 27 19
rect 29 17 30 19
rect 26 12 30 17
<< labels >>
rlabel alu0 29 28 29 28 6 an
rlabel alu0 39 39 39 39 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 36 20 36 6 a
rlabel alu1 12 40 12 40 6 b
rlabel alu1 20 52 20 52 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 40 28 40 6 a
rlabel alu1 24 74 24 74 6 vdd
<< end >>
