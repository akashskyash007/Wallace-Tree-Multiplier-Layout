magic
tech scmos
timestamp 1199202450
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 10 66 12 70
rect 18 66 20 70
rect 28 66 30 70
rect 36 66 38 70
rect 48 58 54 60
rect 48 56 50 58
rect 52 56 54 58
rect 45 54 54 56
rect 45 51 47 54
rect 10 38 12 41
rect 18 38 20 41
rect 28 38 30 41
rect 36 38 38 41
rect 45 39 47 42
rect 9 35 12 38
rect 16 36 22 38
rect 9 27 11 35
rect 16 34 18 36
rect 20 34 22 36
rect 16 32 22 34
rect 26 36 32 38
rect 36 36 40 38
rect 45 37 50 39
rect 26 34 28 36
rect 30 34 32 36
rect 26 32 32 34
rect 38 33 40 36
rect 26 28 28 32
rect 38 31 44 33
rect 38 29 40 31
rect 42 29 44 31
rect 38 28 44 29
rect 2 25 11 27
rect 2 23 4 25
rect 6 23 11 25
rect 2 21 11 23
rect 9 18 11 21
rect 16 26 28 28
rect 35 27 44 28
rect 35 26 41 27
rect 16 18 18 26
rect 35 23 37 26
rect 48 23 50 37
rect 26 18 28 22
rect 45 21 50 23
rect 45 18 47 21
rect 35 8 37 12
rect 9 2 11 6
rect 16 2 18 6
rect 26 4 28 7
rect 45 4 47 12
rect 26 2 47 4
<< ndif >>
rect 30 18 35 23
rect 2 10 9 18
rect 2 8 4 10
rect 6 8 9 10
rect 2 6 9 8
rect 11 6 16 18
rect 18 16 26 18
rect 18 14 21 16
rect 23 14 26 16
rect 18 7 26 14
rect 28 12 35 18
rect 37 18 42 23
rect 37 16 45 18
rect 37 14 40 16
rect 42 14 45 16
rect 37 12 45 14
rect 47 16 54 18
rect 47 14 50 16
rect 52 14 54 16
rect 47 12 54 14
rect 28 7 33 12
rect 18 6 23 7
<< pdif >>
rect 2 64 10 66
rect 2 62 4 64
rect 6 62 10 64
rect 2 57 10 62
rect 2 55 4 57
rect 6 55 10 57
rect 2 41 10 55
rect 12 41 18 66
rect 20 57 28 66
rect 20 55 23 57
rect 25 55 28 57
rect 20 41 28 55
rect 30 41 36 66
rect 38 64 45 66
rect 38 62 41 64
rect 43 62 45 64
rect 38 59 45 62
rect 38 51 43 59
rect 38 42 45 51
rect 47 49 54 51
rect 47 47 50 49
rect 52 47 54 49
rect 47 45 54 47
rect 47 42 52 45
rect 38 41 43 42
<< alu1 >>
rect -2 64 58 72
rect 10 57 27 59
rect 48 58 54 59
rect 10 55 23 57
rect 25 55 27 57
rect 10 54 27 55
rect 32 56 50 58
rect 52 56 54 58
rect 32 54 54 56
rect 10 28 14 54
rect 32 50 36 54
rect 18 46 36 50
rect 18 36 22 46
rect 20 34 22 36
rect 18 32 22 34
rect 50 34 54 43
rect 2 25 6 27
rect 2 23 4 25
rect 2 18 6 23
rect 10 24 23 28
rect 2 14 15 18
rect 19 17 23 24
rect 38 31 54 34
rect 38 29 40 31
rect 42 29 54 31
rect 38 28 54 29
rect 19 16 25 17
rect 19 14 21 16
rect 23 14 25 16
rect 19 13 25 14
rect -2 0 58 8
<< nmos >>
rect 9 6 11 18
rect 16 6 18 18
rect 26 7 28 18
rect 35 12 37 23
rect 45 12 47 18
<< pmos >>
rect 10 41 12 66
rect 18 41 20 66
rect 28 41 30 66
rect 36 41 38 66
rect 45 42 47 51
<< polyct0 >>
rect 28 34 30 36
<< polyct1 >>
rect 50 56 52 58
rect 18 34 20 36
rect 40 29 42 31
rect 4 23 6 25
<< ndifct0 >>
rect 4 8 6 10
rect 40 14 42 16
rect 50 14 52 16
<< ndifct1 >>
rect 21 14 23 16
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 41 62 43 64
rect 50 47 52 49
<< pdifct1 >>
rect 23 55 25 57
<< alu0 >>
rect 3 62 4 64
rect 6 62 7 64
rect 3 57 7 62
rect 39 62 41 64
rect 43 62 45 64
rect 39 61 45 62
rect 3 55 4 57
rect 6 55 7 57
rect 3 53 7 55
rect 42 49 54 50
rect 42 47 50 49
rect 52 47 54 49
rect 42 46 54 47
rect 17 32 18 38
rect 42 42 46 46
rect 30 38 46 42
rect 30 37 34 38
rect 26 36 34 37
rect 26 34 28 36
rect 30 34 34 36
rect 26 33 34 34
rect 6 18 7 27
rect 30 24 34 33
rect 30 20 54 24
rect 38 16 44 17
rect 38 14 40 16
rect 42 14 44 16
rect 2 10 8 11
rect 2 8 4 10
rect 6 8 8 10
rect 38 8 44 14
rect 48 16 54 20
rect 48 14 50 16
rect 52 14 54 16
rect 48 13 54 14
<< labels >>
rlabel alu0 32 31 32 31 6 sn
rlabel alu0 51 18 51 18 6 sn
rlabel alu0 48 48 48 48 6 sn
rlabel alu1 4 24 4 24 6 a0
rlabel alu1 12 16 12 16 6 a0
rlabel alu1 20 40 20 40 6 s
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 48 28 48 6 s
rlabel alu1 36 56 36 56 6 s
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 52 36 52 36 6 a1
rlabel alu1 44 56 44 56 6 s
<< end >>
