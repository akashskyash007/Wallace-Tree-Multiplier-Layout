magic
tech scmos
timestamp 1199469104
<< ab >>
rect 0 0 110 100
<< nwell >>
rect -5 48 115 105
<< pwell >>
rect -5 -5 115 48
<< poly >>
rect 11 93 13 98
rect 23 93 25 98
rect 35 93 37 98
rect 47 93 49 98
rect 59 93 61 98
rect 71 93 73 98
rect 83 93 85 98
rect 95 93 97 98
rect 11 47 13 56
rect 23 53 25 56
rect 35 53 37 56
rect 47 53 49 56
rect 59 53 61 56
rect 71 53 73 56
rect 83 53 85 56
rect 95 53 97 56
rect 23 51 41 53
rect 35 49 37 51
rect 39 49 41 51
rect 35 47 41 49
rect 11 45 23 47
rect 17 43 19 45
rect 21 43 23 45
rect 17 41 23 43
rect 39 39 41 47
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 57 51 63 53
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 67 51 85 53
rect 91 51 97 53
rect 67 49 70 51
rect 72 49 74 51
rect 67 47 74 49
rect 91 49 93 51
rect 95 49 97 51
rect 91 47 97 49
rect 47 39 49 47
rect 59 39 61 47
rect 67 39 69 47
rect 39 2 41 6
rect 47 2 49 6
rect 59 2 61 6
rect 67 2 69 6
<< ndif >>
rect 30 11 39 39
rect 30 9 33 11
rect 35 9 39 11
rect 30 6 39 9
rect 41 6 47 39
rect 49 31 59 39
rect 49 29 53 31
rect 55 29 59 31
rect 49 21 59 29
rect 49 19 53 21
rect 55 19 59 21
rect 49 6 59 19
rect 61 6 67 39
rect 69 21 78 39
rect 69 19 73 21
rect 75 19 78 21
rect 69 11 78 19
rect 69 9 73 11
rect 75 9 78 11
rect 69 6 78 9
<< pdif >>
rect 6 83 11 93
rect 3 81 11 83
rect 3 79 5 81
rect 7 79 11 81
rect 3 77 11 79
rect 6 56 11 77
rect 13 71 23 93
rect 13 69 17 71
rect 19 69 23 71
rect 13 56 23 69
rect 25 81 35 93
rect 25 79 29 81
rect 31 79 35 81
rect 25 56 35 79
rect 37 71 47 93
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 49 81 59 93
rect 49 79 53 81
rect 55 79 59 81
rect 49 71 59 79
rect 49 69 53 71
rect 55 69 59 71
rect 49 56 59 69
rect 61 91 71 93
rect 61 89 65 91
rect 67 89 71 91
rect 61 81 71 89
rect 61 79 65 81
rect 67 79 71 81
rect 61 56 71 79
rect 73 81 83 93
rect 73 79 77 81
rect 79 79 83 81
rect 73 71 83 79
rect 73 69 77 71
rect 79 69 83 71
rect 73 56 83 69
rect 85 91 95 93
rect 85 89 89 91
rect 91 89 95 91
rect 85 81 95 89
rect 85 79 89 81
rect 91 79 95 81
rect 85 56 95 79
rect 97 70 102 93
rect 97 68 105 70
rect 97 66 101 68
rect 103 66 105 68
rect 97 60 105 66
rect 97 58 101 60
rect 103 58 105 60
rect 97 56 105 58
<< alu1 >>
rect -2 91 112 100
rect -2 89 65 91
rect 67 89 89 91
rect 91 89 112 91
rect -2 88 112 89
rect 3 81 57 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 79 53 81
rect 55 79 57 81
rect 3 78 57 79
rect 8 71 45 73
rect 8 69 17 71
rect 19 69 41 71
rect 43 69 45 71
rect 8 68 45 69
rect 51 72 57 78
rect 64 81 68 88
rect 64 79 65 81
rect 67 79 68 81
rect 64 77 68 79
rect 76 81 80 83
rect 76 79 77 81
rect 79 79 80 81
rect 76 72 80 79
rect 88 81 92 88
rect 88 79 89 81
rect 91 79 92 81
rect 88 77 92 79
rect 51 71 104 72
rect 51 69 53 71
rect 55 69 77 71
rect 79 69 104 71
rect 51 68 104 69
rect 8 22 12 68
rect 100 66 101 68
rect 103 66 104 68
rect 17 58 53 62
rect 17 45 23 58
rect 27 51 42 53
rect 27 49 37 51
rect 39 49 42 51
rect 27 48 42 49
rect 47 51 53 58
rect 47 49 49 51
rect 51 49 53 51
rect 47 48 53 49
rect 57 58 93 62
rect 57 51 63 58
rect 57 49 59 51
rect 61 49 63 51
rect 57 48 63 49
rect 68 51 83 53
rect 68 49 70 51
rect 72 49 83 51
rect 68 48 83 49
rect 87 52 93 58
rect 100 60 104 66
rect 100 58 101 60
rect 103 58 104 60
rect 100 56 104 58
rect 87 51 103 52
rect 87 49 93 51
rect 95 49 103 51
rect 87 48 103 49
rect 17 43 19 45
rect 21 43 23 45
rect 17 38 23 43
rect 38 27 42 48
rect 52 31 56 33
rect 52 29 53 31
rect 55 29 56 31
rect 52 22 56 29
rect 68 27 72 48
rect 87 38 93 48
rect 8 21 56 22
rect 8 19 53 21
rect 55 19 56 21
rect 8 17 56 19
rect 72 21 76 23
rect 72 19 73 21
rect 75 19 76 21
rect 72 12 76 19
rect -2 11 112 12
rect -2 9 33 11
rect 35 9 73 11
rect 75 9 112 11
rect -2 7 112 9
rect -2 5 89 7
rect 91 5 99 7
rect 101 5 112 7
rect -2 0 112 5
<< ptie >>
rect 87 7 103 9
rect 87 5 89 7
rect 91 5 99 7
rect 101 5 103 7
rect 87 3 103 5
<< nmos >>
rect 39 6 41 39
rect 47 6 49 39
rect 59 6 61 39
rect 67 6 69 39
<< pmos >>
rect 11 56 13 93
rect 23 56 25 93
rect 35 56 37 93
rect 47 56 49 93
rect 59 56 61 93
rect 71 56 73 93
rect 83 56 85 93
rect 95 56 97 93
<< polyct1 >>
rect 37 49 39 51
rect 19 43 21 45
rect 49 49 51 51
rect 59 49 61 51
rect 70 49 72 51
rect 93 49 95 51
<< ndifct1 >>
rect 33 9 35 11
rect 53 29 55 31
rect 53 19 55 21
rect 73 19 75 21
rect 73 9 75 11
<< ptiect1 >>
rect 89 5 91 7
rect 99 5 101 7
<< pdifct1 >>
rect 5 79 7 81
rect 17 69 19 71
rect 29 79 31 81
rect 41 69 43 71
rect 53 79 55 81
rect 53 69 55 71
rect 65 89 67 91
rect 65 79 67 81
rect 77 79 79 81
rect 77 69 79 71
rect 89 89 91 91
rect 89 79 91 81
rect 101 66 103 68
rect 101 58 103 60
<< labels >>
rlabel pdifct1 6 80 6 80 6 n3
rlabel pdifct1 30 80 30 80 6 n3
rlabel pdifct1 54 70 54 70 6 n3
rlabel pdifct1 54 80 54 80 6 n3
rlabel pdifct1 102 67 102 67 6 n3
rlabel pdifct1 102 59 102 59 6 n3
rlabel pdifct1 78 70 78 70 6 n3
rlabel pdifct1 78 80 78 80 6 n3
rlabel alu1 10 45 10 45 6 z
rlabel alu1 40 20 40 20 6 z
rlabel alu1 30 20 30 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 40 40 40 40 6 b1
rlabel alu1 20 50 20 50 6 b2
rlabel alu1 30 50 30 50 6 b1
rlabel alu1 40 60 40 60 6 b2
rlabel alu1 30 60 30 60 6 b2
rlabel alu1 20 70 20 70 6 z
rlabel alu1 40 70 40 70 6 z
rlabel alu1 30 70 30 70 6 z
rlabel alu1 55 6 55 6 6 vss
rlabel alu1 50 20 50 20 6 z
rlabel alu1 50 55 50 55 6 b2
rlabel alu1 60 55 60 55 6 a2
rlabel alu1 55 94 55 94 6 vdd
rlabel alu1 70 40 70 40 6 a1
rlabel alu1 80 50 80 50 6 a1
rlabel alu1 80 60 80 60 6 a2
rlabel alu1 70 60 70 60 6 a2
rlabel alu1 90 50 90 50 6 a2
rlabel alu1 100 50 100 50 6 a2
<< end >>
