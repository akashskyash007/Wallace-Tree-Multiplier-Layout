magic
tech scmos
timestamp 1199203108
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 12 70 14 74
rect 22 70 24 74
rect 29 70 31 74
rect 12 50 14 56
rect 9 48 15 50
rect 9 46 11 48
rect 13 46 15 48
rect 9 44 15 46
rect 9 22 11 44
rect 22 40 24 43
rect 17 38 24 40
rect 17 36 19 38
rect 21 36 24 38
rect 17 34 24 36
rect 29 39 31 43
rect 29 37 38 39
rect 29 35 34 37
rect 36 35 38 37
rect 19 22 21 34
rect 29 33 38 35
rect 29 22 31 33
rect 9 6 11 10
rect 19 6 21 10
rect 29 6 31 10
<< ndif >>
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 4 10 9 16
rect 11 20 19 22
rect 11 18 14 20
rect 16 18 19 20
rect 11 10 19 18
rect 21 14 29 22
rect 21 12 24 14
rect 26 12 29 14
rect 21 10 29 12
rect 31 20 38 22
rect 31 18 34 20
rect 36 18 38 20
rect 31 16 38 18
rect 31 10 36 16
<< pdif >>
rect 4 68 12 70
rect 4 66 7 68
rect 9 66 12 68
rect 4 56 12 66
rect 14 61 22 70
rect 14 59 17 61
rect 19 59 22 61
rect 14 56 22 59
rect 17 43 22 56
rect 24 43 29 70
rect 31 68 38 70
rect 31 66 34 68
rect 36 66 38 68
rect 31 61 38 66
rect 31 59 34 61
rect 36 59 38 61
rect 31 43 38 59
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 61 23 62
rect 2 59 17 61
rect 19 59 23 61
rect 2 58 23 59
rect 2 22 6 58
rect 10 48 14 50
rect 10 46 11 48
rect 13 46 14 48
rect 25 47 31 54
rect 10 30 14 46
rect 18 42 31 47
rect 25 37 38 38
rect 25 35 34 37
rect 36 35 38 37
rect 25 34 38 35
rect 10 26 23 30
rect 34 25 38 34
rect 2 20 8 22
rect 2 18 4 20
rect 6 18 8 20
rect 2 17 8 18
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 10 11 22
rect 19 10 21 22
rect 29 10 31 22
<< pmos >>
rect 12 56 14 70
rect 22 43 24 70
rect 29 43 31 70
<< polyct0 >>
rect 19 36 21 38
<< polyct1 >>
rect 11 46 13 48
rect 34 35 36 37
<< ndifct0 >>
rect 14 18 16 20
rect 24 12 26 14
rect 34 18 36 20
<< ndifct1 >>
rect 4 18 6 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 7 66 9 68
rect 34 66 36 68
rect 34 59 36 61
<< pdifct1 >>
rect 17 59 19 61
<< alu0 >>
rect 5 66 7 68
rect 9 66 11 68
rect 5 65 11 66
rect 32 66 34 68
rect 36 66 38 68
rect 32 61 38 66
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 18 38 22 42
rect 18 36 19 38
rect 21 36 22 38
rect 18 34 22 36
rect 12 20 38 22
rect 12 18 14 20
rect 16 18 34 20
rect 36 18 38 20
rect 12 17 18 18
rect 32 17 38 18
rect 22 14 28 15
rect 22 12 24 14
rect 26 12 28 14
<< labels >>
rlabel alu0 25 20 25 20 6 n1
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 28 20 28 6 b
rlabel alu1 28 36 28 36 6 a1
rlabel alu1 20 44 20 44 6 a2
rlabel alu1 28 48 28 48 6 a2
rlabel alu1 20 60 20 60 6 z
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 28 36 28 6 a1
<< end >>
