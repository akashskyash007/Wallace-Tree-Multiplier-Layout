magic
tech scmos
timestamp 1199201850
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 51 66 53 70
rect 61 66 63 70
rect 9 36 11 39
rect 9 34 15 36
rect 9 32 11 34
rect 13 32 15 34
rect 9 30 15 32
rect 19 35 21 39
rect 29 35 31 39
rect 19 33 31 35
rect 39 36 41 39
rect 51 36 53 39
rect 61 36 63 39
rect 39 34 54 36
rect 19 31 27 33
rect 29 31 31 33
rect 19 29 31 31
rect 41 33 54 34
rect 41 31 43 33
rect 45 31 54 33
rect 20 25 22 29
rect 35 25 37 30
rect 41 29 54 31
rect 58 34 64 36
rect 58 32 60 34
rect 62 32 64 34
rect 58 30 64 32
rect 42 25 44 29
rect 52 25 54 29
rect 59 25 61 30
rect 20 5 22 10
rect 35 4 37 12
rect 42 8 44 12
rect 52 8 54 12
rect 59 4 61 12
rect 35 2 61 4
<< ndif >>
rect 15 19 20 25
rect 13 17 20 19
rect 13 15 15 17
rect 17 15 20 17
rect 13 13 20 15
rect 15 10 20 13
rect 22 12 35 25
rect 37 12 42 25
rect 44 17 52 25
rect 44 15 47 17
rect 49 15 52 17
rect 44 12 52 15
rect 54 12 59 25
rect 61 12 69 25
rect 22 10 33 12
rect 24 8 27 10
rect 29 8 33 10
rect 24 6 33 8
rect 63 7 69 12
rect 63 5 65 7
rect 67 5 69 7
rect 63 3 69 5
<< pdif >>
rect 43 67 49 69
rect 43 66 45 67
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 39 9 55
rect 11 58 19 66
rect 11 56 14 58
rect 16 56 19 58
rect 11 39 19 56
rect 21 49 29 66
rect 21 47 24 49
rect 26 47 29 49
rect 21 39 29 47
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 50 39 55
rect 31 48 34 50
rect 36 48 39 50
rect 31 39 39 48
rect 41 65 45 66
rect 47 66 49 67
rect 47 65 51 66
rect 41 39 51 65
rect 53 57 61 66
rect 53 55 56 57
rect 58 55 61 57
rect 53 50 61 55
rect 53 48 56 50
rect 58 48 61 50
rect 53 39 61 48
rect 63 64 70 66
rect 63 62 66 64
rect 68 62 70 64
rect 63 56 70 62
rect 63 54 66 56
rect 68 54 70 56
rect 63 39 70 54
<< alu1 >>
rect -2 67 74 72
rect -2 65 45 67
rect 47 65 74 67
rect -2 64 74 65
rect 2 49 28 51
rect 2 47 24 49
rect 26 47 28 49
rect 2 46 28 47
rect 2 18 6 46
rect 42 42 46 51
rect 10 38 63 42
rect 10 34 14 38
rect 57 34 63 38
rect 10 32 11 34
rect 13 32 14 34
rect 10 30 14 32
rect 25 33 31 34
rect 25 31 27 33
rect 29 31 31 33
rect 25 26 31 31
rect 17 22 31 26
rect 41 33 47 34
rect 41 31 43 33
rect 45 31 47 33
rect 41 26 47 31
rect 57 32 60 34
rect 62 32 63 34
rect 57 30 63 32
rect 41 22 55 26
rect 2 17 55 18
rect 2 15 15 17
rect 17 15 47 17
rect 49 15 55 17
rect 2 14 55 15
rect -2 7 74 8
rect -2 5 5 7
rect 7 5 65 7
rect 67 5 74 7
rect -2 0 74 5
<< ptie >>
rect 3 7 9 24
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< nmos >>
rect 20 10 22 25
rect 35 12 37 25
rect 42 12 44 25
rect 52 12 54 25
rect 59 12 61 25
<< pmos >>
rect 9 39 11 66
rect 19 39 21 66
rect 29 39 31 66
rect 39 39 41 66
rect 51 39 53 66
rect 61 39 63 66
<< polyct1 >>
rect 11 32 13 34
rect 27 31 29 33
rect 43 31 45 33
rect 60 32 62 34
<< ndifct0 >>
rect 27 8 29 10
<< ndifct1 >>
rect 15 15 17 17
rect 47 15 49 17
rect 65 5 67 7
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 56 16 58
rect 34 55 36 57
rect 34 48 36 50
rect 56 55 58 57
rect 56 48 58 50
rect 66 62 68 64
rect 66 54 68 56
<< pdifct1 >>
rect 24 47 26 49
rect 45 65 47 67
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 65 62 66 64
rect 68 62 69 64
rect 2 55 4 57
rect 6 55 8 57
rect 12 58 59 59
rect 12 56 14 58
rect 16 57 59 58
rect 16 56 34 57
rect 12 55 34 56
rect 36 55 56 57
rect 58 55 59 57
rect 2 54 8 55
rect 33 50 37 55
rect 33 48 34 50
rect 36 48 37 50
rect 33 46 37 48
rect 55 50 59 55
rect 65 56 69 62
rect 65 54 66 56
rect 68 54 69 56
rect 65 52 69 54
rect 55 48 56 50
rect 58 48 59 50
rect 55 46 59 48
rect 25 10 31 11
rect 25 8 27 10
rect 29 8 31 10
<< labels >>
rlabel alu0 35 52 35 52 6 n1
rlabel alu0 57 52 57 52 6 n1
rlabel alu0 35 57 35 57 6 n1
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 24 20 24 6 b
rlabel alu1 28 28 28 28 6 b
rlabel alu1 28 40 28 40 6 a1
rlabel alu1 20 40 20 40 6 a1
rlabel alu1 20 48 20 48 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 52 24 52 24 6 a2
rlabel alu1 52 40 52 40 6 a1
rlabel alu1 36 40 36 40 6 a1
rlabel alu1 44 44 44 44 6 a1
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 36 60 36 6 a1
<< end >>
