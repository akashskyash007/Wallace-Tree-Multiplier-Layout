magic
tech scmos
timestamp 1199980706
<< ab >>
rect 0 0 32 88
<< nwell >>
rect -8 40 40 97
<< pwell >>
rect -8 -9 40 40
<< poly >>
rect 5 80 14 86
rect 18 80 27 86
rect 9 77 11 80
rect 21 77 23 80
rect 9 48 11 51
rect 21 48 23 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 46 30 48
rect 15 44 17 46
rect 19 44 30 46
rect 15 42 30 44
rect 2 36 17 38
rect 2 34 13 36
rect 15 34 17 36
rect 2 32 17 34
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 9 29 11 32
rect 21 29 23 32
rect 9 8 11 11
rect 21 8 23 11
rect 5 2 14 8
rect 18 2 27 8
<< ndif >>
rect 2 22 9 29
rect 2 20 4 22
rect 6 20 9 22
rect 2 15 9 20
rect 2 13 4 15
rect 6 13 9 15
rect 2 11 9 13
rect 11 24 21 29
rect 11 22 15 24
rect 17 22 21 24
rect 11 17 21 22
rect 11 15 15 17
rect 17 15 21 17
rect 11 11 21 15
rect 23 15 30 29
rect 23 13 26 15
rect 28 13 30 15
rect 23 11 30 13
<< pdif >>
rect 2 74 9 77
rect 2 72 4 74
rect 6 72 9 74
rect 2 67 9 72
rect 2 65 4 67
rect 6 65 9 67
rect 2 51 9 65
rect 11 73 21 77
rect 11 71 15 73
rect 17 71 21 73
rect 11 65 21 71
rect 11 63 15 65
rect 17 63 21 65
rect 11 57 21 63
rect 11 55 15 57
rect 17 55 21 57
rect 11 51 21 55
rect 23 74 30 77
rect 23 72 26 74
rect 28 72 30 74
rect 23 67 30 72
rect 23 65 26 67
rect 28 65 30 67
rect 23 51 30 65
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 81 34 83
rect 3 74 7 81
rect 3 72 4 74
rect 6 72 7 74
rect 3 67 7 72
rect 3 65 4 67
rect 6 65 7 67
rect 3 63 7 65
rect 14 73 18 75
rect 14 71 15 73
rect 17 71 18 73
rect 14 65 18 71
rect 14 63 15 65
rect 17 63 18 65
rect 25 74 29 81
rect 25 72 26 74
rect 28 72 29 74
rect 25 67 29 72
rect 25 65 26 67
rect 28 65 29 67
rect 25 63 29 65
rect 14 58 18 63
rect 5 57 30 58
rect 5 55 15 57
rect 17 55 30 57
rect 5 54 30 55
rect 26 37 30 54
rect 11 36 30 37
rect 11 34 13 36
rect 15 34 23 36
rect 25 34 30 36
rect 11 33 30 34
rect 2 22 8 23
rect 2 20 4 22
rect 6 20 8 22
rect 2 15 8 20
rect 2 13 4 15
rect 6 13 8 15
rect 22 21 26 33
rect 25 15 29 17
rect 25 13 26 15
rect 28 13 29 15
rect 2 7 8 13
rect 25 7 29 13
rect -2 5 34 7
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 34 5
rect -2 -2 2 3
rect 30 -2 34 3
<< alu2 >>
rect -2 85 34 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 80 34 83
rect -2 5 34 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 34 5
rect -2 -2 34 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
<< polyct0 >>
rect 7 44 9 46
rect 17 44 19 46
<< polyct1 >>
rect 13 34 15 36
rect 23 34 25 36
<< ndifct0 >>
rect 15 22 17 24
rect 15 15 17 17
<< ndifct1 >>
rect 4 20 6 22
rect 4 13 6 15
rect 26 13 28 15
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
<< pdifct1 >>
rect 4 72 6 74
rect 4 65 6 67
rect 15 71 17 73
rect 15 63 17 65
rect 15 55 17 57
rect 26 72 28 74
rect 26 65 28 67
<< alu0 >>
rect 4 46 21 47
rect 4 44 7 46
rect 9 44 17 46
rect 19 44 21 46
rect 4 43 21 44
rect 4 30 8 43
rect 4 26 18 30
rect 14 24 18 26
rect 14 22 15 24
rect 17 22 18 24
rect 14 17 18 22
rect 14 15 15 17
rect 17 15 18 17
rect 14 13 18 15
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect -1 3 1 5
rect 31 3 33 5
<< labels >>
rlabel alu1 8 56 8 56 6 z
rlabel pdifct1 16 64 16 64 6 z
rlabel alu1 24 28 24 28 6 z
rlabel alu1 24 56 24 56 6 z
rlabel alu2 16 4 16 4 6 vss
rlabel alu2 16 84 16 84 6 vdd
<< end >>
