magic
tech scmos
timestamp 1199202772
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 9 39 11 50
rect 19 47 21 50
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 19 41 25 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 12 30 14 33
rect 19 30 21 41
rect 29 39 31 50
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 26 33 35 35
rect 26 30 28 33
rect 12 6 14 10
rect 19 6 21 10
rect 26 6 28 10
<< ndif >>
rect 7 22 12 30
rect 5 20 12 22
rect 5 18 7 20
rect 9 18 12 20
rect 5 16 12 18
rect 7 10 12 16
rect 14 10 19 30
rect 21 10 26 30
rect 28 13 36 30
rect 28 11 32 13
rect 34 11 36 13
rect 28 10 36 11
rect 30 8 36 10
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 50 19 59
rect 21 61 29 70
rect 21 59 24 61
rect 26 59 29 61
rect 21 54 29 59
rect 21 52 24 54
rect 26 52 29 54
rect 21 50 29 52
rect 31 68 38 70
rect 31 66 34 68
rect 36 66 38 68
rect 31 61 38 66
rect 31 59 34 61
rect 36 59 38 61
rect 31 50 38 59
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 61 7 63
rect 2 59 4 61
rect 6 59 7 61
rect 2 54 7 59
rect 23 61 27 63
rect 23 59 24 61
rect 26 59 27 61
rect 23 54 27 59
rect 2 52 4 54
rect 6 52 24 54
rect 26 52 27 54
rect 2 50 27 52
rect 2 21 6 50
rect 34 46 38 55
rect 19 45 38 46
rect 19 43 21 45
rect 23 43 38 45
rect 19 42 38 43
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 25 37 38 38
rect 25 35 31 37
rect 33 35 38 37
rect 25 34 38 35
rect 10 25 23 30
rect 2 20 11 21
rect 2 18 7 20
rect 9 18 11 20
rect 2 17 11 18
rect 34 17 38 34
rect -2 11 32 12
rect 34 11 42 12
rect -2 1 42 11
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 26 10 28 30
<< pmos >>
rect 9 50 11 70
rect 19 50 21 70
rect 29 50 31 70
<< polyct1 >>
rect 21 43 23 45
rect 11 35 13 37
rect 31 35 33 37
<< ndifct0 >>
rect 32 12 34 13
<< ndifct1 >>
rect 7 18 9 20
rect 32 11 34 12
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 66 16 68
rect 14 59 16 61
rect 34 66 36 68
rect 34 59 36 61
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
rect 24 59 26 61
rect 24 52 26 54
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 61 18 66
rect 32 66 34 68
rect 36 66 38 68
rect 12 59 14 61
rect 16 59 18 61
rect 12 58 18 59
rect 32 61 38 66
rect 32 59 34 61
rect 36 59 38 61
rect 32 58 38 59
rect 30 13 36 14
rect 30 12 32 13
rect 34 12 36 13
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 32 12 32 6 c
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 28 20 28 6 c
rlabel alu1 28 36 28 36 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 24 36 24 6 a
rlabel alu1 36 52 36 52 6 b
<< end >>
