magic
tech scmos
timestamp 1199541851
<< ab >>
rect 0 0 200 100
<< nwell >>
rect -2 48 202 104
<< pwell >>
rect -2 -4 202 48
<< poly >>
rect 81 95 83 98
rect 93 95 95 98
rect 11 83 13 86
rect 23 83 25 86
rect 35 83 37 86
rect 47 83 49 86
rect 57 83 59 86
rect 11 43 13 65
rect 23 43 25 65
rect 35 53 37 65
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 25 43
rect 17 39 19 41
rect 21 39 25 41
rect 17 37 25 39
rect 33 51 43 53
rect 33 49 39 51
rect 41 49 43 51
rect 33 47 43 49
rect 11 27 13 37
rect 21 29 23 37
rect 33 25 35 47
rect 47 43 49 57
rect 57 53 59 57
rect 121 83 123 86
rect 133 83 135 86
rect 143 83 145 86
rect 155 83 157 86
rect 81 53 83 55
rect 57 51 63 53
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 81 51 89 53
rect 81 49 85 51
rect 87 49 89 51
rect 81 47 89 49
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 45 37 53 39
rect 45 25 47 37
rect 57 25 59 47
rect 81 25 83 47
rect 93 41 95 55
rect 121 43 123 69
rect 133 67 135 69
rect 143 67 145 69
rect 131 65 135 67
rect 141 65 145 67
rect 167 79 169 82
rect 177 79 179 82
rect 187 79 189 82
rect 131 43 133 65
rect 141 43 143 65
rect 155 63 157 65
rect 153 61 157 63
rect 153 43 155 61
rect 167 53 169 65
rect 177 53 179 65
rect 167 51 173 53
rect 167 49 169 51
rect 171 49 173 51
rect 107 41 113 43
rect 93 39 109 41
rect 111 39 113 41
rect 93 25 95 39
rect 107 37 113 39
rect 117 41 123 43
rect 117 39 119 41
rect 121 39 123 41
rect 117 37 123 39
rect 127 41 133 43
rect 127 39 129 41
rect 131 39 133 41
rect 127 37 133 39
rect 137 41 143 43
rect 137 39 139 41
rect 141 39 143 41
rect 137 37 143 39
rect 147 41 155 43
rect 147 39 149 41
rect 151 39 155 41
rect 147 37 155 39
rect 121 25 123 37
rect 131 25 133 37
rect 141 25 143 37
rect 153 27 155 37
rect 165 47 173 49
rect 177 51 183 53
rect 177 49 179 51
rect 181 49 183 51
rect 177 47 183 49
rect 11 14 13 17
rect 21 14 23 17
rect 33 14 35 17
rect 45 14 47 17
rect 57 14 59 17
rect 165 25 167 47
rect 177 29 179 47
rect 175 27 179 29
rect 187 43 189 65
rect 187 41 193 43
rect 187 39 189 41
rect 191 39 193 41
rect 187 37 193 39
rect 175 25 177 27
rect 187 25 189 37
rect 121 14 123 17
rect 131 14 133 17
rect 141 14 143 17
rect 153 14 155 17
rect 165 14 167 17
rect 175 14 177 17
rect 187 14 189 17
rect 81 2 83 5
rect 93 2 95 5
<< ndif >>
rect 17 27 21 29
rect 3 17 11 27
rect 13 17 21 27
rect 23 25 31 29
rect 149 25 153 27
rect 23 21 33 25
rect 23 19 27 21
rect 29 19 33 21
rect 23 17 33 19
rect 35 21 45 25
rect 35 19 39 21
rect 41 19 45 21
rect 35 17 45 19
rect 47 17 57 25
rect 59 21 67 25
rect 59 19 63 21
rect 65 19 67 21
rect 59 17 67 19
rect 73 21 81 25
rect 73 19 75 21
rect 77 19 81 21
rect 3 11 9 17
rect 49 11 55 17
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
rect 73 5 81 19
rect 83 11 93 25
rect 83 9 87 11
rect 89 9 93 11
rect 83 5 93 9
rect 95 21 103 25
rect 95 19 99 21
rect 101 19 103 21
rect 95 5 103 19
rect 113 17 121 25
rect 123 17 131 25
rect 133 17 141 25
rect 143 21 153 25
rect 143 19 147 21
rect 149 19 153 21
rect 143 17 153 19
rect 155 25 159 27
rect 155 21 165 25
rect 155 19 159 21
rect 161 19 165 21
rect 155 17 165 19
rect 167 17 175 25
rect 177 21 187 25
rect 177 19 181 21
rect 183 19 187 21
rect 177 17 187 19
rect 189 21 197 25
rect 189 19 193 21
rect 195 19 197 21
rect 189 17 197 19
rect 113 11 119 17
rect 169 11 173 17
rect 113 9 115 11
rect 117 9 119 11
rect 113 7 119 9
rect 168 9 174 11
rect 168 7 170 9
rect 172 7 174 9
rect 168 5 174 7
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 83 21 89
rect 3 81 11 83
rect 3 79 5 81
rect 7 79 11 81
rect 3 65 11 79
rect 13 65 23 83
rect 25 81 35 83
rect 25 79 29 81
rect 31 79 35 81
rect 25 65 35 79
rect 37 71 47 83
rect 37 69 41 71
rect 43 69 47 71
rect 37 65 47 69
rect 40 57 47 65
rect 49 57 57 83
rect 59 81 67 83
rect 59 79 63 81
rect 65 79 67 81
rect 59 57 67 79
rect 73 61 81 95
rect 73 59 75 61
rect 77 59 81 61
rect 73 55 81 59
rect 83 91 93 95
rect 83 89 87 91
rect 89 89 93 91
rect 83 55 93 89
rect 95 71 103 95
rect 136 93 142 95
rect 95 69 99 71
rect 101 69 103 71
rect 110 91 118 93
rect 110 89 113 91
rect 115 89 118 91
rect 136 91 138 93
rect 140 91 142 93
rect 136 89 142 91
rect 110 83 118 89
rect 137 83 141 89
rect 110 69 121 83
rect 123 81 133 83
rect 123 79 127 81
rect 129 79 133 81
rect 123 69 133 79
rect 135 69 143 83
rect 145 81 155 83
rect 145 79 149 81
rect 151 79 155 81
rect 145 69 155 79
rect 95 61 103 69
rect 95 59 99 61
rect 101 59 103 61
rect 95 55 103 59
rect 147 65 155 69
rect 157 79 164 83
rect 191 81 197 83
rect 191 79 193 81
rect 195 79 197 81
rect 157 71 167 79
rect 157 69 161 71
rect 163 69 167 71
rect 157 65 167 69
rect 169 65 177 79
rect 179 65 187 79
rect 189 65 197 79
<< alu1 >>
rect -2 95 202 100
rect -2 93 31 95
rect 33 93 39 95
rect 41 93 47 95
rect 49 93 55 95
rect 57 93 63 95
rect 65 93 151 95
rect 153 93 159 95
rect 161 93 167 95
rect 169 93 175 95
rect 177 93 183 95
rect 185 93 202 95
rect -2 91 138 93
rect 140 91 202 93
rect -2 89 17 91
rect 19 89 87 91
rect 89 89 113 91
rect 115 89 202 91
rect -2 88 202 89
rect 4 81 8 82
rect 28 81 32 82
rect 62 81 66 82
rect 126 81 130 82
rect 148 81 152 82
rect 192 81 196 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 63 81
rect 65 79 66 81
rect 4 78 8 79
rect 28 78 32 79
rect 62 78 66 79
rect 87 79 113 81
rect 8 41 12 72
rect 8 39 9 41
rect 11 39 12 41
rect 8 18 12 39
rect 18 41 22 72
rect 40 71 44 72
rect 87 71 89 79
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 29 69 41 71
rect 43 69 89 71
rect 29 22 31 69
rect 40 68 44 69
rect 38 51 42 62
rect 38 49 39 51
rect 41 49 42 51
rect 38 28 42 49
rect 48 41 52 62
rect 48 39 49 41
rect 51 39 52 41
rect 48 28 52 39
rect 58 51 62 62
rect 58 49 59 51
rect 61 49 62 51
rect 58 28 62 49
rect 68 61 78 62
rect 68 59 75 61
rect 77 59 78 61
rect 68 58 78 59
rect 68 32 72 58
rect 87 52 89 69
rect 84 51 89 52
rect 84 49 85 51
rect 87 49 89 51
rect 98 71 102 72
rect 98 69 99 71
rect 101 69 102 71
rect 111 71 113 79
rect 126 79 127 81
rect 129 79 149 81
rect 151 79 193 81
rect 195 79 196 81
rect 126 78 130 79
rect 148 78 152 79
rect 192 78 196 79
rect 159 71 164 72
rect 111 69 151 71
rect 98 61 102 69
rect 98 59 99 61
rect 101 59 102 61
rect 84 48 88 49
rect 68 28 82 32
rect 78 22 82 28
rect 26 21 31 22
rect 26 19 27 21
rect 29 19 31 21
rect 38 21 42 22
rect 62 21 66 22
rect 38 19 39 21
rect 41 19 63 21
rect 65 19 66 21
rect 26 18 30 19
rect 38 18 42 19
rect 62 18 66 19
rect 74 21 82 22
rect 74 19 75 21
rect 77 19 82 21
rect 74 18 82 19
rect 98 21 102 59
rect 108 41 112 42
rect 108 39 109 41
rect 111 39 112 41
rect 108 38 112 39
rect 118 41 122 62
rect 118 39 119 41
rect 121 39 122 41
rect 98 19 99 21
rect 101 19 102 21
rect 109 21 111 38
rect 118 28 122 39
rect 128 41 132 62
rect 128 39 129 41
rect 131 39 132 41
rect 128 28 132 39
rect 138 41 142 62
rect 149 42 151 69
rect 159 69 161 71
rect 163 69 164 71
rect 159 68 164 69
rect 138 39 139 41
rect 141 39 142 41
rect 138 28 142 39
rect 148 41 152 42
rect 148 39 149 41
rect 151 39 152 41
rect 148 38 152 39
rect 159 31 161 68
rect 149 29 161 31
rect 168 51 172 62
rect 168 49 169 51
rect 171 49 172 51
rect 149 22 151 29
rect 168 28 172 49
rect 178 51 182 72
rect 178 49 179 51
rect 181 49 182 51
rect 178 28 182 49
rect 188 41 192 72
rect 188 39 189 41
rect 191 39 192 41
rect 188 28 192 39
rect 146 21 151 22
rect 109 19 147 21
rect 149 19 151 21
rect 98 18 102 19
rect 146 18 151 19
rect 158 21 162 22
rect 180 21 184 22
rect 158 19 159 21
rect 161 19 181 21
rect 183 19 184 21
rect 158 18 162 19
rect 180 18 184 19
rect 192 21 196 22
rect 192 19 193 21
rect 195 19 196 21
rect 192 12 196 19
rect -2 11 202 12
rect -2 9 5 11
rect 7 9 51 11
rect 53 9 87 11
rect 89 9 115 11
rect 117 9 202 11
rect -2 7 19 9
rect 21 7 29 9
rect 31 7 39 9
rect 41 7 127 9
rect 129 7 137 9
rect 139 7 147 9
rect 149 7 158 9
rect 160 7 170 9
rect 172 7 183 9
rect 185 7 191 9
rect 193 7 202 9
rect -2 0 202 7
<< ptie >>
rect 17 9 43 11
rect 17 7 19 9
rect 21 7 29 9
rect 31 7 39 9
rect 41 7 43 9
rect 17 5 43 7
rect 125 9 162 11
rect 125 7 127 9
rect 129 7 137 9
rect 139 7 147 9
rect 149 7 158 9
rect 160 7 162 9
rect 125 5 162 7
rect 181 9 195 11
rect 181 7 183 9
rect 185 7 191 9
rect 193 7 195 9
rect 181 5 195 7
<< ntie >>
rect 29 95 67 97
rect 149 95 187 97
rect 29 93 31 95
rect 33 93 39 95
rect 41 93 47 95
rect 49 93 55 95
rect 57 93 63 95
rect 65 93 67 95
rect 29 91 67 93
rect 149 93 151 95
rect 153 93 159 95
rect 161 93 167 95
rect 169 93 175 95
rect 177 93 183 95
rect 185 93 187 95
rect 149 91 187 93
<< nmos >>
rect 11 17 13 27
rect 21 17 23 29
rect 33 17 35 25
rect 45 17 47 25
rect 57 17 59 25
rect 81 5 83 25
rect 93 5 95 25
rect 121 17 123 25
rect 131 17 133 25
rect 141 17 143 25
rect 153 17 155 27
rect 165 17 167 25
rect 175 17 177 25
rect 187 17 189 25
<< pmos >>
rect 11 65 13 83
rect 23 65 25 83
rect 35 65 37 83
rect 47 57 49 83
rect 57 57 59 83
rect 81 55 83 95
rect 93 55 95 95
rect 121 69 123 83
rect 133 69 135 83
rect 143 69 145 83
rect 155 65 157 83
rect 167 65 169 79
rect 177 65 179 79
rect 187 65 189 79
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 39 49 41 51
rect 59 49 61 51
rect 85 49 87 51
rect 49 39 51 41
rect 169 49 171 51
rect 109 39 111 41
rect 119 39 121 41
rect 129 39 131 41
rect 139 39 141 41
rect 149 39 151 41
rect 179 49 181 51
rect 189 39 191 41
<< ndifct1 >>
rect 27 19 29 21
rect 39 19 41 21
rect 63 19 65 21
rect 75 19 77 21
rect 5 9 7 11
rect 51 9 53 11
rect 87 9 89 11
rect 99 19 101 21
rect 147 19 149 21
rect 159 19 161 21
rect 181 19 183 21
rect 193 19 195 21
rect 115 9 117 11
rect 170 7 172 9
<< ntiect1 >>
rect 31 93 33 95
rect 39 93 41 95
rect 47 93 49 95
rect 55 93 57 95
rect 63 93 65 95
rect 151 93 153 95
rect 159 93 161 95
rect 167 93 169 95
rect 175 93 177 95
rect 183 93 185 95
<< ptiect1 >>
rect 19 7 21 9
rect 29 7 31 9
rect 39 7 41 9
rect 127 7 129 9
rect 137 7 139 9
rect 147 7 149 9
rect 158 7 160 9
rect 183 7 185 9
rect 191 7 193 9
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 29 79 31 81
rect 41 69 43 71
rect 63 79 65 81
rect 75 59 77 61
rect 87 89 89 91
rect 99 69 101 71
rect 113 89 115 91
rect 138 91 140 93
rect 127 79 129 81
rect 149 79 151 81
rect 99 59 101 61
rect 193 79 195 81
rect 161 69 163 71
<< labels >>
rlabel alu1 10 45 10 45 6 a1
rlabel alu1 20 50 20 50 6 b1
rlabel alu1 60 45 60 45 6 b2
rlabel alu1 50 45 50 45 6 a2
rlabel alu1 70 45 70 45 6 cout
rlabel alu1 40 45 40 45 6 cin1
rlabel alu1 100 6 100 6 6 vss
rlabel alu1 80 25 80 25 6 cout
rlabel alu1 100 45 100 45 6 sout
rlabel alu1 100 94 100 94 6 vdd
rlabel alu1 140 45 140 45 6 cin2
rlabel alu1 130 45 130 45 6 b3
rlabel alu1 120 45 120 45 6 a3
rlabel alu1 170 45 170 45 6 cin3
rlabel polyct1 180 50 180 50 6 a4
rlabel alu1 190 50 190 50 6 b4
<< end >>
