magic
tech scmos
timestamp 1199201699
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 9 57 11 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 33 41 35
rect 49 33 51 39
rect 59 36 61 39
rect 58 34 64 36
rect 9 26 11 33
rect 19 26 21 33
rect 29 31 33 33
rect 35 31 37 33
rect 29 29 37 31
rect 48 31 54 33
rect 48 29 50 31
rect 52 29 54 31
rect 29 26 31 29
rect 41 27 54 29
rect 58 32 60 34
rect 62 32 64 34
rect 58 30 64 32
rect 9 11 11 15
rect 41 18 43 27
rect 58 23 60 30
rect 68 25 74 27
rect 68 23 70 25
rect 72 23 74 25
rect 48 21 60 23
rect 48 18 50 21
rect 58 18 60 21
rect 65 21 74 23
rect 65 18 67 21
rect 19 2 21 6
rect 29 2 31 6
rect 41 2 43 7
rect 48 2 50 7
rect 58 2 60 7
rect 65 2 67 7
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 4 15 9 20
rect 11 19 19 26
rect 11 17 14 19
rect 16 17 19 19
rect 11 15 19 17
rect 13 6 19 15
rect 21 24 29 26
rect 21 22 24 24
rect 26 22 29 24
rect 21 17 29 22
rect 21 15 24 17
rect 26 15 29 17
rect 21 6 29 15
rect 31 18 39 26
rect 31 16 34 18
rect 36 16 41 18
rect 31 10 41 16
rect 31 8 34 10
rect 36 8 41 10
rect 31 7 41 8
rect 43 7 48 18
rect 50 16 58 18
rect 50 14 53 16
rect 55 14 58 16
rect 50 7 58 14
rect 60 7 65 18
rect 67 11 75 18
rect 67 9 70 11
rect 72 9 75 11
rect 67 7 75 9
rect 31 6 39 7
<< pdif >>
rect 14 57 19 66
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 48 9 53
rect 2 46 4 48
rect 6 46 9 48
rect 2 38 9 46
rect 11 55 19 57
rect 11 53 14 55
rect 16 53 19 55
rect 11 48 19 53
rect 11 46 14 48
rect 16 46 19 48
rect 11 38 19 46
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 50 39 55
rect 31 48 34 50
rect 36 48 39 50
rect 31 38 39 48
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 39 49 55
rect 51 57 59 66
rect 51 55 54 57
rect 56 55 59 57
rect 51 50 59 55
rect 51 48 54 50
rect 56 48 59 50
rect 51 39 59 48
rect 61 59 67 66
rect 61 57 69 59
rect 61 55 64 57
rect 66 55 69 57
rect 61 50 69 55
rect 61 48 64 50
rect 66 48 69 50
rect 61 39 69 48
rect 41 38 47 39
<< alu1 >>
rect -2 67 82 72
rect -2 65 5 67
rect 7 65 73 67
rect 75 65 82 67
rect -2 64 82 65
rect 12 55 18 56
rect 12 53 14 55
rect 16 53 18 55
rect 33 57 38 59
rect 33 55 34 57
rect 36 55 38 57
rect 12 50 18 53
rect 33 50 38 55
rect 12 48 34 50
rect 36 48 38 50
rect 12 46 14 48
rect 16 46 38 48
rect 12 45 22 46
rect 18 35 22 45
rect 2 34 22 35
rect 2 30 27 34
rect 2 24 7 30
rect 2 22 4 24
rect 6 22 7 24
rect 2 20 7 22
rect 23 24 27 30
rect 23 22 24 24
rect 26 22 27 24
rect 23 17 27 22
rect 23 15 24 17
rect 26 15 27 17
rect 23 13 27 15
rect 49 31 54 35
rect 49 29 50 31
rect 52 29 54 31
rect 58 34 63 43
rect 58 32 60 34
rect 62 32 71 34
rect 58 30 71 32
rect 49 26 54 29
rect 49 25 74 26
rect 49 23 70 25
rect 72 23 74 25
rect 49 22 74 23
rect -2 7 82 8
rect -2 5 5 7
rect 7 5 82 7
rect -2 0 82 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 71 67 77 69
rect 3 63 9 65
rect 71 65 73 67
rect 75 65 77 67
rect 71 63 77 65
<< nmos >>
rect 9 15 11 26
rect 19 6 21 26
rect 29 6 31 26
rect 41 7 43 18
rect 48 7 50 18
rect 58 7 60 18
rect 65 7 67 18
<< pmos >>
rect 9 38 11 57
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 39 51 66
rect 59 39 61 66
<< polyct0 >>
rect 33 31 35 33
<< polyct1 >>
rect 50 29 52 31
rect 60 32 62 34
rect 70 23 72 25
<< ndifct0 >>
rect 14 17 16 19
rect 34 16 36 18
rect 34 8 36 10
rect 53 14 55 16
rect 70 9 72 11
<< ndifct1 >>
rect 4 22 6 24
rect 24 22 26 24
rect 24 15 26 17
<< ntiect1 >>
rect 5 65 7 67
rect 73 65 75 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 4 53 6 55
rect 4 46 6 48
rect 24 62 26 64
rect 24 55 26 57
rect 44 62 46 64
rect 44 55 46 57
rect 54 55 56 57
rect 54 48 56 50
rect 64 55 66 57
rect 64 48 66 50
<< pdifct1 >>
rect 14 53 16 55
rect 14 46 16 48
rect 34 55 36 57
rect 34 48 36 50
<< alu0 >>
rect 3 55 7 64
rect 22 62 24 64
rect 26 62 28 64
rect 22 57 28 62
rect 42 62 44 64
rect 46 62 48 64
rect 3 53 4 55
rect 6 53 7 55
rect 3 48 7 53
rect 3 46 4 48
rect 6 46 7 48
rect 3 44 7 46
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 42 57 48 62
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 53 57 57 59
rect 53 55 54 57
rect 56 55 57 57
rect 53 50 57 55
rect 41 48 54 50
rect 56 48 57 50
rect 41 46 57 48
rect 63 57 67 64
rect 63 55 64 57
rect 66 55 67 57
rect 63 50 67 55
rect 63 48 64 50
rect 66 48 67 50
rect 63 46 67 48
rect 41 34 45 46
rect 31 33 45 34
rect 31 31 33 33
rect 35 31 45 33
rect 31 30 45 31
rect 13 19 17 21
rect 13 17 14 19
rect 16 17 17 19
rect 13 8 17 17
rect 33 18 37 20
rect 33 16 34 18
rect 36 16 37 18
rect 33 10 37 16
rect 41 17 45 30
rect 41 16 57 17
rect 41 14 53 16
rect 55 14 57 16
rect 41 13 57 14
rect 33 8 34 10
rect 36 8 37 10
rect 69 11 73 13
rect 69 9 70 11
rect 72 9 73 11
rect 69 8 73 9
<< labels >>
rlabel alu0 49 15 49 15 6 zn
rlabel alu0 38 32 38 32 6 zn
rlabel alu0 55 52 55 52 6 zn
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 32 12 32 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 52 28 52 28 6 a
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 60 24 60 24 6 a
rlabel alu1 68 32 68 32 6 b
rlabel alu1 68 24 68 24 6 a
rlabel alu1 60 40 60 40 6 b
<< end >>
