magic
tech scmos
timestamp 1199203585
<< ab >>
rect 0 0 112 72
<< nwell >>
rect -5 32 117 77
<< pwell >>
rect -5 -5 117 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 61 66 63 70
rect 71 66 73 70
rect 29 59 31 64
rect 39 59 41 64
rect 48 42 54 44
rect 48 40 50 42
rect 52 40 54 42
rect 48 38 54 40
rect 81 59 83 64
rect 91 59 93 64
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 48 35 50 38
rect 9 33 25 35
rect 29 33 50 35
rect 61 35 63 38
rect 71 35 73 38
rect 81 35 83 38
rect 91 35 93 38
rect 61 33 73 35
rect 78 33 103 35
rect 16 31 21 33
rect 23 31 25 33
rect 16 29 25 31
rect 9 24 11 29
rect 16 27 28 29
rect 16 24 18 27
rect 26 24 28 27
rect 33 24 35 33
rect 65 31 67 33
rect 69 31 71 33
rect 65 29 71 31
rect 78 29 80 33
rect 97 31 99 33
rect 101 31 103 33
rect 97 29 103 31
rect 65 24 67 29
rect 75 27 80 29
rect 75 24 77 27
rect 85 25 91 27
rect 9 4 11 12
rect 16 8 18 12
rect 26 8 28 12
rect 33 4 35 12
rect 9 2 35 4
rect 85 23 87 25
rect 89 23 91 25
rect 85 21 97 23
rect 85 18 87 21
rect 95 18 97 21
rect 65 2 67 6
rect 75 2 77 6
rect 85 4 87 9
rect 95 4 97 9
<< ndif >>
rect 2 16 9 24
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 12 16 24
rect 18 22 26 24
rect 18 20 21 22
rect 23 20 26 22
rect 18 12 26 20
rect 28 12 33 24
rect 35 12 44 24
rect 37 7 44 12
rect 37 5 39 7
rect 41 5 44 7
rect 37 3 44 5
rect 60 19 65 24
rect 58 17 65 19
rect 58 15 60 17
rect 62 15 65 17
rect 58 13 65 15
rect 60 6 65 13
rect 67 22 75 24
rect 67 20 70 22
rect 72 20 75 22
rect 67 6 75 20
rect 77 18 83 24
rect 77 13 85 18
rect 77 11 80 13
rect 82 11 85 13
rect 77 9 85 11
rect 87 16 95 18
rect 87 14 90 16
rect 92 14 95 16
rect 87 9 95 14
rect 97 9 105 18
rect 77 6 83 9
rect 99 7 105 9
rect 99 5 101 7
rect 103 5 105 7
rect 99 3 105 5
<< pdif >>
rect 4 59 9 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 4 38 9 46
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 59 26 66
rect 54 64 61 66
rect 54 62 56 64
rect 58 62 61 64
rect 21 57 29 59
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 42 39 59
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 57 48 59
rect 41 55 44 57
rect 46 55 48 57
rect 41 53 48 55
rect 54 57 61 62
rect 54 55 56 57
rect 58 55 61 57
rect 54 53 61 55
rect 41 38 46 53
rect 56 38 61 53
rect 63 56 71 66
rect 63 54 66 56
rect 68 54 71 56
rect 63 49 71 54
rect 63 47 66 49
rect 68 47 71 49
rect 63 38 71 47
rect 73 59 79 66
rect 73 57 81 59
rect 73 55 76 57
rect 78 55 81 57
rect 73 38 81 55
rect 83 42 91 59
rect 83 40 86 42
rect 88 40 91 42
rect 83 38 91 40
rect 93 57 100 59
rect 93 55 96 57
rect 98 55 100 57
rect 93 38 100 55
<< alu1 >>
rect -2 67 114 72
rect -2 65 105 67
rect 107 65 114 67
rect -2 64 114 65
rect 2 57 48 58
rect 2 55 4 57
rect 6 55 24 57
rect 26 55 44 57
rect 46 55 48 57
rect 2 54 48 55
rect 2 50 7 54
rect 2 48 4 50
rect 6 48 7 50
rect 2 46 7 48
rect 2 26 6 46
rect 97 34 103 42
rect 65 33 82 34
rect 65 31 67 33
rect 69 31 82 33
rect 65 30 82 31
rect 89 33 103 34
rect 89 31 99 33
rect 101 31 103 33
rect 89 30 103 31
rect 78 26 82 30
rect 2 22 24 26
rect 78 25 91 26
rect 78 23 87 25
rect 89 23 91 25
rect 78 22 91 23
rect 20 20 21 22
rect 23 20 24 22
rect 20 18 24 20
rect 20 17 64 18
rect 20 15 60 17
rect 62 15 64 17
rect 20 14 64 15
rect -2 7 114 8
rect -2 5 39 7
rect 41 5 50 7
rect 52 5 101 7
rect 103 5 114 7
rect -2 0 114 5
<< ptie >>
rect 48 7 54 24
rect 48 5 50 7
rect 52 5 54 7
rect 48 3 54 5
<< ntie >>
rect 103 67 109 69
rect 103 65 105 67
rect 107 65 109 67
rect 103 63 109 65
<< nmos >>
rect 9 12 11 24
rect 16 12 18 24
rect 26 12 28 24
rect 33 12 35 24
rect 65 6 67 24
rect 75 6 77 24
rect 85 9 87 18
rect 95 9 97 18
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 59
rect 39 38 41 59
rect 61 38 63 66
rect 71 38 73 66
rect 81 38 83 59
rect 91 38 93 59
<< polyct0 >>
rect 50 40 52 42
rect 21 31 23 33
<< polyct1 >>
rect 67 31 69 33
rect 99 31 101 33
rect 87 23 89 25
<< ndifct0 >>
rect 4 14 6 16
rect 70 20 72 22
rect 80 11 82 13
rect 90 14 92 16
<< ndifct1 >>
rect 21 20 23 22
rect 39 5 41 7
rect 60 15 62 17
rect 101 5 103 7
<< ntiect1 >>
rect 105 65 107 67
<< ptiect1 >>
rect 50 5 52 7
<< pdifct0 >>
rect 14 47 16 49
rect 14 40 16 42
rect 56 62 58 64
rect 34 40 36 42
rect 56 55 58 57
rect 66 54 68 56
rect 66 47 68 49
rect 76 55 78 57
rect 86 40 88 42
rect 96 55 98 57
<< pdifct1 >>
rect 4 55 6 57
rect 4 48 6 50
rect 24 55 26 57
rect 44 55 46 57
<< alu0 >>
rect 54 62 56 64
rect 58 62 60 64
rect 54 57 60 62
rect 54 55 56 57
rect 58 55 60 57
rect 54 54 60 55
rect 65 56 69 58
rect 65 54 66 56
rect 68 54 69 56
rect 74 57 80 64
rect 74 55 76 57
rect 78 55 80 57
rect 74 54 80 55
rect 94 57 100 64
rect 94 55 96 57
rect 98 55 100 57
rect 94 54 100 55
rect 65 50 69 54
rect 12 49 110 50
rect 12 47 14 49
rect 16 47 66 49
rect 68 47 110 49
rect 12 46 110 47
rect 12 42 17 46
rect 12 40 14 42
rect 16 40 17 42
rect 12 38 17 40
rect 32 42 38 43
rect 32 40 34 42
rect 36 40 38 42
rect 32 34 38 40
rect 49 42 53 46
rect 84 42 90 43
rect 49 40 50 42
rect 52 40 53 42
rect 49 38 53 40
rect 57 40 86 42
rect 88 40 90 42
rect 57 38 90 40
rect 57 34 61 38
rect 19 33 61 34
rect 19 31 21 33
rect 23 31 61 33
rect 19 30 61 31
rect 57 26 61 30
rect 57 22 73 26
rect 69 20 70 22
rect 72 20 73 22
rect 69 18 73 20
rect 3 16 7 18
rect 3 14 4 16
rect 6 14 7 16
rect 106 17 110 46
rect 88 16 110 17
rect 3 8 7 14
rect 79 13 83 15
rect 88 14 90 16
rect 92 14 110 16
rect 88 13 110 14
rect 79 11 80 13
rect 82 11 83 13
rect 79 8 83 11
<< labels >>
rlabel alu0 14 44 14 44 6 bn
rlabel alu0 51 44 51 44 6 bn
rlabel alu0 35 36 35 36 6 an
rlabel alu0 71 22 71 22 6 an
rlabel alu0 40 32 40 32 6 an
rlabel alu0 67 52 67 52 6 bn
rlabel alu0 99 15 99 15 6 bn
rlabel alu0 87 40 87 40 6 an
rlabel alu0 61 48 61 48 6 bn
rlabel alu1 20 24 20 24 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 56 12 56 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 56 4 56 4 6 vss
rlabel alu1 60 16 60 16 6 z
rlabel polyct1 68 32 68 32 6 b
rlabel alu1 76 32 76 32 6 b
rlabel alu1 56 68 56 68 6 vdd
rlabel alu1 84 24 84 24 6 b
rlabel alu1 92 32 92 32 6 a
rlabel alu1 100 36 100 36 6 a
<< end >>
