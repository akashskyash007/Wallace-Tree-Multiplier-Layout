magic
tech scmos
timestamp 1199469842
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 11 53 13 56
rect 23 53 25 56
rect 11 51 25 53
rect 17 49 19 51
rect 21 49 25 51
rect 17 47 25 49
rect 35 53 37 56
rect 47 53 49 56
rect 35 51 49 53
rect 35 49 37 51
rect 39 49 41 51
rect 35 47 41 49
rect 17 38 19 47
rect 35 43 39 47
rect 47 45 53 47
rect 47 44 49 45
rect 25 41 39 43
rect 25 38 27 41
rect 37 38 39 41
rect 45 43 49 44
rect 51 43 53 45
rect 45 41 53 43
rect 45 38 47 41
rect 17 2 19 6
rect 25 2 27 6
rect 37 2 39 6
rect 45 2 47 6
<< ndif >>
rect 8 21 17 38
rect 8 19 11 21
rect 13 19 17 21
rect 8 11 17 19
rect 8 9 11 11
rect 13 9 17 11
rect 8 6 17 9
rect 19 6 25 38
rect 27 31 37 38
rect 27 29 31 31
rect 33 29 37 31
rect 27 21 37 29
rect 27 19 31 21
rect 33 19 37 21
rect 27 6 37 19
rect 39 6 45 38
rect 47 21 55 38
rect 47 19 51 21
rect 53 19 55 21
rect 47 11 55 19
rect 47 9 51 11
rect 53 9 55 11
rect 47 6 55 9
<< pdif >>
rect 3 91 11 94
rect 3 89 5 91
rect 7 89 11 91
rect 3 81 11 89
rect 3 79 5 81
rect 7 79 11 81
rect 3 56 11 79
rect 13 71 23 94
rect 13 69 17 71
rect 19 69 23 71
rect 13 61 23 69
rect 13 59 17 61
rect 19 59 23 61
rect 13 56 23 59
rect 25 91 35 94
rect 25 89 29 91
rect 31 89 35 91
rect 25 81 35 89
rect 25 79 29 81
rect 31 79 35 81
rect 25 56 35 79
rect 37 81 47 94
rect 37 79 41 81
rect 43 79 47 81
rect 37 72 47 79
rect 37 70 41 72
rect 43 70 47 72
rect 37 56 47 70
rect 49 91 57 94
rect 49 89 53 91
rect 55 89 57 91
rect 49 81 57 89
rect 49 79 53 81
rect 55 79 57 81
rect 49 56 57 79
<< alu1 >>
rect -2 91 62 100
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 53 91
rect 55 89 62 91
rect -2 88 62 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 77 8 79
rect 28 81 32 88
rect 28 79 29 81
rect 31 79 32 81
rect 28 77 32 79
rect 38 81 44 83
rect 38 79 41 81
rect 43 79 44 81
rect 38 73 44 79
rect 52 81 56 88
rect 52 79 53 81
rect 55 79 56 81
rect 52 77 56 79
rect 16 72 44 73
rect 16 71 41 72
rect 16 69 17 71
rect 19 70 41 71
rect 43 70 44 72
rect 19 69 44 70
rect 16 68 44 69
rect 16 63 22 68
rect 8 61 22 63
rect 8 59 17 61
rect 19 59 22 61
rect 8 57 22 59
rect 36 58 53 62
rect 8 33 12 57
rect 18 51 22 53
rect 18 49 19 51
rect 21 49 22 51
rect 18 42 22 49
rect 36 51 42 58
rect 36 49 37 51
rect 39 49 42 51
rect 36 47 42 49
rect 48 45 52 53
rect 48 43 49 45
rect 51 43 52 45
rect 48 42 52 43
rect 18 37 52 42
rect 8 31 34 33
rect 8 29 31 31
rect 33 29 34 31
rect 8 27 34 29
rect 10 21 14 23
rect 10 19 11 21
rect 13 19 14 21
rect 10 12 14 19
rect 28 21 34 27
rect 28 19 31 21
rect 33 19 34 21
rect 28 17 34 19
rect 50 21 54 23
rect 50 19 51 21
rect 53 19 54 21
rect 50 12 54 19
rect -2 11 62 12
rect -2 9 11 11
rect 13 9 51 11
rect 53 9 62 11
rect -2 0 62 9
<< nmos >>
rect 17 6 19 38
rect 25 6 27 38
rect 37 6 39 38
rect 45 6 47 38
<< pmos >>
rect 11 56 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 47 56 49 94
<< polyct1 >>
rect 19 49 21 51
rect 37 49 39 51
rect 49 43 51 45
<< ndifct1 >>
rect 11 19 13 21
rect 11 9 13 11
rect 31 29 33 31
rect 31 19 33 21
rect 51 19 53 21
rect 51 9 53 11
<< pdifct1 >>
rect 5 89 7 91
rect 5 79 7 81
rect 17 69 19 71
rect 17 59 19 61
rect 29 89 31 91
rect 29 79 31 81
rect 41 79 43 81
rect 41 70 43 72
rect 53 89 55 91
rect 53 79 55 81
<< labels >>
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 45 20 45 6 a
rlabel alu1 20 30 20 30 6 z
rlabel alu1 20 65 20 65 6 z
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 30 25 30 25 6 z
rlabel alu1 30 40 30 40 6 a
rlabel alu1 40 40 40 40 6 a
rlabel alu1 30 70 30 70 6 z
rlabel alu1 40 55 40 55 6 b
rlabel alu1 40 75 40 75 6 z
rlabel alu1 30 94 30 94 6 vdd
rlabel alu1 50 45 50 45 6 a
rlabel alu1 50 60 50 60 6 b
<< end >>
