magic
tech scmos
timestamp 1199201963
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 57 11 62
rect 21 62 27 64
rect 21 60 23 62
rect 25 60 27 62
rect 21 58 27 60
rect 21 55 23 58
rect 9 39 11 45
rect 9 37 16 39
rect 9 35 12 37
rect 14 35 16 37
rect 9 33 16 35
rect 9 30 11 33
rect 21 30 23 45
rect 9 19 11 24
rect 21 18 23 23
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 11 27 21 30
rect 11 25 15 27
rect 17 25 21 27
rect 11 24 21 25
rect 13 23 21 24
rect 23 28 30 30
rect 23 26 26 28
rect 28 26 30 28
rect 23 23 30 26
<< pdif >>
rect 13 71 19 73
rect 13 69 15 71
rect 17 69 19 71
rect 13 57 19 69
rect 4 51 9 57
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 11 55 19 57
rect 11 45 21 55
rect 23 51 28 55
rect 23 49 30 51
rect 23 47 26 49
rect 28 47 30 49
rect 23 45 30 47
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 71 34 79
rect -2 69 15 71
rect 17 69 34 71
rect -2 68 34 69
rect 18 62 30 63
rect 18 60 23 62
rect 25 60 30 62
rect 18 57 30 60
rect 2 49 14 55
rect 18 49 22 57
rect 2 47 4 49
rect 6 47 7 49
rect 2 45 7 47
rect 2 29 6 45
rect 2 28 8 29
rect 2 26 4 28
rect 6 26 8 28
rect 2 25 8 26
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 24 11 30
rect 21 23 23 30
<< pmos >>
rect 9 45 11 57
rect 21 45 23 55
<< polyct0 >>
rect 12 35 14 37
<< polyct1 >>
rect 23 60 25 62
<< ndifct0 >>
rect 15 25 17 27
rect 26 26 28 28
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 26 47 28 49
<< pdifct1 >>
rect 15 69 17 71
rect 4 47 6 49
<< alu0 >>
rect 25 49 29 51
rect 25 47 26 49
rect 28 47 29 49
rect 25 38 29 47
rect 10 37 30 38
rect 10 35 12 37
rect 14 35 30 37
rect 10 34 30 35
rect 14 27 18 29
rect 14 25 15 27
rect 17 25 18 27
rect 24 28 30 34
rect 24 26 26 28
rect 28 26 30 28
rect 24 25 30 26
rect 14 12 18 25
<< labels >>
rlabel alu0 27 38 27 38 6 an
rlabel alu0 20 36 20 36 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 20 56 20 56 6 a
rlabel alu1 28 60 28 60 6 a
<< end >>
