magic
tech scmos
timestamp 1199202212
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 20 71 26 73
rect 20 69 22 71
rect 24 69 26 71
rect 20 67 26 69
rect 9 57 11 65
rect 9 47 11 50
rect 9 45 18 47
rect 12 43 14 45
rect 16 43 18 45
rect 12 33 18 43
rect 22 45 26 67
rect 36 66 38 71
rect 43 66 45 71
rect 36 55 38 58
rect 43 55 45 58
rect 32 53 38 55
rect 32 51 34 53
rect 36 51 38 53
rect 32 49 38 51
rect 42 53 48 55
rect 42 51 44 53
rect 46 51 48 53
rect 42 49 48 51
rect 22 41 37 45
rect 9 31 18 33
rect 23 35 29 37
rect 23 33 25 35
rect 27 33 29 35
rect 23 31 29 33
rect 33 35 37 41
rect 33 31 49 35
rect 9 28 11 31
rect 16 28 18 31
rect 26 28 28 31
rect 33 28 35 31
rect 40 28 42 31
rect 47 28 49 31
rect 9 6 11 22
rect 16 6 18 22
rect 26 17 28 22
rect 33 17 35 22
rect 40 17 42 22
rect 47 17 49 22
<< ndif >>
rect 2 26 9 28
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 11 22 16 28
rect 18 26 26 28
rect 18 24 21 26
rect 23 24 26 26
rect 18 22 26 24
rect 28 22 33 28
rect 35 22 40 28
rect 42 22 47 28
rect 49 26 56 28
rect 49 24 52 26
rect 54 24 56 26
rect 49 22 56 24
<< pdif >>
rect 2 54 9 57
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 11 54 18 57
rect 11 52 14 54
rect 16 52 18 54
rect 11 50 18 52
rect 28 71 34 73
rect 28 69 30 71
rect 32 69 34 71
rect 28 66 34 69
rect 28 58 36 66
rect 38 58 43 66
rect 45 62 56 66
rect 45 60 52 62
rect 54 60 56 62
rect 45 58 56 60
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 22 71
rect 24 69 30 71
rect 32 69 66 71
rect -2 68 66 69
rect 2 54 8 63
rect 2 52 4 54
rect 6 52 8 54
rect 2 38 8 52
rect 12 54 18 68
rect 12 52 14 54
rect 16 52 18 54
rect 12 50 18 52
rect 22 62 56 63
rect 22 60 52 62
rect 54 60 56 62
rect 22 59 56 60
rect 22 46 28 59
rect 12 45 28 46
rect 12 43 14 45
rect 16 43 28 45
rect 12 42 28 43
rect 33 53 39 55
rect 33 51 34 53
rect 36 51 39 53
rect 33 38 39 51
rect 2 32 19 38
rect 23 35 39 38
rect 23 33 25 35
rect 27 33 39 35
rect 23 32 39 33
rect 2 26 8 32
rect 2 24 4 26
rect 6 24 8 26
rect 2 17 8 24
rect 19 26 25 28
rect 19 24 21 26
rect 23 24 25 26
rect 19 12 25 24
rect 50 26 56 59
rect 50 24 52 26
rect 54 24 56 26
rect 50 17 56 24
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 22 11 28
rect 16 22 18 28
rect 26 22 28 28
rect 33 22 35 28
rect 40 22 42 28
rect 47 22 49 28
<< pmos >>
rect 9 50 11 57
rect 36 58 38 66
rect 43 58 45 66
<< polyct0 >>
rect 44 51 46 53
<< polyct1 >>
rect 22 69 24 71
rect 14 43 16 45
rect 34 51 36 53
rect 25 33 27 35
<< ndifct1 >>
rect 4 24 6 26
rect 21 24 23 26
rect 52 24 54 26
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct1 >>
rect 4 52 6 54
rect 14 52 16 54
rect 30 69 32 71
rect 52 60 54 62
<< alu0 >>
rect 43 53 47 55
rect 43 51 44 53
rect 46 51 47 53
rect 43 12 47 51
<< labels >>
rlabel polyct1 15 44 15 44 6 an
rlabel ndifct1 53 25 53 25 6 an
rlabel pdifct1 53 61 53 61 6 an
rlabel alu1 12 36 12 36 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 36 28 36 6 a
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 44 36 44 6 a
rlabel alu1 32 74 32 74 6 vdd
<< end >>
