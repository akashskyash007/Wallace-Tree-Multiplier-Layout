magic
tech scmos
timestamp 1199202588
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 10 61 16 63
rect 10 59 12 61
rect 14 59 16 61
rect 10 57 16 59
rect 10 50 12 57
rect 20 50 22 55
rect 10 39 12 42
rect 20 39 22 42
rect 9 36 12 39
rect 16 37 23 39
rect 9 30 11 36
rect 16 35 19 37
rect 21 35 23 37
rect 16 33 23 35
rect 16 30 18 33
rect 9 18 11 23
rect 16 18 18 23
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 23 9 26
rect 11 23 16 30
rect 18 23 27 30
rect 20 20 27 23
rect 20 18 22 20
rect 24 18 27 20
rect 20 16 27 18
<< pdif >>
rect 2 71 8 73
rect 2 69 4 71
rect 6 69 8 71
rect 2 50 8 69
rect 2 42 10 50
rect 12 46 20 50
rect 12 44 15 46
rect 17 44 20 46
rect 12 42 20 44
rect 22 48 30 50
rect 22 46 26 48
rect 28 46 30 48
rect 22 42 30 46
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 71 34 79
rect -2 69 4 71
rect 6 69 34 71
rect -2 68 34 69
rect 2 61 16 63
rect 2 59 12 61
rect 14 59 16 61
rect 2 58 16 59
rect 2 49 6 58
rect 10 46 19 47
rect 10 44 15 46
rect 17 44 19 46
rect 2 43 19 44
rect 2 40 14 43
rect 2 30 6 40
rect 18 37 30 39
rect 18 35 19 37
rect 21 35 30 37
rect 18 33 30 35
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 24 7 26
rect 26 25 30 33
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 23 11 30
rect 16 23 18 30
<< pmos >>
rect 10 42 12 50
rect 20 42 22 50
<< polyct1 >>
rect 12 59 14 61
rect 19 35 21 37
<< ndifct0 >>
rect 22 18 24 20
<< ndifct1 >>
rect 4 26 6 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 26 46 28 48
<< pdifct1 >>
rect 4 69 6 71
rect 15 44 17 46
<< alu0 >>
rect 25 48 29 68
rect 25 46 26 48
rect 28 46 29 48
rect 25 44 29 46
rect 20 20 26 21
rect 20 18 22 20
rect 24 18 26 20
rect 20 12 26 18
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 4 56 4 56 6 b
rlabel alu1 12 44 12 44 6 z
rlabel alu1 12 60 12 60 6 b
rlabel alu1 16 6 16 6 6 vss
rlabel polyct1 20 36 20 36 6 a
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 32 28 32 6 a
<< end >>
