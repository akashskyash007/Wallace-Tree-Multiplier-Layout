magic
tech scmos
timestamp 1199203467
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 11 71 34 73
rect 11 65 13 71
rect 9 62 13 65
rect 22 63 24 67
rect 32 63 34 71
rect 42 69 44 74
rect 49 69 51 74
rect 9 59 11 62
rect 22 48 24 51
rect 9 44 11 47
rect 22 46 27 48
rect 32 46 34 51
rect 42 46 44 51
rect 49 48 51 51
rect 9 42 15 44
rect 9 40 11 42
rect 13 40 15 42
rect 9 38 15 40
rect 13 35 15 38
rect 25 39 27 46
rect 39 44 44 46
rect 48 46 54 48
rect 48 44 50 46
rect 52 44 54 46
rect 25 37 31 39
rect 25 35 27 37
rect 29 35 31 37
rect 13 33 19 35
rect 25 33 31 35
rect 17 30 19 33
rect 29 30 31 33
rect 39 30 41 44
rect 48 42 54 44
rect 49 30 51 42
rect 7 20 13 22
rect 7 18 9 20
rect 11 18 13 20
rect 17 19 19 24
rect 7 16 13 18
rect 29 19 31 24
rect 11 14 13 16
rect 39 14 41 24
rect 49 19 51 24
rect 55 20 61 22
rect 55 18 57 20
rect 59 18 61 20
rect 55 16 61 18
rect 55 14 57 16
rect 11 12 57 14
<< ndif >>
rect 9 28 17 30
rect 9 26 11 28
rect 13 26 17 28
rect 9 24 17 26
rect 19 24 29 30
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 24 39 26
rect 41 28 49 30
rect 41 26 44 28
rect 46 26 49 28
rect 41 24 49 26
rect 51 28 58 30
rect 51 26 54 28
rect 56 26 58 28
rect 51 24 58 26
rect 21 20 27 24
rect 21 18 23 20
rect 25 18 27 20
rect 21 16 27 18
<< pdif >>
rect 53 71 60 73
rect 53 69 55 71
rect 57 69 60 71
rect 37 63 42 69
rect 15 61 22 63
rect 15 59 17 61
rect 19 59 22 61
rect 4 53 9 59
rect 2 51 9 53
rect 2 49 4 51
rect 6 49 9 51
rect 2 47 9 49
rect 11 51 22 59
rect 24 55 32 63
rect 24 53 27 55
rect 29 53 32 55
rect 24 51 32 53
rect 34 61 42 63
rect 34 59 37 61
rect 39 59 42 61
rect 34 51 42 59
rect 44 51 49 69
rect 51 51 60 69
rect 11 47 20 51
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 55 71
rect 57 69 66 71
rect -2 68 66 69
rect 35 61 62 62
rect 35 59 37 61
rect 39 59 62 61
rect 35 58 62 59
rect 17 47 23 54
rect 10 42 23 47
rect 10 40 11 42
rect 13 40 14 42
rect 10 38 14 40
rect 18 37 31 38
rect 18 35 27 37
rect 29 35 31 37
rect 18 34 31 35
rect 18 25 22 34
rect 58 38 62 58
rect 42 34 62 38
rect 42 28 47 34
rect 42 26 44 28
rect 46 26 47 28
rect 42 24 47 26
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 17 24 19 30
rect 29 24 31 30
rect 39 24 41 30
rect 49 24 51 30
<< pmos >>
rect 9 47 11 59
rect 22 51 24 63
rect 32 51 34 63
rect 42 51 44 69
rect 49 51 51 69
<< polyct0 >>
rect 50 44 52 46
rect 9 18 11 20
rect 57 18 59 20
<< polyct1 >>
rect 11 40 13 42
rect 27 35 29 37
<< ndifct0 >>
rect 11 26 13 28
rect 34 26 36 28
rect 54 26 56 28
rect 23 18 25 20
<< ndifct1 >>
rect 44 26 46 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 17 59 19 61
rect 4 49 6 51
rect 27 53 29 55
<< pdifct1 >>
rect 55 69 57 71
rect 37 59 39 61
<< alu0 >>
rect 15 61 21 68
rect 15 59 17 61
rect 19 59 21 61
rect 15 58 21 59
rect 26 55 30 57
rect 2 51 7 53
rect 2 49 4 51
rect 6 49 7 51
rect 2 47 7 49
rect 26 53 27 55
rect 29 54 30 55
rect 29 53 38 54
rect 26 50 38 53
rect 2 30 6 47
rect 34 47 38 50
rect 34 46 54 47
rect 34 44 50 46
rect 52 44 54 46
rect 34 43 54 44
rect 2 28 14 30
rect 2 26 11 28
rect 13 26 14 28
rect 7 24 14 26
rect 34 30 38 43
rect 33 28 38 30
rect 33 26 34 28
rect 36 26 38 28
rect 33 24 38 26
rect 53 28 57 30
rect 53 26 54 28
rect 56 26 57 28
rect 7 20 13 24
rect 53 21 57 26
rect 7 18 9 20
rect 11 18 13 20
rect 7 17 13 18
rect 21 20 27 21
rect 21 18 23 20
rect 25 18 27 20
rect 21 12 27 18
rect 53 20 61 21
rect 53 18 57 20
rect 59 18 61 20
rect 53 17 61 18
<< labels >>
rlabel alu0 10 23 10 23 6 bn
rlabel alu0 10 27 10 27 6 bn
rlabel alu0 4 50 4 50 6 bn
rlabel alu0 36 39 36 39 6 an
rlabel alu0 32 52 32 52 6 an
rlabel alu0 57 19 57 19 6 bn
rlabel alu0 55 23 55 23 6 bn
rlabel alu0 44 45 44 45 6 an
rlabel alu1 12 44 12 44 6 b
rlabel polyct1 28 36 28 36 6 a
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 48 20 48 6 b
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 28 44 28 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 36 52 36 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 52 60 52 60 6 z
<< end >>
