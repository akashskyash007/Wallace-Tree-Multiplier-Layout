magic
tech scmos
timestamp 1199203715
<< ab >>
rect 0 0 168 80
<< nwell >>
rect -5 36 173 88
<< pwell >>
rect -5 -8 173 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 72 53 74
rect 29 69 31 72
rect 39 69 41 72
rect 51 55 53 72
rect 62 70 64 74
rect 72 70 74 74
rect 82 70 84 74
rect 92 70 94 74
rect 112 70 114 74
rect 122 70 124 74
rect 132 70 134 74
rect 48 53 54 55
rect 48 51 50 53
rect 52 51 54 53
rect 48 49 54 51
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 62 41 64 44
rect 72 41 74 44
rect 143 64 156 66
rect 143 61 145 64
rect 152 62 158 64
rect 152 60 154 62
rect 156 60 158 62
rect 152 58 158 60
rect 153 55 155 58
rect 143 42 145 46
rect 9 37 22 39
rect 29 37 41 39
rect 61 39 74 41
rect 82 39 84 42
rect 92 39 94 42
rect 112 39 114 42
rect 122 39 124 42
rect 61 37 67 39
rect 16 35 18 37
rect 20 35 22 37
rect 16 33 22 35
rect 9 28 11 33
rect 16 31 28 33
rect 16 28 18 31
rect 26 28 28 31
rect 33 28 35 37
rect 61 35 63 37
rect 65 35 67 37
rect 79 37 108 39
rect 79 35 81 37
rect 45 30 47 35
rect 55 33 67 35
rect 55 30 57 33
rect 65 30 67 33
rect 75 33 81 35
rect 102 35 104 37
rect 106 35 108 37
rect 102 33 108 35
rect 112 37 118 39
rect 112 35 114 37
rect 116 35 118 37
rect 112 33 118 35
rect 122 37 128 39
rect 122 35 124 37
rect 126 35 128 37
rect 132 38 134 42
rect 132 36 146 38
rect 122 33 128 35
rect 140 34 142 36
rect 144 34 146 36
rect 75 30 77 33
rect 85 31 91 33
rect 85 29 87 31
rect 89 29 91 31
rect 85 27 97 29
rect 85 24 87 27
rect 95 24 97 27
rect 113 24 115 33
rect 122 29 124 33
rect 140 32 146 34
rect 140 29 142 32
rect 153 30 155 42
rect 120 27 124 29
rect 120 24 122 27
rect 130 24 132 29
rect 9 8 11 16
rect 16 12 18 16
rect 26 12 28 16
rect 33 8 35 16
rect 9 6 35 8
rect 45 8 47 16
rect 55 12 57 16
rect 65 12 67 16
rect 75 8 77 16
rect 45 6 77 8
rect 85 7 87 12
rect 95 7 97 12
rect 140 12 142 16
rect 113 6 115 11
rect 120 6 122 11
rect 130 8 132 11
rect 153 8 155 19
rect 130 6 155 8
<< ndif >>
rect 37 28 45 30
rect 2 20 9 28
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 16 16 28
rect 18 26 26 28
rect 18 24 21 26
rect 23 24 26 26
rect 18 16 26 24
rect 28 16 33 28
rect 35 16 45 28
rect 47 28 55 30
rect 47 26 50 28
rect 52 26 55 28
rect 47 16 55 26
rect 57 21 65 30
rect 57 19 60 21
rect 62 19 65 21
rect 57 16 65 19
rect 67 28 75 30
rect 67 26 70 28
rect 72 26 75 28
rect 67 21 75 26
rect 67 19 70 21
rect 72 19 75 21
rect 67 16 75 19
rect 77 24 82 30
rect 148 29 153 30
rect 135 24 140 29
rect 77 20 85 24
rect 77 18 80 20
rect 82 18 85 20
rect 77 16 85 18
rect 37 11 43 16
rect 37 9 39 11
rect 41 9 43 11
rect 37 7 43 9
rect 80 12 85 16
rect 87 21 95 24
rect 87 19 90 21
rect 92 19 95 21
rect 87 12 95 19
rect 97 14 113 24
rect 97 12 104 14
rect 106 12 113 14
rect 99 11 113 12
rect 115 11 120 24
rect 122 21 130 24
rect 122 19 125 21
rect 127 19 130 21
rect 122 11 130 19
rect 132 22 140 24
rect 132 20 135 22
rect 137 20 140 22
rect 132 16 140 20
rect 142 21 153 29
rect 142 19 147 21
rect 149 19 153 21
rect 155 28 162 30
rect 155 26 158 28
rect 160 26 162 28
rect 155 24 162 26
rect 155 19 160 24
rect 142 16 151 19
rect 132 11 137 16
rect 99 9 111 11
<< pdif >>
rect 4 62 9 69
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 53 9 58
rect 2 51 4 53
rect 6 51 9 53
rect 2 49 9 51
rect 4 42 9 49
rect 11 53 19 69
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 61 29 69
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 46 39 69
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 63 46 69
rect 41 61 49 63
rect 41 59 45 61
rect 47 59 49 61
rect 41 57 49 59
rect 41 42 46 57
rect 55 68 62 70
rect 55 66 57 68
rect 59 66 62 68
rect 55 61 62 66
rect 55 59 57 61
rect 59 59 62 61
rect 55 57 62 59
rect 56 44 62 57
rect 64 60 72 70
rect 64 58 67 60
rect 69 58 72 60
rect 64 53 72 58
rect 64 51 67 53
rect 69 51 72 53
rect 64 44 72 51
rect 74 68 82 70
rect 74 66 77 68
rect 79 66 82 68
rect 74 61 82 66
rect 74 59 77 61
rect 79 59 82 61
rect 74 44 82 59
rect 77 42 82 44
rect 84 46 92 70
rect 84 44 87 46
rect 89 44 92 46
rect 84 42 92 44
rect 94 68 101 70
rect 94 66 97 68
rect 99 66 101 68
rect 94 61 101 66
rect 107 63 112 70
rect 94 59 97 61
rect 99 59 101 61
rect 94 42 101 59
rect 105 61 112 63
rect 105 59 107 61
rect 109 59 112 61
rect 105 57 112 59
rect 107 42 112 57
rect 114 54 122 70
rect 114 52 117 54
rect 119 52 122 54
rect 114 42 122 52
rect 124 53 132 70
rect 124 51 127 53
rect 129 51 132 53
rect 124 46 132 51
rect 124 44 127 46
rect 129 44 132 46
rect 124 42 132 44
rect 134 68 141 70
rect 134 66 137 68
rect 139 66 141 68
rect 134 61 141 66
rect 134 46 143 61
rect 145 55 150 61
rect 145 50 153 55
rect 145 48 148 50
rect 150 48 153 50
rect 145 46 153 48
rect 134 42 141 46
rect 148 42 153 46
rect 155 53 166 55
rect 155 51 162 53
rect 164 51 166 53
rect 155 42 166 51
<< alu1 >>
rect -2 81 170 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 170 81
rect -2 68 170 79
rect 2 61 49 62
rect 2 60 24 61
rect 2 58 4 60
rect 6 59 24 60
rect 26 59 45 61
rect 47 59 49 61
rect 6 58 49 59
rect 146 62 158 63
rect 2 53 6 58
rect 2 51 4 53
rect 2 30 6 51
rect 57 37 87 38
rect 57 35 63 37
rect 65 35 87 37
rect 57 34 87 35
rect 2 26 24 30
rect 20 24 21 26
rect 23 24 24 26
rect 81 26 87 34
rect 20 22 24 24
rect 20 21 64 22
rect 20 19 60 21
rect 62 19 64 21
rect 20 18 64 19
rect 146 60 154 62
rect 156 60 158 62
rect 146 57 158 60
rect 154 49 158 57
rect 145 33 158 39
rect 145 26 151 33
rect -2 11 170 12
rect -2 9 39 11
rect 41 9 170 11
rect -2 1 170 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 170 1
rect -2 -2 170 -1
<< ptie >>
rect 0 1 168 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 168 1
rect 0 -3 168 -1
<< ntie >>
rect 0 81 168 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 168 81
rect 0 77 168 79
<< nmos >>
rect 9 16 11 28
rect 16 16 18 28
rect 26 16 28 28
rect 33 16 35 28
rect 45 16 47 30
rect 55 16 57 30
rect 65 16 67 30
rect 75 16 77 30
rect 85 12 87 24
rect 95 12 97 24
rect 113 11 115 24
rect 120 11 122 24
rect 130 11 132 24
rect 140 16 142 29
rect 153 19 155 30
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 69
rect 62 44 64 70
rect 72 44 74 70
rect 82 42 84 70
rect 92 42 94 70
rect 112 42 114 70
rect 122 42 124 70
rect 132 42 134 70
rect 143 46 145 61
rect 153 42 155 55
<< polyct0 >>
rect 50 51 52 53
rect 18 35 20 37
rect 104 35 106 37
rect 114 35 116 37
rect 124 35 126 37
rect 142 34 144 36
rect 87 29 89 31
<< polyct1 >>
rect 154 60 156 62
rect 63 35 65 37
<< ndifct0 >>
rect 4 18 6 20
rect 50 26 52 28
rect 70 26 72 28
rect 70 19 72 21
rect 80 18 82 20
rect 90 19 92 21
rect 104 12 106 14
rect 125 19 127 21
rect 135 20 137 22
rect 147 19 149 21
rect 158 26 160 28
<< ndifct1 >>
rect 21 24 23 26
rect 60 19 62 21
rect 39 9 41 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
<< pdifct0 >>
rect 14 51 16 53
rect 14 44 16 46
rect 34 44 36 46
rect 57 66 59 68
rect 57 59 59 61
rect 67 58 69 60
rect 67 51 69 53
rect 77 66 79 68
rect 77 59 79 61
rect 87 44 89 46
rect 97 66 99 68
rect 97 59 99 61
rect 107 59 109 61
rect 117 52 119 54
rect 127 51 129 53
rect 127 44 129 46
rect 137 66 139 68
rect 148 48 150 50
rect 162 51 164 53
<< pdifct1 >>
rect 4 58 6 60
rect 4 51 6 53
rect 24 59 26 61
rect 45 59 47 61
<< alu0 >>
rect 55 66 57 68
rect 59 66 61 68
rect 55 61 61 66
rect 75 66 77 68
rect 79 66 81 68
rect 55 59 57 61
rect 59 59 61 61
rect 55 58 61 59
rect 66 60 70 62
rect 66 58 67 60
rect 69 58 70 60
rect 75 61 81 66
rect 75 59 77 61
rect 79 59 81 61
rect 75 58 81 59
rect 95 66 97 68
rect 99 66 101 68
rect 95 61 101 66
rect 135 66 137 68
rect 139 66 141 68
rect 135 65 141 66
rect 95 59 97 61
rect 99 59 101 61
rect 95 58 101 59
rect 105 61 138 62
rect 105 59 107 61
rect 109 59 138 61
rect 105 58 138 59
rect 6 49 7 58
rect 66 54 70 58
rect 115 54 121 55
rect 12 53 99 54
rect 12 51 14 53
rect 16 51 50 53
rect 52 51 67 53
rect 69 51 99 53
rect 12 50 99 51
rect 12 46 17 50
rect 12 44 14 46
rect 16 44 17 46
rect 12 42 17 44
rect 32 46 38 47
rect 85 46 91 47
rect 32 44 34 46
rect 36 44 38 46
rect 32 38 38 44
rect 48 44 87 46
rect 89 44 91 46
rect 48 42 91 44
rect 48 38 52 42
rect 16 37 52 38
rect 16 35 18 37
rect 20 35 52 37
rect 16 34 52 35
rect 48 30 52 34
rect 48 28 73 30
rect 48 26 50 28
rect 52 26 70 28
rect 72 26 73 28
rect 87 31 91 32
rect 89 29 91 31
rect 87 28 91 29
rect 48 25 54 26
rect 3 20 7 22
rect 3 18 4 20
rect 6 18 7 20
rect 69 21 73 26
rect 95 22 99 50
rect 69 19 70 21
rect 72 19 73 21
rect 3 12 7 18
rect 69 17 73 19
rect 79 20 83 22
rect 79 18 80 20
rect 82 18 83 20
rect 88 21 99 22
rect 88 19 90 21
rect 92 19 99 21
rect 88 18 99 19
rect 103 52 117 54
rect 119 52 121 54
rect 103 50 121 52
rect 126 53 130 55
rect 126 51 127 53
rect 129 51 130 53
rect 103 37 107 50
rect 126 46 130 51
rect 103 35 104 37
rect 106 35 107 37
rect 103 22 107 35
rect 113 44 127 46
rect 129 44 130 46
rect 113 42 130 44
rect 134 46 138 58
rect 147 50 151 52
rect 147 48 148 50
rect 150 48 151 50
rect 161 53 165 68
rect 161 51 162 53
rect 164 51 165 53
rect 161 49 165 51
rect 147 46 151 48
rect 134 42 166 46
rect 113 37 117 42
rect 134 38 138 42
rect 113 35 114 37
rect 116 35 117 37
rect 113 30 117 35
rect 122 37 138 38
rect 122 35 124 37
rect 126 35 138 37
rect 122 34 138 35
rect 141 36 145 38
rect 141 34 142 36
rect 144 34 145 36
rect 141 32 145 34
rect 113 26 138 30
rect 162 29 166 42
rect 156 28 166 29
rect 156 26 158 28
rect 160 26 166 28
rect 134 22 138 26
rect 156 25 166 26
rect 103 21 129 22
rect 103 19 125 21
rect 127 19 129 21
rect 103 18 129 19
rect 134 20 135 22
rect 137 20 138 22
rect 134 18 138 20
rect 145 21 151 22
rect 145 19 147 21
rect 149 19 151 21
rect 79 12 83 18
rect 102 14 108 15
rect 102 12 104 14
rect 106 12 108 14
rect 145 12 151 19
<< labels >>
rlabel alu0 14 48 14 48 6 cn
rlabel alu0 35 40 35 40 6 zn
rlabel alu0 60 28 60 28 6 zn
rlabel alu0 71 23 71 23 6 zn
rlabel alu0 93 20 93 20 6 cn
rlabel alu0 69 44 69 44 6 zn
rlabel alu0 68 56 68 56 6 cn
rlabel alu0 55 52 55 52 6 cn
rlabel alu0 116 20 116 20 6 iz
rlabel polyct0 115 36 115 36 6 an
rlabel alu0 128 48 128 48 6 an
rlabel alu0 118 52 118 52 6 iz
rlabel polyct0 105 36 105 36 6 iz
rlabel alu0 136 24 136 24 6 an
rlabel alu0 161 27 161 27 6 bn
rlabel alu0 130 36 130 36 6 bn
rlabel alu0 149 47 149 47 6 bn
rlabel alu0 121 60 121 60 6 bn
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 20 28 20 28 6 z
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 44 20 44 20 6 z
rlabel alu1 76 36 76 36 6 c
rlabel alu1 68 36 68 36 6 c
rlabel alu1 60 36 60 36 6 c
rlabel alu1 44 60 44 60 6 z
rlabel alu1 84 6 84 6 6 vss
rlabel alu1 84 32 84 32 6 c
rlabel alu1 84 74 84 74 6 vdd
rlabel alu1 156 36 156 36 6 a
rlabel alu1 148 32 148 32 6 a
rlabel alu1 156 56 156 56 6 b
rlabel alu1 148 60 148 60 6 b
<< end >>
