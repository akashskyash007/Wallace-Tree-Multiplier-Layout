magic
tech scmos
timestamp 1199201792
<< ab >>
rect 0 0 88 72
<< nwell >>
rect -5 32 93 77
<< pwell >>
rect -5 -5 93 32
<< poly >>
rect 9 66 11 70
rect 16 66 18 70
rect 26 66 28 70
rect 33 66 35 70
rect 43 66 45 70
rect 53 66 55 70
rect 63 66 65 70
rect 73 66 75 70
rect 9 29 11 38
rect 16 35 18 38
rect 26 35 28 38
rect 16 33 28 35
rect 20 31 24 33
rect 26 31 28 33
rect 20 29 28 31
rect 9 27 15 29
rect 9 25 11 27
rect 13 25 15 27
rect 9 23 15 25
rect 10 20 12 23
rect 20 20 22 29
rect 33 27 35 38
rect 43 35 45 38
rect 53 35 55 38
rect 63 35 65 38
rect 43 33 49 35
rect 43 31 45 33
rect 47 31 49 33
rect 43 29 49 31
rect 53 33 65 35
rect 73 35 75 38
rect 73 33 79 35
rect 53 31 55 33
rect 57 31 59 33
rect 53 29 59 31
rect 73 31 75 33
rect 77 31 79 33
rect 73 29 79 31
rect 33 25 39 27
rect 47 26 49 29
rect 54 26 56 29
rect 33 23 35 25
rect 37 23 39 25
rect 33 21 39 23
rect 10 5 12 10
rect 20 5 22 10
rect 47 4 49 9
rect 54 4 56 9
<< ndif >>
rect 2 10 10 20
rect 12 17 20 20
rect 12 15 15 17
rect 17 15 20 17
rect 12 10 20 15
rect 22 10 31 20
rect 42 19 47 26
rect 40 17 47 19
rect 40 15 42 17
rect 44 15 47 17
rect 40 13 47 15
rect 2 7 8 10
rect 2 5 4 7
rect 6 5 8 7
rect 24 7 31 10
rect 42 9 47 13
rect 49 9 54 26
rect 56 20 63 26
rect 56 18 59 20
rect 61 18 63 20
rect 56 13 63 18
rect 56 11 59 13
rect 61 11 63 13
rect 56 9 63 11
rect 24 5 26 7
rect 28 5 31 7
rect 2 3 8 5
rect 24 3 31 5
<< pdif >>
rect 4 60 9 66
rect 2 58 9 60
rect 2 56 4 58
rect 6 56 9 58
rect 2 54 9 56
rect 4 38 9 54
rect 11 38 16 66
rect 18 50 26 66
rect 18 48 21 50
rect 23 48 26 50
rect 18 43 26 48
rect 18 41 21 43
rect 23 41 26 43
rect 18 38 26 41
rect 28 38 33 66
rect 35 57 43 66
rect 35 55 38 57
rect 40 55 43 57
rect 35 50 43 55
rect 35 48 38 50
rect 40 48 43 50
rect 35 38 43 48
rect 45 64 53 66
rect 45 62 48 64
rect 50 62 53 64
rect 45 57 53 62
rect 45 55 48 57
rect 50 55 53 57
rect 45 38 53 55
rect 55 56 63 66
rect 55 54 58 56
rect 60 54 63 56
rect 55 49 63 54
rect 55 47 58 49
rect 60 47 63 49
rect 55 38 63 47
rect 65 64 73 66
rect 65 62 68 64
rect 70 62 73 64
rect 65 57 73 62
rect 65 55 68 57
rect 70 55 73 57
rect 65 38 73 55
rect 75 59 80 66
rect 75 57 82 59
rect 75 55 78 57
rect 80 55 82 57
rect 75 50 82 55
rect 75 48 78 50
rect 80 48 82 50
rect 75 46 82 48
rect 75 38 80 46
<< alu1 >>
rect -2 64 90 72
rect 2 50 25 51
rect 2 48 21 50
rect 23 48 25 50
rect 2 47 25 48
rect 2 18 6 47
rect 18 46 25 47
rect 19 43 25 46
rect 10 27 14 43
rect 19 41 21 43
rect 23 41 25 43
rect 19 40 25 41
rect 33 34 39 42
rect 22 33 39 34
rect 22 31 24 33
rect 26 31 39 33
rect 22 30 39 31
rect 43 38 78 42
rect 43 33 49 38
rect 43 31 45 33
rect 47 31 49 33
rect 43 30 49 31
rect 53 33 70 34
rect 53 31 55 33
rect 57 31 70 33
rect 53 30 70 31
rect 10 25 11 27
rect 13 26 14 27
rect 13 25 39 26
rect 10 23 35 25
rect 37 23 39 25
rect 10 22 39 23
rect 2 17 47 18
rect 2 15 15 17
rect 17 15 42 17
rect 44 15 47 17
rect 2 14 47 15
rect 66 13 70 30
rect 74 33 78 38
rect 74 31 75 33
rect 77 31 78 33
rect 74 21 78 31
rect -2 7 90 8
rect -2 5 4 7
rect 6 5 26 7
rect 28 5 69 7
rect 71 5 77 7
rect 79 5 90 7
rect -2 0 90 5
<< ptie >>
rect 67 7 81 9
rect 67 5 69 7
rect 71 5 77 7
rect 79 5 81 7
rect 67 3 81 5
<< nmos >>
rect 10 10 12 20
rect 20 10 22 20
rect 47 9 49 26
rect 54 9 56 26
<< pmos >>
rect 9 38 11 66
rect 16 38 18 66
rect 26 38 28 66
rect 33 38 35 66
rect 43 38 45 66
rect 53 38 55 66
rect 63 38 65 66
rect 73 38 75 66
<< polyct1 >>
rect 24 31 26 33
rect 11 25 13 27
rect 45 31 47 33
rect 55 31 57 33
rect 75 31 77 33
rect 35 23 37 25
<< ndifct0 >>
rect 59 18 61 20
rect 59 11 61 13
<< ndifct1 >>
rect 15 15 17 17
rect 42 15 44 17
rect 4 5 6 7
rect 26 5 28 7
<< ptiect1 >>
rect 69 5 71 7
rect 77 5 79 7
<< pdifct0 >>
rect 4 56 6 58
rect 38 55 40 57
rect 38 48 40 50
rect 48 62 50 64
rect 48 55 50 57
rect 58 54 60 56
rect 58 47 60 49
rect 68 62 70 64
rect 68 55 70 57
rect 78 55 80 57
rect 78 48 80 50
<< pdifct1 >>
rect 21 48 23 50
rect 21 41 23 43
<< alu0 >>
rect 46 62 48 64
rect 50 62 52 64
rect 2 58 41 59
rect 2 56 4 58
rect 6 57 41 58
rect 6 56 38 57
rect 2 55 38 56
rect 40 55 41 57
rect 6 46 18 47
rect 37 50 41 55
rect 46 57 52 62
rect 66 62 68 64
rect 70 62 72 64
rect 46 55 48 57
rect 50 55 52 57
rect 46 54 52 55
rect 57 56 61 58
rect 57 54 58 56
rect 60 54 61 56
rect 66 57 72 62
rect 66 55 68 57
rect 70 55 72 57
rect 66 54 72 55
rect 77 57 81 59
rect 77 55 78 57
rect 80 55 81 57
rect 57 50 61 54
rect 77 50 81 55
rect 37 48 38 50
rect 40 49 78 50
rect 40 48 58 49
rect 37 47 58 48
rect 60 48 78 49
rect 80 48 81 50
rect 60 47 81 48
rect 37 46 81 47
rect 58 20 62 22
rect 58 18 59 20
rect 61 18 62 20
rect 58 13 62 18
rect 58 11 59 13
rect 61 11 62 13
rect 58 8 62 11
<< labels >>
rlabel alu0 39 52 39 52 6 n1
rlabel alu0 21 57 21 57 6 n1
rlabel alu0 79 52 79 52 6 n1
rlabel alu0 59 52 59 52 6 n1
rlabel alu1 12 16 12 16 6 z
rlabel alu1 12 36 12 36 6 b
rlabel alu1 4 36 4 36 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 24 20 24 6 b
rlabel polyct1 36 24 36 24 6 b
rlabel alu1 28 32 28 32 6 c
rlabel alu1 28 24 28 24 6 b
rlabel alu1 36 36 36 36 6 c
rlabel alu1 20 48 20 48 6 z
rlabel alu1 44 4 44 4 6 vss
rlabel alu1 44 16 44 16 6 z
rlabel alu1 60 32 60 32 6 a1
rlabel alu1 52 40 52 40 6 a2
rlabel alu1 60 40 60 40 6 a2
rlabel alu1 44 68 44 68 6 vdd
rlabel alu1 68 20 68 20 6 a1
rlabel alu1 76 28 76 28 6 a2
rlabel alu1 68 40 68 40 6 a2
<< end >>
