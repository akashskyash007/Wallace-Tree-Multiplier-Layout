magic
tech scmos
timestamp 1199469589
<< ab >>
rect 0 0 30 100
<< nwell >>
rect -5 48 35 105
<< pwell >>
rect -5 -5 35 48
<< poly >>
rect 15 75 17 80
rect 15 50 17 55
rect 15 48 23 50
rect 15 46 19 48
rect 21 46 23 48
rect 15 44 23 46
rect 15 33 17 44
rect 15 18 17 23
<< ndif >>
rect 7 31 15 33
rect 7 29 9 31
rect 11 29 15 31
rect 7 27 15 29
rect 10 23 15 27
rect 17 23 26 33
rect 19 21 26 23
rect 19 19 21 21
rect 23 19 26 21
rect 19 17 26 19
<< pdif >>
rect 10 71 15 75
rect 7 69 15 71
rect 7 67 9 69
rect 11 67 15 69
rect 7 61 15 67
rect 7 59 9 61
rect 11 59 15 61
rect 7 57 15 59
rect 10 55 15 57
rect 17 71 26 75
rect 17 69 21 71
rect 23 69 26 71
rect 17 55 26 69
<< alu1 >>
rect -2 95 32 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 32 95
rect -2 88 32 93
rect 8 69 12 73
rect 8 67 9 69
rect 11 67 12 69
rect 20 71 24 88
rect 20 69 21 71
rect 23 69 24 71
rect 20 67 24 69
rect 8 61 12 67
rect 8 59 9 61
rect 11 59 12 61
rect 8 32 12 59
rect 18 48 22 63
rect 18 46 19 48
rect 21 46 22 48
rect 18 37 22 46
rect 8 31 23 32
rect 8 29 9 31
rect 11 29 23 31
rect 8 27 23 29
rect 20 21 24 23
rect 20 19 21 21
rect 23 19 24 21
rect 20 12 24 19
rect -2 7 32 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 32 7
rect -2 0 32 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 15 23 17 33
<< pmos >>
rect 15 55 17 75
<< polyct1 >>
rect 19 46 21 48
<< ndifct1 >>
rect 9 29 11 31
rect 21 19 23 21
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 9 67 11 69
rect 9 59 11 61
rect 21 69 23 71
<< labels >>
rlabel alu1 15 6 15 6 6 vss
rlabel alu1 10 50 10 50 6 z
rlabel alu1 15 94 15 94 6 vdd
rlabel alu1 20 30 20 30 6 z
rlabel alu1 20 50 20 50 6 a
<< end >>
