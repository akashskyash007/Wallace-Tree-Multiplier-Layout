magic
tech scmos
timestamp 1199543315
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 45 95 47 98
rect 57 95 59 98
rect 11 85 13 88
rect 19 85 21 88
rect 27 85 29 88
rect 11 33 13 55
rect 19 43 21 55
rect 27 53 29 55
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 7 31 13 33
rect 7 29 9 31
rect 11 29 13 31
rect 7 27 13 29
rect 19 29 21 37
rect 31 29 33 47
rect 45 43 47 55
rect 57 43 59 55
rect 37 41 59 43
rect 37 39 39 41
rect 41 39 59 41
rect 37 37 59 39
rect 19 27 25 29
rect 31 27 37 29
rect 11 25 13 27
rect 23 25 25 27
rect 35 25 37 27
rect 45 25 47 37
rect 57 25 59 37
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 45 2 47 5
rect 57 2 59 5
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 15 35 19
rect 37 15 45 25
rect 15 11 21 15
rect 15 9 17 11
rect 19 9 21 11
rect 39 9 45 15
rect 15 7 21 9
rect 37 7 45 9
rect 37 5 39 7
rect 41 5 45 7
rect 47 21 57 25
rect 47 19 51 21
rect 53 19 57 21
rect 47 5 57 19
rect 59 21 67 25
rect 59 19 63 21
rect 65 19 67 21
rect 59 11 67 19
rect 59 9 63 11
rect 65 9 67 11
rect 59 5 67 9
rect 37 3 43 5
<< pdif >>
rect 31 91 45 95
rect 31 89 39 91
rect 41 89 45 91
rect 31 85 45 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 55 19 85
rect 21 55 27 85
rect 29 55 45 85
rect 47 81 57 95
rect 47 79 51 81
rect 53 79 57 81
rect 47 71 57 79
rect 47 69 51 71
rect 53 69 57 71
rect 47 61 57 69
rect 47 59 51 61
rect 53 59 57 61
rect 47 55 57 59
rect 59 91 67 95
rect 59 89 63 91
rect 65 89 67 91
rect 59 81 67 89
rect 59 79 63 81
rect 65 79 67 81
rect 59 71 67 79
rect 59 69 63 71
rect 65 69 67 71
rect 59 61 67 69
rect 59 59 63 61
rect 65 59 67 61
rect 59 55 67 59
<< alu1 >>
rect -2 95 72 100
rect -2 93 5 95
rect 7 93 21 95
rect 23 93 72 95
rect -2 91 72 93
rect -2 89 39 91
rect 41 89 63 91
rect 65 89 72 91
rect -2 88 72 89
rect 4 81 8 82
rect 48 81 54 82
rect 4 79 5 81
rect 7 79 41 81
rect 4 78 8 79
rect 8 31 12 72
rect 8 29 9 31
rect 11 29 12 31
rect 8 28 12 29
rect 18 41 22 72
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 28 51 32 72
rect 28 49 29 51
rect 31 49 32 51
rect 28 28 32 49
rect 39 42 41 79
rect 48 79 51 81
rect 53 79 54 81
rect 48 78 54 79
rect 62 81 66 88
rect 62 79 63 81
rect 65 79 66 81
rect 48 72 52 78
rect 48 71 54 72
rect 48 69 51 71
rect 53 69 54 71
rect 48 68 54 69
rect 62 71 66 79
rect 62 69 63 71
rect 65 69 66 71
rect 48 62 52 68
rect 48 61 54 62
rect 48 59 51 61
rect 53 59 54 61
rect 48 58 54 59
rect 62 61 66 69
rect 62 59 63 61
rect 65 59 66 61
rect 62 58 66 59
rect 38 41 42 42
rect 38 39 39 41
rect 41 39 42 41
rect 38 38 42 39
rect 4 21 8 22
rect 28 21 32 22
rect 39 21 41 38
rect 4 19 5 21
rect 7 19 29 21
rect 31 19 41 21
rect 48 22 52 58
rect 48 21 54 22
rect 48 19 51 21
rect 53 19 54 21
rect 4 18 8 19
rect 28 18 32 19
rect 48 18 54 19
rect 62 21 66 22
rect 62 19 63 21
rect 65 19 66 21
rect 62 12 66 19
rect -2 11 72 12
rect -2 9 17 11
rect 19 9 63 11
rect 65 9 72 11
rect -2 7 72 9
rect -2 5 39 7
rect 41 5 72 7
rect -2 0 72 5
<< ntie >>
rect 3 95 25 97
rect 3 93 5 95
rect 7 93 21 95
rect 23 93 25 95
rect 3 91 25 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 45 5 47 25
rect 57 5 59 25
<< pmos >>
rect 11 55 13 85
rect 19 55 21 85
rect 27 55 29 85
rect 45 55 47 95
rect 57 55 59 95
<< polyct1 >>
rect 29 49 31 51
rect 19 39 21 41
rect 9 29 11 31
rect 39 39 41 41
<< ndifct1 >>
rect 5 19 7 21
rect 29 19 31 21
rect 17 9 19 11
rect 39 5 41 7
rect 51 19 53 21
rect 63 19 65 21
rect 63 9 65 11
<< ntiect1 >>
rect 5 93 7 95
rect 21 93 23 95
<< pdifct1 >>
rect 39 89 41 91
rect 5 79 7 81
rect 51 79 53 81
rect 51 69 53 71
rect 51 59 53 61
rect 63 89 65 91
rect 63 79 65 81
rect 63 69 65 71
rect 63 59 65 61
<< labels >>
rlabel alu1 10 50 10 50 6 i2
rlabel polyct1 30 50 30 50 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 50 50 50 50 6 q
rlabel alu1 35 94 35 94 6 vdd
<< end >>
