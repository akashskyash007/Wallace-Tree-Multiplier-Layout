magic
tech scmos
timestamp 1199203103
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 12 66 14 71
rect 22 66 24 71
rect 29 66 31 71
rect 12 49 14 58
rect 9 47 15 49
rect 9 45 11 47
rect 13 45 15 47
rect 9 43 15 45
rect 9 30 11 43
rect 22 39 24 50
rect 18 37 24 39
rect 18 35 20 37
rect 22 35 24 37
rect 18 33 24 35
rect 29 47 31 50
rect 29 45 35 47
rect 29 43 31 45
rect 33 43 35 45
rect 29 41 35 43
rect 19 30 21 33
rect 9 18 11 23
rect 19 18 21 23
rect 29 22 31 41
rect 29 10 31 15
<< ndif >>
rect 2 27 9 30
rect 2 25 4 27
rect 6 25 9 27
rect 2 23 9 25
rect 11 27 19 30
rect 11 25 14 27
rect 16 25 19 27
rect 11 23 19 25
rect 21 23 27 30
rect 23 22 27 23
rect 23 16 29 22
rect 21 15 29 16
rect 31 20 38 22
rect 31 18 34 20
rect 36 18 38 20
rect 31 15 38 18
rect 21 11 27 15
rect 21 9 23 11
rect 25 9 27 11
rect 21 7 27 9
<< pdif >>
rect 3 71 10 73
rect 3 69 6 71
rect 8 69 10 71
rect 3 66 10 69
rect 3 58 12 66
rect 14 62 22 66
rect 14 60 17 62
rect 19 60 22 62
rect 14 58 22 60
rect 17 50 22 58
rect 24 50 29 66
rect 31 62 38 66
rect 31 60 34 62
rect 36 60 38 62
rect 31 50 38 60
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 71 42 79
rect -2 69 6 71
rect 8 69 42 71
rect -2 68 42 69
rect 2 62 23 63
rect 2 60 17 62
rect 19 60 23 62
rect 2 58 23 60
rect 2 27 6 58
rect 10 50 23 54
rect 10 47 14 50
rect 10 45 11 47
rect 13 45 14 47
rect 34 46 38 55
rect 10 33 14 45
rect 25 45 38 46
rect 25 43 31 45
rect 33 43 38 45
rect 25 42 38 43
rect 18 37 31 38
rect 18 35 20 37
rect 22 35 31 37
rect 18 34 31 35
rect 25 31 31 34
rect 2 25 4 27
rect 2 17 6 25
rect 25 25 38 31
rect -2 11 42 12
rect -2 9 23 11
rect 25 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 23 11 30
rect 19 23 21 30
rect 29 15 31 22
<< pmos >>
rect 12 58 14 66
rect 22 50 24 66
rect 29 50 31 66
<< polyct1 >>
rect 11 45 13 47
rect 20 35 22 37
rect 31 43 33 45
<< ndifct0 >>
rect 14 25 16 27
rect 34 18 36 20
<< ndifct1 >>
rect 4 25 6 27
rect 23 9 25 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 34 60 36 62
<< pdifct1 >>
rect 6 69 8 71
rect 17 60 19 62
<< alu0 >>
rect 32 62 38 68
rect 32 60 34 62
rect 36 60 38 62
rect 32 59 38 60
rect 6 23 7 29
rect 13 27 17 29
rect 13 25 14 27
rect 16 25 17 27
rect 13 21 17 25
rect 13 20 38 21
rect 13 18 34 20
rect 36 18 38 20
rect 13 17 38 18
<< labels >>
rlabel alu0 15 23 15 23 6 n1
rlabel alu0 25 19 25 19 6 n1
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 28 32 28 32 6 a2
rlabel alu1 28 44 28 44 6 a1
rlabel alu1 20 52 20 52 6 b
rlabel alu1 20 60 20 60 6 z
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 36 52 36 52 6 a1
<< end >>
