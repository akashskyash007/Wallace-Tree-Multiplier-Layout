magic
tech scmos
timestamp 1199202032
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 19 65 21 70
rect 29 65 31 70
rect 9 61 11 65
rect 9 39 11 43
rect 19 39 21 43
rect 9 37 21 39
rect 9 35 16 37
rect 18 36 21 37
rect 18 35 20 36
rect 9 33 20 35
rect 9 30 11 33
rect 29 32 31 43
rect 24 30 31 32
rect 24 28 26 30
rect 28 28 31 30
rect 24 26 31 28
rect 29 23 31 26
rect 9 6 11 10
rect 29 7 31 12
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 23 22 30
rect 11 21 29 23
rect 11 19 17 21
rect 19 19 29 21
rect 11 14 29 19
rect 11 12 17 14
rect 19 12 29 14
rect 31 21 38 23
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
rect 31 12 36 17
rect 11 10 27 12
<< pdif >>
rect 14 61 19 65
rect 2 59 9 61
rect 2 57 4 59
rect 6 57 9 59
rect 2 52 9 57
rect 2 50 4 52
rect 6 50 9 52
rect 2 43 9 50
rect 11 54 19 61
rect 11 52 14 54
rect 16 52 19 54
rect 11 47 19 52
rect 11 45 14 47
rect 16 45 19 47
rect 11 43 19 45
rect 21 63 29 65
rect 21 61 24 63
rect 26 61 29 63
rect 21 56 29 61
rect 21 54 24 56
rect 26 54 29 56
rect 21 43 29 54
rect 31 56 36 65
rect 31 54 38 56
rect 31 52 34 54
rect 36 52 38 54
rect 31 47 38 52
rect 31 45 34 47
rect 36 45 38 47
rect 31 43 38 45
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 13 54 17 56
rect 13 52 14 54
rect 16 52 17 54
rect 13 47 17 52
rect 13 46 14 47
rect 2 45 14 46
rect 16 46 17 47
rect 16 45 23 46
rect 2 42 23 45
rect 2 30 6 42
rect 17 30 30 31
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 17 28 26 30
rect 28 28 30 30
rect 17 26 30 28
rect 2 21 7 26
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect 26 17 30 26
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 10 11 30
rect 29 12 31 23
<< pmos >>
rect 9 43 11 61
rect 19 43 21 65
rect 29 43 31 65
<< polyct0 >>
rect 16 35 18 37
<< polyct1 >>
rect 26 28 28 30
<< ndifct0 >>
rect 17 19 19 21
rect 17 12 19 14
rect 34 19 36 21
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 4 57 6 59
rect 4 50 6 52
rect 24 61 26 63
rect 24 54 26 56
rect 34 52 36 54
rect 34 45 36 47
<< pdifct1 >>
rect 14 52 16 54
rect 14 45 16 47
<< alu0 >>
rect 2 59 8 68
rect 2 57 4 59
rect 6 57 8 59
rect 2 52 8 57
rect 23 63 27 68
rect 23 61 24 63
rect 26 61 27 63
rect 23 56 27 61
rect 2 50 4 52
rect 6 50 8 52
rect 2 49 8 50
rect 23 54 24 56
rect 26 54 27 56
rect 23 52 27 54
rect 33 54 37 56
rect 33 52 34 54
rect 36 52 37 54
rect 33 47 37 52
rect 33 45 34 47
rect 36 45 37 47
rect 33 38 37 45
rect 14 37 37 38
rect 14 35 16 37
rect 18 35 37 37
rect 14 34 37 35
rect 15 21 21 22
rect 15 19 17 21
rect 19 19 21 21
rect 15 14 21 19
rect 33 21 37 34
rect 33 19 34 21
rect 36 19 37 21
rect 33 17 37 19
rect 15 12 17 14
rect 19 12 21 14
<< labels >>
rlabel alu0 25 36 25 36 6 an
rlabel alu0 35 36 35 36 6 an
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 28 20 28 6 a
rlabel alu1 28 24 28 24 6 a
rlabel alu1 20 44 20 44 6 z
rlabel alu1 20 74 20 74 6 vdd
<< end >>
