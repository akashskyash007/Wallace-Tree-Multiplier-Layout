magic
tech scmos
timestamp 1199470161
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -5 48 95 105
<< pwell >>
rect -5 -5 95 48
<< poly >>
rect 17 94 19 98
rect 25 94 27 98
rect 33 94 35 98
rect 41 94 43 98
rect 53 94 55 98
rect 61 94 63 98
rect 69 94 71 98
rect 77 94 79 98
rect 17 52 19 55
rect 7 50 19 52
rect 7 48 9 50
rect 11 48 15 50
rect 7 46 15 48
rect 13 24 15 46
rect 25 33 27 55
rect 33 42 35 55
rect 41 52 43 55
rect 53 52 55 55
rect 41 50 55 52
rect 45 48 47 50
rect 49 48 51 50
rect 45 46 51 48
rect 33 40 43 42
rect 37 38 39 40
rect 41 38 43 40
rect 37 36 43 38
rect 25 31 33 33
rect 25 29 29 31
rect 31 29 33 31
rect 25 27 33 29
rect 25 24 27 27
rect 37 24 39 36
rect 49 24 51 46
rect 61 43 63 55
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 69 33 71 55
rect 77 52 79 55
rect 77 50 83 52
rect 77 48 79 50
rect 81 48 83 50
rect 77 46 83 48
rect 65 31 71 33
rect 65 29 67 31
rect 69 29 71 31
rect 65 27 71 29
rect 13 8 15 13
rect 25 8 27 13
rect 37 8 39 13
rect 49 8 51 13
<< ndif >>
rect 4 21 13 24
rect 4 19 7 21
rect 9 19 13 21
rect 4 13 13 19
rect 15 21 25 24
rect 15 19 19 21
rect 21 19 25 21
rect 15 13 25 19
rect 27 13 37 24
rect 39 21 49 24
rect 39 19 43 21
rect 45 19 49 21
rect 39 13 49 19
rect 51 21 60 24
rect 51 19 55 21
rect 57 19 60 21
rect 51 13 60 19
rect 29 11 35 13
rect 29 9 31 11
rect 33 9 35 11
rect 29 7 35 9
<< pdif >>
rect 9 91 17 94
rect 9 89 11 91
rect 13 89 17 91
rect 9 55 17 89
rect 19 55 25 94
rect 27 55 33 94
rect 35 55 41 94
rect 43 71 53 94
rect 43 69 47 71
rect 49 69 53 71
rect 43 61 53 69
rect 43 59 47 61
rect 49 59 53 61
rect 43 55 53 59
rect 55 55 61 94
rect 63 55 69 94
rect 71 55 77 94
rect 79 91 87 94
rect 79 89 83 91
rect 85 89 87 91
rect 79 81 87 89
rect 79 79 83 81
rect 85 79 87 81
rect 79 71 87 79
rect 79 69 83 71
rect 85 69 87 71
rect 79 55 87 69
<< alu1 >>
rect -2 91 92 100
rect -2 89 11 91
rect 13 89 83 91
rect 85 89 92 91
rect -2 88 92 89
rect 7 78 73 82
rect 7 50 12 78
rect 7 48 9 50
rect 11 48 12 50
rect 7 46 12 48
rect 18 71 52 73
rect 18 69 47 71
rect 49 69 52 71
rect 18 68 52 69
rect 6 21 10 23
rect 6 19 7 21
rect 9 19 10 21
rect 6 12 10 19
rect 18 22 22 68
rect 28 52 32 63
rect 46 61 52 68
rect 46 59 47 61
rect 49 59 52 61
rect 46 57 52 59
rect 28 50 53 52
rect 28 48 47 50
rect 49 48 53 50
rect 28 47 53 48
rect 28 37 32 47
rect 58 42 62 63
rect 68 52 73 78
rect 82 81 86 88
rect 82 79 83 81
rect 85 79 86 81
rect 82 71 86 79
rect 82 69 83 71
rect 85 69 86 71
rect 82 67 86 69
rect 68 50 83 52
rect 68 48 79 50
rect 81 48 83 50
rect 68 47 83 48
rect 37 41 62 42
rect 37 40 59 41
rect 37 38 39 40
rect 41 39 59 40
rect 61 39 62 41
rect 41 38 62 39
rect 37 37 62 38
rect 68 32 72 43
rect 27 31 72 32
rect 27 29 29 31
rect 31 29 67 31
rect 69 29 72 31
rect 27 28 72 29
rect 18 21 47 22
rect 18 19 19 21
rect 21 19 43 21
rect 45 19 47 21
rect 18 17 47 19
rect 54 21 58 23
rect 54 19 55 21
rect 57 19 58 21
rect 54 12 58 19
rect 68 17 72 28
rect -2 11 92 12
rect -2 9 31 11
rect 33 9 92 11
rect -2 7 92 9
rect -2 5 69 7
rect 71 5 79 7
rect 81 5 92 7
rect -2 0 92 5
<< ptie >>
rect 67 7 83 9
rect 67 5 69 7
rect 71 5 79 7
rect 81 5 83 7
rect 67 3 83 5
<< nmos >>
rect 13 13 15 24
rect 25 13 27 24
rect 37 13 39 24
rect 49 13 51 24
<< pmos >>
rect 17 55 19 94
rect 25 55 27 94
rect 33 55 35 94
rect 41 55 43 94
rect 53 55 55 94
rect 61 55 63 94
rect 69 55 71 94
rect 77 55 79 94
<< polyct1 >>
rect 9 48 11 50
rect 47 48 49 50
rect 39 38 41 40
rect 29 29 31 31
rect 59 39 61 41
rect 79 48 81 50
rect 67 29 69 31
<< ndifct1 >>
rect 7 19 9 21
rect 19 19 21 21
rect 43 19 45 21
rect 55 19 57 21
rect 31 9 33 11
<< ptiect1 >>
rect 69 5 71 7
rect 79 5 81 7
<< pdifct1 >>
rect 11 89 13 91
rect 47 69 49 71
rect 47 59 49 61
rect 83 89 85 91
rect 83 79 85 81
rect 83 69 85 71
<< labels >>
rlabel alu1 10 65 10 65 6 d
rlabel alu1 30 20 30 20 6 z
rlabel polyct1 30 30 30 30 6 b
rlabel alu1 20 45 20 45 6 z
rlabel alu1 30 50 30 50 6 a
rlabel alu1 30 70 30 70 6 z
rlabel alu1 30 80 30 80 6 d
rlabel alu1 20 80 20 80 6 d
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 40 20 40 20 6 z
rlabel alu1 40 30 40 30 6 b
rlabel alu1 50 30 50 30 6 b
rlabel alu1 50 40 50 40 6 c
rlabel alu1 40 40 40 40 6 c
rlabel alu1 50 50 50 50 6 a
rlabel alu1 40 50 40 50 6 a
rlabel alu1 40 70 40 70 6 z
rlabel alu1 50 65 50 65 6 z
rlabel alu1 50 80 50 80 6 d
rlabel alu1 40 80 40 80 6 d
rlabel alu1 45 94 45 94 6 vdd
rlabel alu1 70 30 70 30 6 b
rlabel alu1 60 30 60 30 6 b
rlabel alu1 60 50 60 50 6 c
rlabel alu1 70 65 70 65 6 d
rlabel alu1 60 80 60 80 6 d
rlabel alu1 80 50 80 50 6 d
<< end >>
