magic
tech scmos
timestamp 1199973047
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -5 40 101 97
<< pwell >>
rect -5 -9 101 40
<< poly >>
rect 2 77 11 83
rect 9 74 11 77
rect 21 77 30 83
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 77 75 83
rect 53 74 55 77
rect 73 74 75 77
rect 85 81 94 83
rect 85 79 87 81
rect 89 79 94 81
rect 85 77 94 79
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 41 14 43
rect 2 39 7 41
rect 9 39 14 41
rect 2 37 14 39
rect 18 41 30 43
rect 18 39 23 41
rect 25 39 30 41
rect 18 37 30 39
rect 34 41 46 43
rect 34 39 39 41
rect 41 39 46 41
rect 34 37 46 39
rect 50 41 62 43
rect 50 39 55 41
rect 57 39 62 41
rect 50 37 62 39
rect 66 41 78 43
rect 66 39 71 41
rect 73 39 78 41
rect 66 37 78 39
rect 82 37 94 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 5 62 11
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndif >>
rect 2 27 9 34
rect 2 25 4 27
rect 6 25 9 27
rect 2 20 9 25
rect 2 18 4 20
rect 6 18 9 20
rect 2 14 9 18
rect 11 14 21 34
rect 23 29 30 34
rect 23 27 26 29
rect 28 27 30 29
rect 23 14 30 27
rect 34 28 41 34
rect 34 26 36 28
rect 38 26 41 28
rect 34 21 41 26
rect 34 19 36 21
rect 38 19 41 21
rect 34 14 41 19
rect 43 32 53 34
rect 43 30 47 32
rect 49 30 53 32
rect 43 14 53 30
rect 55 18 62 34
rect 55 16 58 18
rect 60 16 62 18
rect 55 14 62 16
rect 66 32 73 34
rect 66 30 68 32
rect 70 30 73 32
rect 66 25 73 30
rect 66 23 68 25
rect 70 23 73 25
rect 66 14 73 23
rect 75 25 85 34
rect 75 23 79 25
rect 81 23 85 25
rect 75 17 85 23
rect 75 15 79 17
rect 81 15 85 17
rect 75 14 85 15
rect 87 14 94 34
rect 13 12 15 14
rect 17 12 19 14
rect 13 6 19 12
rect 13 4 15 6
rect 17 4 19 6
rect 13 2 19 4
rect 45 2 51 14
rect 77 2 83 14
<< pdif >>
rect 13 84 19 86
rect 13 82 15 84
rect 17 82 19 84
rect 13 76 19 82
rect 13 74 15 76
rect 17 74 19 76
rect 45 74 51 86
rect 77 74 83 86
rect 2 68 9 74
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 46 9 59
rect 11 46 21 74
rect 23 61 30 74
rect 23 59 26 61
rect 28 59 30 61
rect 23 46 30 59
rect 34 72 41 74
rect 34 70 36 72
rect 38 70 41 72
rect 34 46 41 70
rect 43 50 53 74
rect 43 48 47 50
rect 49 48 53 50
rect 43 46 53 48
rect 55 72 62 74
rect 55 70 58 72
rect 60 70 62 72
rect 55 65 62 70
rect 55 63 58 65
rect 60 63 62 65
rect 55 46 62 63
rect 66 65 73 74
rect 66 63 68 65
rect 70 63 73 65
rect 66 58 73 63
rect 66 56 68 58
rect 70 56 73 58
rect 66 46 73 56
rect 75 73 85 74
rect 75 71 79 73
rect 81 71 85 73
rect 75 66 85 71
rect 75 64 79 66
rect 81 64 85 66
rect 75 46 85 64
rect 87 46 94 74
<< alu1 >>
rect -2 89 98 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 73 87 87 89
rect 89 87 91 89
rect 93 87 98 89
rect -2 86 98 87
rect 14 84 18 86
rect 14 82 15 84
rect 17 82 18 84
rect 14 81 18 82
rect 14 79 15 81
rect 17 79 18 81
rect 14 76 18 79
rect 14 74 15 76
rect 17 74 18 76
rect 14 72 18 74
rect 78 81 82 86
rect 78 79 79 81
rect 81 79 82 81
rect 78 73 82 79
rect 86 81 90 86
rect 86 79 87 81
rect 89 79 90 81
rect 86 77 90 79
rect 78 71 79 73
rect 81 71 82 73
rect 6 41 10 55
rect 6 39 7 41
rect 9 39 10 41
rect 6 33 10 39
rect 78 66 82 71
rect 78 64 79 66
rect 81 64 82 66
rect 78 62 82 64
rect 22 41 26 55
rect 22 39 23 41
rect 25 39 26 41
rect 22 33 26 39
rect 46 50 50 52
rect 46 48 47 50
rect 49 48 50 50
rect 46 32 50 48
rect 46 30 47 32
rect 49 30 50 32
rect 14 14 18 16
rect 14 12 15 14
rect 17 12 18 14
rect 14 9 18 12
rect 46 17 50 30
rect 54 42 74 47
rect 54 41 58 42
rect 54 39 55 41
rect 57 39 58 41
rect 54 25 58 39
rect 70 41 74 42
rect 70 39 71 41
rect 73 39 74 41
rect 70 37 74 39
rect 78 25 82 27
rect 78 23 79 25
rect 81 23 82 25
rect 78 17 82 23
rect 78 15 79 17
rect 81 15 82 17
rect 78 9 82 15
rect 14 7 15 9
rect 17 7 18 9
rect 14 6 18 7
rect 14 4 15 6
rect 17 4 18 6
rect 14 2 18 4
rect 78 7 79 9
rect 81 7 82 9
rect 78 2 82 7
rect -2 1 98 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 73 -1 87 1
rect 89 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< alu2 >>
rect -2 89 98 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 71 89
rect 73 87 87 89
rect 89 87 98 89
rect -2 81 98 87
rect -2 79 15 81
rect 17 79 79 81
rect 81 79 98 81
rect -2 76 98 79
rect -2 9 98 12
rect -2 7 15 9
rect 17 7 79 9
rect 81 7 98 9
rect -2 1 98 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 71 1
rect 73 -1 87 1
rect 89 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 71 3
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 57 -3 71 -1
rect 89 1 96 3
rect 89 -1 91 1
rect 93 -1 96 1
rect 89 -3 96 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 71 91
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 57 85 71 87
rect 89 89 96 91
rect 89 87 91 89
rect 93 87 96 89
rect 89 85 96 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polyct0 >>
rect 39 39 41 41
<< polyct1 >>
rect 87 79 89 81
rect 7 39 9 41
rect 23 39 25 41
rect 55 39 57 41
rect 71 39 73 41
<< ndifct0 >>
rect 4 25 6 27
rect 4 18 6 20
rect 26 27 28 29
rect 36 26 38 28
rect 36 19 38 21
rect 58 16 60 18
rect 68 30 70 32
rect 68 23 70 25
<< ndifct1 >>
rect 47 30 49 32
rect 79 23 81 25
rect 79 15 81 17
rect 15 12 17 14
rect 15 4 17 6
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
rect 67 87 69 89
rect 91 87 93 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 26 59 28 61
rect 36 70 38 72
rect 58 70 60 72
rect 58 63 60 65
rect 68 63 70 65
rect 68 56 70 58
<< pdifct1 >>
rect 15 82 17 84
rect 15 74 17 76
rect 47 48 49 50
rect 79 71 81 73
rect 79 64 81 66
<< alu0 >>
rect 22 72 40 73
rect 22 70 36 72
rect 38 70 40 72
rect 22 69 40 70
rect 56 72 62 73
rect 56 70 58 72
rect 60 70 62 72
rect 2 68 26 69
rect 2 66 4 68
rect 6 66 26 68
rect 56 66 62 70
rect 2 65 26 66
rect 30 65 62 66
rect 2 61 8 65
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 14 29 18 65
rect 30 63 58 65
rect 60 63 62 65
rect 30 62 62 63
rect 67 65 71 67
rect 67 63 68 65
rect 70 63 71 65
rect 24 61 34 62
rect 24 59 26 61
rect 28 59 34 61
rect 67 59 71 63
rect 24 58 34 59
rect 30 30 34 58
rect 38 58 82 59
rect 38 56 68 58
rect 70 56 82 58
rect 38 55 82 56
rect 38 41 42 55
rect 38 39 39 41
rect 41 39 42 41
rect 38 37 42 39
rect 3 27 18 29
rect 3 25 4 27
rect 6 25 18 27
rect 24 29 39 30
rect 24 27 26 29
rect 28 28 39 29
rect 28 27 36 28
rect 24 26 36 27
rect 38 26 39 28
rect 3 20 7 25
rect 3 18 4 20
rect 6 18 7 20
rect 14 23 18 25
rect 14 19 26 23
rect 3 16 7 18
rect 22 13 26 19
rect 35 21 39 26
rect 35 19 36 21
rect 38 19 39 21
rect 35 17 39 19
rect 78 34 82 55
rect 67 32 82 34
rect 67 30 68 32
rect 70 30 82 32
rect 67 25 71 30
rect 67 23 68 25
rect 70 23 71 25
rect 67 21 71 23
rect 57 18 61 20
rect 57 16 58 18
rect 60 16 61 18
rect 57 13 61 16
rect 22 9 61 13
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 71 87 73 89
rect 87 87 89 89
rect 15 79 17 81
rect 79 79 81 81
rect 15 7 17 9
rect 79 7 81 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
rect 71 -1 73 1
rect 87 -1 89 1
<< labels >>
rlabel alu1 8 44 8 44 6 a1
rlabel alu1 24 44 24 44 6 a0
rlabel alu1 48 32 48 32 6 z
rlabel alu1 56 36 56 36 6 s
rlabel alu1 64 44 64 44 6 s
rlabel alu1 72 44 72 44 6 s
rlabel alu2 48 6 48 6 6 vss
rlabel alu2 48 82 48 82 6 vdd
<< end >>
