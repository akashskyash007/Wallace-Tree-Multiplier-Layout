magic
tech scmos
timestamp 1199203146
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 13 64 15 69
rect 21 64 23 69
rect 31 64 33 69
rect 39 64 41 69
rect 13 43 15 48
rect 21 43 23 48
rect 9 41 15 43
rect 9 39 11 41
rect 13 39 15 41
rect 9 37 15 39
rect 20 41 26 43
rect 20 39 22 41
rect 24 39 26 41
rect 20 37 26 39
rect 9 19 11 37
rect 20 26 22 37
rect 31 35 33 48
rect 39 45 41 48
rect 39 43 46 45
rect 39 41 42 43
rect 44 41 46 43
rect 39 39 46 41
rect 30 33 36 35
rect 30 31 32 33
rect 34 31 36 33
rect 30 29 36 31
rect 30 26 32 29
rect 20 14 22 19
rect 30 14 32 19
rect 41 18 43 39
rect 9 7 11 12
rect 41 6 43 11
<< ndif >>
rect 13 24 20 26
rect 13 22 15 24
rect 17 22 20 24
rect 13 19 20 22
rect 22 23 30 26
rect 22 21 25 23
rect 27 21 30 23
rect 22 19 30 21
rect 32 19 39 26
rect 2 16 9 19
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 12 17 19
rect 34 18 39 19
rect 34 11 41 18
rect 43 16 50 18
rect 43 14 46 16
rect 48 14 50 16
rect 43 11 50 14
rect 34 9 39 11
rect 33 7 39 9
rect 33 5 35 7
rect 37 5 39 7
rect 33 3 39 5
<< pdif >>
rect 4 67 11 69
rect 4 65 7 67
rect 9 65 11 67
rect 4 64 11 65
rect 4 48 13 64
rect 15 48 21 64
rect 23 58 31 64
rect 23 56 26 58
rect 28 56 31 58
rect 23 48 31 56
rect 33 48 39 64
rect 41 62 48 64
rect 41 60 44 62
rect 46 60 48 62
rect 41 48 48 60
<< alu1 >>
rect -2 67 58 72
rect -2 65 7 67
rect 9 65 58 67
rect -2 64 58 65
rect 2 58 30 59
rect 2 56 26 58
rect 28 56 30 58
rect 2 55 30 56
rect 2 53 14 55
rect 2 26 6 53
rect 10 41 14 43
rect 10 39 11 41
rect 13 39 14 41
rect 10 34 14 39
rect 18 42 22 51
rect 34 50 38 59
rect 34 46 47 50
rect 41 43 47 46
rect 18 41 31 42
rect 18 39 22 41
rect 24 39 31 41
rect 18 38 31 39
rect 41 41 42 43
rect 44 41 47 43
rect 41 38 47 41
rect 10 30 23 34
rect 30 33 39 34
rect 30 31 32 33
rect 34 31 39 33
rect 30 30 39 31
rect 33 27 39 30
rect 2 24 19 26
rect 2 22 15 24
rect 17 22 19 24
rect 2 21 19 22
rect 33 21 46 27
rect -2 7 58 8
rect -2 5 24 7
rect 26 5 35 7
rect 37 5 58 7
rect -2 0 58 5
<< ptie >>
rect 21 7 29 9
rect 21 5 24 7
rect 26 5 29 7
rect 21 3 29 5
<< nmos >>
rect 20 19 22 26
rect 30 19 32 26
rect 9 12 11 19
rect 41 11 43 18
<< pmos >>
rect 13 48 15 64
rect 21 48 23 64
rect 31 48 33 64
rect 39 48 41 64
<< polyct1 >>
rect 11 39 13 41
rect 22 39 24 41
rect 42 41 44 43
rect 32 31 34 33
<< ndifct0 >>
rect 25 21 27 23
rect 4 14 6 16
rect 46 14 48 16
<< ndifct1 >>
rect 15 22 17 24
rect 35 5 37 7
<< ptiect1 >>
rect 24 5 26 7
<< pdifct0 >>
rect 44 60 46 62
<< pdifct1 >>
rect 7 65 9 67
rect 26 56 28 58
<< alu0 >>
rect 43 62 47 64
rect 43 60 44 62
rect 46 60 47 62
rect 43 58 47 60
rect 24 23 28 25
rect 24 21 25 23
rect 27 21 28 23
rect 24 17 28 21
rect 2 16 50 17
rect 2 14 4 16
rect 6 14 46 16
rect 48 14 50 16
rect 2 13 50 14
<< labels >>
rlabel alu0 26 19 26 19 6 n3
rlabel alu0 26 15 26 15 6 n3
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 20 32 20 32 6 b1
rlabel polyct1 12 40 12 40 6 b1
rlabel alu1 20 48 20 48 6 b2
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 28 40 28 40 6 b2
rlabel alu1 36 56 36 56 6 a1
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 24 44 24 6 a2
rlabel alu1 44 44 44 44 6 a1
<< end >>
