magic
tech scmos
timestamp 1199203662
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 20 65 22 70
rect 30 65 32 70
rect 40 65 42 70
rect 50 65 52 70
rect 2 56 8 58
rect 2 54 4 56
rect 6 54 8 56
rect 2 52 11 54
rect 9 49 11 52
rect 61 51 63 56
rect 9 35 11 38
rect 20 35 22 38
rect 30 35 32 38
rect 9 33 22 35
rect 26 33 32 35
rect 9 24 11 33
rect 26 31 28 33
rect 30 31 32 33
rect 26 29 32 31
rect 40 35 42 38
rect 50 35 52 38
rect 61 35 63 40
rect 40 33 46 35
rect 40 31 42 33
rect 44 31 46 33
rect 40 29 46 31
rect 50 33 70 35
rect 19 27 28 29
rect 19 24 21 27
rect 40 26 42 29
rect 50 26 52 33
rect 61 31 66 33
rect 68 31 70 33
rect 61 29 70 31
rect 61 26 63 29
rect 9 4 11 18
rect 29 19 31 23
rect 19 8 21 12
rect 61 15 63 20
rect 40 9 42 14
rect 50 9 52 14
rect 29 4 31 7
rect 9 2 31 4
<< ndif >>
rect 33 24 40 26
rect 2 22 9 24
rect 2 20 4 22
rect 6 20 9 22
rect 2 18 9 20
rect 11 22 19 24
rect 11 20 14 22
rect 16 20 19 22
rect 11 18 19 20
rect 13 12 19 18
rect 21 19 26 24
rect 33 22 35 24
rect 37 22 40 24
rect 33 19 40 22
rect 21 16 29 19
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 24 7 29 12
rect 31 14 40 19
rect 42 18 50 26
rect 42 16 45 18
rect 47 16 50 18
rect 42 14 50 16
rect 52 20 61 26
rect 63 24 70 26
rect 63 22 66 24
rect 68 22 70 24
rect 63 20 70 22
rect 52 18 59 20
rect 52 16 55 18
rect 57 16 59 18
rect 52 14 59 16
rect 31 7 36 14
<< pdif >>
rect 13 61 20 65
rect 13 59 15 61
rect 17 59 20 61
rect 13 49 20 59
rect 4 44 9 49
rect 2 42 9 44
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 38 20 49
rect 22 58 30 65
rect 22 56 25 58
rect 27 56 30 58
rect 22 38 30 56
rect 32 49 40 65
rect 32 47 35 49
rect 37 47 40 49
rect 32 42 40 47
rect 32 40 35 42
rect 37 40 40 42
rect 32 38 40 40
rect 42 58 50 65
rect 42 56 45 58
rect 47 56 50 58
rect 42 38 50 56
rect 52 57 59 65
rect 52 55 55 57
rect 57 55 59 57
rect 52 51 59 55
rect 52 40 61 51
rect 63 49 70 51
rect 63 47 66 49
rect 68 47 70 49
rect 63 45 70 47
rect 63 40 68 45
rect 52 38 59 40
<< alu1 >>
rect -2 67 74 72
rect -2 65 5 67
rect 7 65 65 67
rect 67 65 74 67
rect -2 64 74 65
rect 2 56 7 59
rect 2 54 4 56
rect 6 54 7 56
rect 2 50 14 54
rect 10 45 14 50
rect 26 49 38 51
rect 26 47 35 49
rect 37 47 38 49
rect 26 45 38 47
rect 34 42 38 45
rect 34 40 35 42
rect 37 40 38 42
rect 34 24 38 40
rect 57 38 70 42
rect 65 33 70 38
rect 65 31 66 33
rect 68 31 70 33
rect 65 29 70 31
rect 34 22 35 24
rect 37 22 38 24
rect 34 20 38 22
rect -2 7 74 8
rect -2 5 65 7
rect 67 5 74 7
rect -2 0 74 5
<< ptie >>
rect 63 7 69 13
rect 63 5 65 7
rect 67 5 69 7
rect 63 3 69 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 63 67 69 69
rect 63 65 65 67
rect 67 65 69 67
rect 3 63 9 65
rect 63 59 69 65
<< nmos >>
rect 9 18 11 24
rect 19 12 21 24
rect 29 7 31 19
rect 40 14 42 26
rect 50 14 52 26
rect 61 20 63 26
<< pmos >>
rect 9 38 11 49
rect 20 38 22 65
rect 30 38 32 65
rect 40 38 42 65
rect 50 38 52 65
rect 61 40 63 51
<< polyct0 >>
rect 28 31 30 33
rect 42 31 44 33
<< polyct1 >>
rect 4 54 6 56
rect 66 31 68 33
<< ndifct0 >>
rect 4 20 6 22
rect 14 20 16 22
rect 24 14 26 16
rect 45 16 47 18
rect 66 22 68 24
rect 55 16 57 18
<< ndifct1 >>
rect 35 22 37 24
<< ntiect1 >>
rect 5 65 7 67
rect 65 65 67 67
<< ptiect1 >>
rect 65 5 67 7
<< pdifct0 >>
rect 15 59 17 61
rect 4 40 6 42
rect 25 56 27 58
rect 45 56 47 58
rect 55 55 57 57
rect 66 47 68 49
<< pdifct1 >>
rect 35 47 37 49
rect 35 40 37 42
<< alu0 >>
rect 13 61 19 64
rect 13 59 15 61
rect 17 59 19 61
rect 13 58 19 59
rect 23 58 49 59
rect 23 56 25 58
rect 27 56 45 58
rect 47 56 49 58
rect 23 55 49 56
rect 53 57 59 64
rect 53 55 55 57
rect 57 55 59 57
rect 53 54 59 55
rect 3 42 7 44
rect 3 40 4 42
rect 6 40 7 42
rect 3 33 7 40
rect 27 33 31 35
rect 3 31 28 33
rect 30 31 31 33
rect 3 29 31 31
rect 3 22 7 29
rect 50 49 70 50
rect 50 47 66 49
rect 68 47 70 49
rect 50 46 70 47
rect 50 35 54 46
rect 41 33 54 35
rect 41 31 42 33
rect 44 31 54 33
rect 41 29 54 31
rect 3 20 4 22
rect 6 20 7 22
rect 3 18 7 20
rect 13 22 17 24
rect 13 20 14 22
rect 16 20 17 22
rect 50 26 54 29
rect 50 24 70 26
rect 50 22 66 24
rect 68 22 70 24
rect 64 21 70 22
rect 13 8 17 20
rect 43 18 49 19
rect 43 17 45 18
rect 22 16 45 17
rect 47 16 49 18
rect 22 14 24 16
rect 26 14 49 16
rect 22 13 49 14
rect 53 18 59 19
rect 53 16 55 18
rect 57 16 59 18
rect 53 8 59 16
<< labels >>
rlabel alu0 17 31 17 31 6 bn
rlabel polyct0 29 32 29 32 6 bn
rlabel alu0 35 15 35 15 6 n2
rlabel alu0 46 16 46 16 6 n2
rlabel alu0 36 57 36 57 6 n1
rlabel alu0 47 32 47 32 6 an
rlabel ndifct0 67 23 67 23 6 an
rlabel alu0 60 48 60 48 6 an
rlabel alu1 12 48 12 48 6 b
rlabel alu1 4 56 4 56 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 36 36 36 36 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 68 32 68 32 6 a
rlabel alu1 60 40 60 40 6 a
<< end >>
