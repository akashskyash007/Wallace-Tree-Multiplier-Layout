magic
tech scmos
timestamp 1199202358
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 69 11 73
rect 19 69 21 73
rect 29 69 31 73
rect 39 61 41 65
rect 9 39 11 43
rect 19 39 21 43
rect 29 39 31 43
rect 39 39 41 43
rect 9 37 41 39
rect 14 30 16 37
rect 24 35 29 37
rect 31 35 37 37
rect 39 35 41 37
rect 24 33 41 35
rect 24 30 26 33
rect 14 13 16 18
rect 24 13 26 18
<< ndif >>
rect 6 22 14 30
rect 6 20 9 22
rect 11 20 14 22
rect 6 18 14 20
rect 16 28 24 30
rect 16 26 19 28
rect 21 26 24 28
rect 16 18 24 26
rect 26 22 34 30
rect 26 20 29 22
rect 31 20 34 22
rect 26 18 34 20
<< pdif >>
rect 2 67 9 69
rect 2 65 4 67
rect 6 65 9 67
rect 2 60 9 65
rect 2 58 4 60
rect 6 58 9 60
rect 2 43 9 58
rect 11 54 19 69
rect 11 52 14 54
rect 16 52 19 54
rect 11 47 19 52
rect 11 45 14 47
rect 16 45 19 47
rect 11 43 19 45
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 43 29 58
rect 31 61 36 69
rect 31 54 39 61
rect 31 52 34 54
rect 36 52 39 54
rect 31 47 39 52
rect 31 45 34 47
rect 36 45 39 47
rect 31 43 39 45
rect 41 59 48 61
rect 41 57 44 59
rect 46 57 48 59
rect 41 52 48 57
rect 41 50 44 52
rect 46 50 48 52
rect 41 43 48 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 33 54 39 56
rect 33 52 34 54
rect 36 52 39 54
rect 33 47 39 52
rect 33 46 34 47
rect 9 45 14 46
rect 16 45 34 46
rect 36 45 39 47
rect 9 42 39 45
rect 18 28 22 42
rect 27 37 47 38
rect 27 35 29 37
rect 31 35 37 37
rect 39 35 47 37
rect 27 34 47 35
rect 18 26 19 28
rect 21 26 22 28
rect 41 26 47 34
rect 18 24 22 26
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 14 18 16 30
rect 24 18 26 30
<< pmos >>
rect 9 43 11 69
rect 19 43 21 69
rect 29 43 31 69
rect 39 43 41 61
<< polyct1 >>
rect 29 35 31 37
rect 37 35 39 37
<< ndifct0 >>
rect 9 20 11 22
rect 29 20 31 22
<< ndifct1 >>
rect 19 26 21 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 65 6 67
rect 4 58 6 60
rect 14 52 16 54
rect 14 46 16 47
rect 24 65 26 67
rect 24 58 26 60
rect 44 57 46 59
rect 44 50 46 52
<< pdifct1 >>
rect 14 45 16 46
rect 34 52 36 54
rect 34 45 36 47
<< alu0 >>
rect 3 67 7 68
rect 3 65 4 67
rect 6 65 7 67
rect 3 60 7 65
rect 3 58 4 60
rect 6 58 7 60
rect 3 56 7 58
rect 23 67 27 68
rect 23 65 24 67
rect 26 65 27 67
rect 23 60 27 65
rect 23 58 24 60
rect 26 58 27 60
rect 23 56 27 58
rect 42 59 48 68
rect 42 57 44 59
rect 46 57 48 59
rect 13 54 17 56
rect 13 52 14 54
rect 16 52 17 54
rect 13 47 17 52
rect 13 46 14 47
rect 16 46 17 47
rect 42 52 48 57
rect 42 50 44 52
rect 46 50 48 52
rect 42 49 48 50
rect 8 22 12 24
rect 8 20 9 22
rect 11 20 12 22
rect 8 12 12 20
rect 28 22 32 24
rect 28 20 29 22
rect 31 20 32 22
rect 28 12 32 20
<< labels >>
rlabel alu1 20 36 20 36 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 36 36 36 6 a
rlabel alu1 28 44 28 44 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 a
<< end >>
