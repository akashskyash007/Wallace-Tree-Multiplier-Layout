magic
tech scmos
timestamp 1199201837
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 29 62 31 67
rect 9 54 11 59
rect 19 54 21 59
rect 29 43 31 46
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 9 35 11 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 31 21 38
rect 29 37 35 39
rect 19 29 25 31
rect 12 21 14 29
rect 19 27 21 29
rect 23 27 25 29
rect 19 25 25 27
rect 22 22 24 25
rect 29 22 31 37
rect 12 11 14 15
rect 22 11 24 15
rect 29 11 31 15
<< ndif >>
rect 17 21 22 22
rect 3 15 12 21
rect 14 19 22 21
rect 14 17 17 19
rect 19 17 22 19
rect 14 15 22 17
rect 24 15 29 22
rect 31 15 38 22
rect 3 7 10 15
rect 33 9 38 15
rect 3 5 6 7
rect 8 5 10 7
rect 3 3 10 5
rect 32 7 38 9
rect 32 5 34 7
rect 36 5 38 7
rect 32 3 38 5
<< pdif >>
rect 21 67 27 69
rect 21 65 23 67
rect 25 65 27 67
rect 21 62 27 65
rect 21 61 29 62
rect 23 54 29 61
rect 4 51 9 54
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 52 19 54
rect 11 50 14 52
rect 16 50 19 52
rect 11 38 19 50
rect 21 46 29 54
rect 31 59 36 62
rect 31 57 38 59
rect 31 55 34 57
rect 36 55 38 57
rect 31 50 38 55
rect 31 48 34 50
rect 36 48 38 50
rect 31 46 38 48
rect 21 38 27 46
<< alu1 >>
rect -2 67 42 72
rect -2 65 5 67
rect 7 65 13 67
rect 15 65 23 67
rect 25 65 42 67
rect -2 64 42 65
rect 2 49 6 51
rect 2 47 4 49
rect 2 42 6 47
rect 2 40 4 42
rect 2 19 6 40
rect 26 43 30 51
rect 10 37 22 43
rect 26 41 38 43
rect 26 39 31 41
rect 33 39 38 41
rect 26 37 38 39
rect 10 33 14 37
rect 10 31 11 33
rect 13 31 14 33
rect 10 29 14 31
rect 19 29 25 30
rect 19 27 21 29
rect 23 27 30 29
rect 19 25 30 27
rect 26 19 30 25
rect 2 17 17 19
rect 19 17 22 19
rect 2 13 22 17
rect 26 13 38 19
rect -2 7 42 8
rect -2 5 6 7
rect 8 5 16 7
rect 18 5 24 7
rect 26 5 34 7
rect 36 5 42 7
rect -2 0 42 5
<< ptie >>
rect 14 7 28 9
rect 14 5 16 7
rect 18 5 24 7
rect 26 5 28 7
rect 14 3 28 5
<< ntie >>
rect 3 67 17 69
rect 3 65 5 67
rect 7 65 13 67
rect 15 65 17 67
rect 3 63 17 65
<< nmos >>
rect 12 15 14 21
rect 22 15 24 22
rect 29 15 31 22
<< pmos >>
rect 9 38 11 54
rect 19 38 21 54
rect 29 46 31 62
<< polyct1 >>
rect 31 39 33 41
rect 11 31 13 33
rect 21 27 23 29
<< ndifct1 >>
rect 17 17 19 19
rect 6 5 8 7
rect 34 5 36 7
<< ntiect1 >>
rect 5 65 7 67
rect 13 65 15 67
<< ptiect1 >>
rect 16 5 18 7
rect 24 5 26 7
<< pdifct0 >>
rect 14 50 16 52
rect 34 55 36 57
rect 34 48 36 50
<< pdifct1 >>
rect 23 65 25 67
rect 4 47 6 49
rect 4 40 6 42
<< alu0 >>
rect 13 57 37 59
rect 13 55 34 57
rect 36 55 37 57
rect 13 52 17 55
rect 6 38 7 51
rect 13 50 14 52
rect 16 50 17 52
rect 13 48 17 50
rect 33 50 37 55
rect 33 48 34 50
rect 36 48 37 50
rect 33 46 37 48
rect 16 19 20 21
<< labels >>
rlabel alu0 15 53 15 53 6 n1
rlabel alu0 35 52 35 52 6 n1
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 12 36 12 36 6 b
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 28 20 28 20 6 a2
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 40 20 40 6 b
rlabel alu1 28 44 28 44 6 a1
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 36 16 36 16 6 a2
rlabel alu1 36 40 36 40 6 a1
<< end >>
