magic
tech scmos
timestamp 1199202869
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 10 70 12 74
rect 17 70 19 74
rect 27 70 29 74
rect 34 70 36 74
rect 44 66 46 71
rect 10 39 12 42
rect 17 39 19 42
rect 27 39 29 42
rect 34 39 36 42
rect 4 37 13 39
rect 4 35 6 37
rect 8 35 13 37
rect 4 33 13 35
rect 17 37 29 39
rect 33 37 39 39
rect 17 35 19 37
rect 21 35 23 37
rect 17 33 23 35
rect 33 35 35 37
rect 37 35 39 37
rect 33 33 39 35
rect 11 30 13 33
rect 21 30 23 33
rect 44 31 46 42
rect 44 29 50 31
rect 44 27 46 29
rect 48 27 50 29
rect 33 25 50 27
rect 33 22 35 25
rect 11 10 13 15
rect 21 10 23 15
rect 33 6 35 10
<< ndif >>
rect 2 15 11 30
rect 13 28 21 30
rect 13 26 16 28
rect 18 26 21 28
rect 13 15 21 26
rect 23 22 31 30
rect 23 15 33 22
rect 2 11 9 15
rect 2 9 5 11
rect 7 9 9 11
rect 25 11 33 15
rect 2 7 9 9
rect 25 9 27 11
rect 29 10 33 11
rect 35 20 42 22
rect 35 18 38 20
rect 40 18 42 20
rect 35 16 42 18
rect 35 10 40 16
rect 29 9 31 10
rect 25 7 31 9
<< pdif >>
rect 2 68 10 70
rect 2 66 5 68
rect 7 66 10 68
rect 2 61 10 66
rect 2 59 5 61
rect 7 59 10 61
rect 2 42 10 59
rect 12 42 17 70
rect 19 60 27 70
rect 19 58 22 60
rect 24 58 27 60
rect 19 53 27 58
rect 19 51 22 53
rect 24 51 27 53
rect 19 42 27 51
rect 29 42 34 70
rect 36 66 42 70
rect 36 64 44 66
rect 36 62 39 64
rect 41 62 44 64
rect 36 56 44 62
rect 36 54 39 56
rect 41 54 44 56
rect 36 42 44 54
rect 46 55 51 66
rect 46 53 53 55
rect 46 51 49 53
rect 51 51 53 53
rect 46 46 53 51
rect 46 44 49 46
rect 51 44 53 46
rect 46 42 53 44
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 17 53 30 55
rect 17 51 22 53
rect 24 51 30 53
rect 17 50 30 51
rect 9 42 22 46
rect 18 37 22 42
rect 18 35 19 37
rect 21 35 22 37
rect 18 33 22 35
rect 26 29 30 50
rect 14 28 30 29
rect 14 26 16 28
rect 18 26 30 28
rect 14 25 30 26
rect 42 29 54 31
rect 42 27 46 29
rect 48 27 54 29
rect 42 25 54 27
rect 50 17 54 25
rect -2 11 58 12
rect -2 9 5 11
rect 7 9 27 11
rect 29 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 11 15 13 30
rect 21 15 23 30
rect 33 10 35 22
<< pmos >>
rect 10 42 12 70
rect 17 42 19 70
rect 27 42 29 70
rect 34 42 36 70
rect 44 42 46 66
<< polyct0 >>
rect 6 35 8 37
rect 35 35 37 37
<< polyct1 >>
rect 19 35 21 37
rect 46 27 48 29
<< ndifct0 >>
rect 38 18 40 20
<< ndifct1 >>
rect 16 26 18 28
rect 5 9 7 11
rect 27 9 29 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 5 66 7 68
rect 5 59 7 61
rect 22 58 24 60
rect 39 62 41 64
rect 39 54 41 56
rect 49 51 51 53
rect 49 44 51 46
<< pdifct1 >>
rect 22 51 24 53
<< alu0 >>
rect 3 66 5 68
rect 7 66 9 68
rect 3 61 9 66
rect 38 64 42 68
rect 38 62 39 64
rect 41 62 42 64
rect 3 59 5 61
rect 7 59 9 61
rect 3 58 9 59
rect 21 60 25 62
rect 21 58 22 60
rect 24 58 25 60
rect 21 55 25 58
rect 38 56 42 62
rect 38 54 39 56
rect 41 54 42 56
rect 38 52 42 54
rect 48 53 52 55
rect 5 37 9 39
rect 5 35 6 37
rect 8 35 9 37
rect 5 21 9 35
rect 48 51 49 53
rect 51 51 52 53
rect 48 46 52 51
rect 48 44 49 46
rect 51 44 52 46
rect 48 39 52 44
rect 34 37 52 39
rect 34 35 35 37
rect 37 35 52 37
rect 34 21 38 35
rect 5 20 42 21
rect 5 18 38 20
rect 40 18 42 20
rect 5 17 42 18
<< labels >>
rlabel alu0 7 28 7 28 6 an
rlabel alu0 36 28 36 28 6 an
rlabel alu0 23 19 23 19 6 an
rlabel pdifct0 50 45 50 45 6 an
rlabel alu1 12 44 12 44 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 40 28 40 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a
rlabel alu1 52 24 52 24 6 a
<< end >>
