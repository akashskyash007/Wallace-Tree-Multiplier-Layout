magic
tech scmos
timestamp 1199201665
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 39 58 41 63
rect 49 58 51 63
rect 59 58 61 63
rect 69 58 71 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 9 37 32 39
rect 20 35 27 37
rect 29 35 32 37
rect 20 33 32 35
rect 39 37 45 39
rect 39 35 41 37
rect 43 35 45 37
rect 39 33 45 35
rect 49 37 61 39
rect 69 37 71 42
rect 49 35 57 37
rect 59 35 61 37
rect 49 33 61 35
rect 20 30 22 33
rect 30 30 32 33
rect 42 30 44 33
rect 49 30 51 33
rect 59 30 61 33
rect 66 35 71 37
rect 66 30 68 35
rect 20 6 22 10
rect 30 6 32 10
rect 42 8 44 17
rect 49 12 51 17
rect 59 12 61 17
rect 66 8 68 17
rect 42 6 68 8
<< ndif >>
rect 13 21 20 30
rect 13 19 15 21
rect 17 19 20 21
rect 13 14 20 19
rect 13 12 15 14
rect 17 12 20 14
rect 13 10 20 12
rect 22 28 30 30
rect 22 26 25 28
rect 27 26 30 28
rect 22 21 30 26
rect 22 19 25 21
rect 27 19 30 21
rect 22 10 30 19
rect 32 17 42 30
rect 44 17 49 30
rect 51 21 59 30
rect 51 19 54 21
rect 56 19 59 21
rect 51 17 59 19
rect 61 17 66 30
rect 68 28 75 30
rect 68 26 71 28
rect 73 26 75 28
rect 68 21 75 26
rect 68 19 71 21
rect 73 19 75 21
rect 68 17 75 19
rect 32 14 39 17
rect 32 12 35 14
rect 37 12 39 14
rect 32 10 39 12
<< pdif >>
rect 4 55 9 69
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 67 19 69
rect 11 65 14 67
rect 16 65 19 67
rect 11 60 19 65
rect 11 58 14 60
rect 16 58 19 60
rect 11 42 19 58
rect 21 53 29 69
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 58 37 69
rect 31 56 39 58
rect 31 54 34 56
rect 36 54 39 56
rect 31 42 39 54
rect 41 53 49 58
rect 41 51 44 53
rect 46 51 49 53
rect 41 46 49 51
rect 41 44 44 46
rect 46 44 49 46
rect 41 42 49 44
rect 51 56 59 58
rect 51 54 54 56
rect 56 54 59 56
rect 51 42 59 54
rect 61 54 69 58
rect 61 52 64 54
rect 66 52 69 54
rect 61 47 69 52
rect 61 45 64 47
rect 66 45 69 47
rect 61 42 69 45
rect 71 56 78 58
rect 71 54 74 56
rect 76 54 78 56
rect 71 42 78 54
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 23 53 27 55
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 2 44 4 46
rect 6 44 24 46
rect 26 44 27 46
rect 2 42 27 44
rect 9 30 14 42
rect 74 38 78 47
rect 39 37 47 38
rect 39 35 41 37
rect 43 35 47 37
rect 39 34 47 35
rect 55 37 78 38
rect 55 35 57 37
rect 59 35 78 37
rect 55 34 78 35
rect 9 28 28 30
rect 9 26 25 28
rect 27 26 28 28
rect 24 21 28 26
rect 24 19 25 21
rect 27 19 28 21
rect 24 17 28 19
rect 41 30 47 34
rect 41 26 55 30
rect -2 1 82 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 20 10 22 30
rect 30 10 32 30
rect 42 17 44 30
rect 49 17 51 30
rect 59 17 61 30
rect 66 17 68 30
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
rect 39 42 41 58
rect 49 42 51 58
rect 59 42 61 58
rect 69 42 71 58
<< polyct0 >>
rect 27 35 29 37
<< polyct1 >>
rect 41 35 43 37
rect 57 35 59 37
<< ndifct0 >>
rect 15 19 17 21
rect 15 12 17 14
rect 54 19 56 21
rect 71 26 73 28
rect 71 19 73 21
rect 35 12 37 14
<< ndifct1 >>
rect 25 26 27 28
rect 25 19 27 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 14 65 16 67
rect 14 58 16 60
rect 34 54 36 56
rect 44 51 46 53
rect 44 44 46 46
rect 54 54 56 56
rect 64 52 66 54
rect 64 45 66 47
rect 74 54 76 56
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 51 26 53
rect 24 44 26 46
<< alu0 >>
rect 13 67 17 68
rect 13 65 14 67
rect 16 65 17 67
rect 13 60 17 65
rect 13 58 14 60
rect 16 58 17 60
rect 13 56 17 58
rect 33 56 37 68
rect 33 54 34 56
rect 36 54 37 56
rect 53 56 57 68
rect 73 56 77 68
rect 33 52 37 54
rect 43 53 47 55
rect 43 51 44 53
rect 46 51 47 53
rect 53 54 54 56
rect 56 54 57 56
rect 53 52 57 54
rect 63 54 67 56
rect 63 52 64 54
rect 66 52 67 54
rect 73 54 74 56
rect 76 54 77 56
rect 73 52 77 54
rect 43 47 47 51
rect 63 47 67 52
rect 31 46 64 47
rect 31 44 44 46
rect 46 45 64 46
rect 66 45 67 47
rect 46 44 67 45
rect 31 43 67 44
rect 31 38 35 43
rect 25 37 35 38
rect 25 35 27 37
rect 29 35 35 37
rect 25 34 35 35
rect 13 21 19 22
rect 13 19 15 21
rect 17 19 19 21
rect 13 14 19 19
rect 31 22 35 34
rect 70 28 74 30
rect 70 26 71 28
rect 73 26 74 28
rect 31 21 58 22
rect 31 19 54 21
rect 56 19 58 21
rect 31 18 58 19
rect 70 21 74 26
rect 70 19 71 21
rect 73 19 74 21
rect 13 12 15 14
rect 17 12 19 14
rect 33 14 39 15
rect 33 12 35 14
rect 37 12 39 14
rect 70 12 74 19
<< labels >>
rlabel alu0 30 36 30 36 6 zn
rlabel alu0 44 20 44 20 6 zn
rlabel alu0 45 49 45 49 6 zn
rlabel alu0 49 45 49 45 6 zn
rlabel alu0 65 49 65 49 6 zn
rlabel alu1 12 36 12 36 6 z
rlabel alu1 4 52 4 52 6 z
rlabel alu1 20 28 20 28 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 44 32 44 32 6 a
rlabel alu1 52 28 52 28 6 a
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 36 60 36 6 b
rlabel alu1 68 36 68 36 6 b
rlabel alu1 76 44 76 44 6 b
<< end >>
