magic
tech scmos
timestamp 1199201810
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 12 32 14 43
rect 19 40 21 43
rect 29 40 31 43
rect 39 40 41 43
rect 19 38 25 40
rect 19 36 21 38
rect 23 36 25 38
rect 19 34 25 36
rect 29 38 35 40
rect 29 36 31 38
rect 33 36 35 38
rect 29 34 35 36
rect 39 38 47 40
rect 39 36 43 38
rect 45 36 47 38
rect 39 34 47 36
rect 9 30 15 32
rect 9 28 11 30
rect 13 28 15 30
rect 9 26 15 28
rect 10 23 12 26
rect 20 23 22 34
rect 32 26 34 34
rect 39 26 41 34
rect 10 12 12 17
rect 20 12 22 17
rect 32 12 34 17
rect 39 12 41 17
<< ndif >>
rect 24 23 32 26
rect 2 17 10 23
rect 12 21 20 23
rect 12 19 15 21
rect 17 19 20 21
rect 12 17 20 19
rect 22 17 32 23
rect 34 17 39 26
rect 41 23 46 26
rect 41 21 48 23
rect 41 19 44 21
rect 46 19 48 21
rect 41 17 48 19
rect 2 11 8 17
rect 2 9 4 11
rect 6 9 8 11
rect 2 7 8 9
rect 24 11 30 17
rect 24 9 26 11
rect 28 9 30 11
rect 24 7 30 9
<< pdif >>
rect 7 64 12 70
rect 5 62 12 64
rect 5 60 7 62
rect 9 60 12 62
rect 5 54 12 60
rect 5 52 7 54
rect 9 52 12 54
rect 5 50 12 52
rect 7 43 12 50
rect 14 43 19 70
rect 21 61 29 70
rect 21 59 24 61
rect 26 59 29 61
rect 21 43 29 59
rect 31 68 39 70
rect 31 66 34 68
rect 36 66 39 68
rect 31 43 39 66
rect 41 63 46 70
rect 41 61 48 63
rect 41 59 44 61
rect 46 59 48 61
rect 41 57 48 59
rect 41 43 46 57
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 62 11 63
rect 2 60 7 62
rect 9 60 11 62
rect 2 59 11 60
rect 2 22 6 59
rect 18 49 30 55
rect 34 49 46 55
rect 10 30 14 47
rect 18 41 24 49
rect 20 38 24 41
rect 20 36 21 38
rect 23 36 24 38
rect 20 34 24 36
rect 29 38 38 39
rect 29 36 31 38
rect 33 36 38 38
rect 29 35 38 36
rect 33 30 38 35
rect 42 38 46 49
rect 42 36 43 38
rect 45 36 46 38
rect 42 34 46 36
rect 10 28 11 30
rect 13 28 23 30
rect 10 26 23 28
rect 33 26 47 30
rect 2 21 48 22
rect 2 19 15 21
rect 17 19 44 21
rect 46 19 48 21
rect 2 18 48 19
rect -2 11 58 12
rect -2 9 4 11
rect 6 9 26 11
rect 28 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 10 17 12 23
rect 20 17 22 23
rect 32 17 34 26
rect 39 17 41 26
<< pmos >>
rect 12 43 14 70
rect 19 43 21 70
rect 29 43 31 70
rect 39 43 41 70
<< polyct1 >>
rect 21 36 23 38
rect 31 36 33 38
rect 43 36 45 38
rect 11 28 13 30
<< ndifct1 >>
rect 15 19 17 21
rect 44 19 46 21
rect 4 9 6 11
rect 26 9 28 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 7 52 9 54
rect 24 59 26 61
rect 34 66 36 68
rect 44 59 46 61
<< pdifct1 >>
rect 7 60 9 62
<< alu0 >>
rect 32 66 34 68
rect 36 66 38 68
rect 32 65 38 66
rect 22 61 48 62
rect 22 59 24 61
rect 26 59 44 61
rect 46 59 48 61
rect 22 58 48 59
rect 6 54 11 55
rect 6 52 7 54
rect 9 52 11 54
rect 6 51 11 52
<< labels >>
rlabel alu0 35 60 35 60 6 n1
rlabel alu1 4 44 4 44 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 28 20 28 6 c
rlabel alu1 12 40 12 40 6 c
rlabel alu1 20 48 20 48 6 b
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 32 36 32 6 a1
rlabel alu1 28 52 28 52 6 b
rlabel alu1 36 52 36 52 6 a2
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 20 44 20 6 z
rlabel alu1 44 28 44 28 6 a1
rlabel alu1 44 48 44 48 6 a2
<< end >>
