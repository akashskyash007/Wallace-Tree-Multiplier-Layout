magic
tech scmos
timestamp 1199203292
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 64 11 69
rect 22 59 24 64
rect 29 59 31 64
rect 36 59 38 64
rect 9 35 11 52
rect 22 46 24 49
rect 17 44 24 46
rect 17 42 19 44
rect 21 42 24 44
rect 17 40 24 42
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 9 25 11 29
rect 19 25 21 40
rect 29 39 31 49
rect 36 46 38 49
rect 36 44 43 46
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 29 25 31 33
rect 41 31 43 44
rect 41 29 47 31
rect 41 27 43 29
rect 45 27 47 29
rect 41 25 47 27
rect 41 22 43 25
rect 9 14 11 19
rect 19 15 21 19
rect 29 15 31 19
rect 41 11 43 16
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 23 19 25
rect 11 21 14 23
rect 16 21 19 23
rect 11 19 19 21
rect 21 23 29 25
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 31 22 39 25
rect 31 19 41 22
rect 33 16 41 19
rect 43 20 50 22
rect 43 18 46 20
rect 48 18 50 20
rect 43 16 50 18
rect 33 11 39 16
rect 33 9 35 11
rect 37 9 39 11
rect 33 7 39 9
<< pdif >>
rect 13 71 20 73
rect 13 69 15 71
rect 17 69 20 71
rect 13 64 20 69
rect 2 62 9 64
rect 2 60 4 62
rect 6 60 9 62
rect 2 58 9 60
rect 4 52 9 58
rect 11 59 20 64
rect 11 52 22 59
rect 13 49 22 52
rect 24 49 29 59
rect 31 49 36 59
rect 38 55 43 59
rect 38 53 45 55
rect 38 51 41 53
rect 43 51 45 53
rect 38 49 45 51
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 15 71
rect 17 69 58 71
rect -2 68 58 69
rect 2 62 15 63
rect 2 60 4 62
rect 6 60 15 62
rect 2 58 15 60
rect 2 23 6 58
rect 17 44 31 46
rect 17 42 19 44
rect 21 42 31 44
rect 17 34 23 42
rect 41 38 47 46
rect 29 37 47 38
rect 29 35 31 37
rect 33 35 47 37
rect 29 34 47 35
rect 2 21 4 23
rect 2 17 6 21
rect 33 29 47 30
rect 33 27 43 29
rect 45 27 47 29
rect 33 26 47 27
rect -2 11 58 12
rect -2 9 35 11
rect 37 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 19 31 25
rect 41 16 43 22
<< pmos >>
rect 9 52 11 64
rect 22 49 24 59
rect 29 49 31 59
rect 36 49 38 59
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 19 42 21 44
rect 31 35 33 37
rect 43 27 45 29
<< ndifct0 >>
rect 14 21 16 23
rect 24 21 26 23
rect 46 18 48 20
<< ndifct1 >>
rect 4 21 6 23
rect 35 9 37 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 41 51 43 53
<< pdifct1 >>
rect 15 69 17 71
rect 4 60 6 62
<< alu0 >>
rect 10 53 45 54
rect 10 51 41 53
rect 43 51 45 53
rect 10 50 45 51
rect 10 33 14 50
rect 10 31 11 33
rect 13 31 14 33
rect 10 27 27 31
rect 6 19 7 25
rect 12 23 18 24
rect 12 21 14 23
rect 16 21 18 23
rect 12 12 18 21
rect 23 23 27 27
rect 23 21 24 23
rect 26 21 27 23
rect 23 20 50 21
rect 23 18 46 20
rect 48 18 50 20
rect 23 17 50 18
<< labels >>
rlabel alu0 12 40 12 40 6 zn
rlabel alu0 25 24 25 24 6 zn
rlabel alu0 36 19 36 19 6 zn
rlabel alu0 27 52 27 52 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 40 20 40 6 a
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 28 36 28 6 c
rlabel alu1 36 36 36 36 6 b
rlabel alu1 28 44 28 44 6 a
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 28 44 28 6 c
rlabel alu1 44 40 44 40 6 b
<< end >>
