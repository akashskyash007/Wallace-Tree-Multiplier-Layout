magic
tech scmos
timestamp 1199201736
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 66 11 70
rect 19 63 21 68
rect 29 63 31 68
rect 41 63 43 68
rect 19 43 21 54
rect 29 51 31 54
rect 29 49 37 51
rect 29 47 33 49
rect 35 47 37 49
rect 29 45 37 47
rect 19 41 25 43
rect 19 39 21 41
rect 23 39 25 41
rect 9 35 11 38
rect 19 37 25 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 9 26 11 29
rect 22 22 24 37
rect 29 22 31 45
rect 41 31 43 54
rect 40 29 46 31
rect 40 27 42 29
rect 44 27 46 29
rect 36 25 46 27
rect 36 22 38 25
rect 9 8 11 12
rect 22 8 24 13
rect 29 8 31 13
rect 36 8 38 13
<< ndif >>
rect 4 19 9 26
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 12 9 15
rect 11 22 20 26
rect 11 13 22 22
rect 24 13 29 22
rect 31 13 36 22
rect 38 19 43 22
rect 38 17 45 19
rect 38 15 41 17
rect 43 15 45 17
rect 38 13 45 15
rect 11 12 20 13
rect 13 7 20 12
rect 13 5 15 7
rect 17 5 20 7
rect 13 3 20 5
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 63 16 66
rect 33 67 39 69
rect 33 65 35 67
rect 37 65 39 67
rect 33 63 39 65
rect 11 61 19 63
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 21 58 29 63
rect 21 56 24 58
rect 26 56 29 58
rect 21 54 29 56
rect 31 54 41 63
rect 43 60 48 63
rect 43 58 50 60
rect 43 56 46 58
rect 48 56 50 58
rect 43 54 50 56
rect 11 38 17 54
<< alu1 >>
rect -2 67 58 72
rect -2 65 35 67
rect 37 65 58 67
rect -2 64 58 65
rect 2 49 7 59
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 2 40 4 42
rect 6 40 7 42
rect 2 38 7 40
rect 31 49 47 50
rect 31 47 33 49
rect 35 47 47 49
rect 31 46 47 47
rect 2 18 6 38
rect 17 41 31 42
rect 17 39 21 41
rect 23 39 31 41
rect 17 38 31 39
rect 41 38 47 46
rect 25 30 31 38
rect 41 29 47 34
rect 41 27 42 29
rect 44 27 47 29
rect 41 26 47 27
rect 25 22 47 26
rect 2 17 15 18
rect 2 15 4 17
rect 6 15 15 17
rect 2 14 15 15
rect -2 7 58 8
rect -2 5 15 7
rect 17 5 58 7
rect -2 0 58 5
<< nmos >>
rect 9 12 11 26
rect 22 13 24 22
rect 29 13 31 22
rect 36 13 38 22
<< pmos >>
rect 9 38 11 66
rect 19 54 21 63
rect 29 54 31 63
rect 41 54 43 63
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 33 47 35 49
rect 21 39 23 41
rect 42 27 44 29
<< ndifct0 >>
rect 41 15 43 17
<< ndifct1 >>
rect 4 15 6 17
rect 15 5 17 7
<< pdifct0 >>
rect 14 59 16 61
rect 24 56 26 58
rect 46 56 48 58
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 35 65 37 67
<< alu0 >>
rect 13 61 17 64
rect 13 59 14 61
rect 16 59 17 61
rect 13 57 17 59
rect 22 58 50 59
rect 22 56 24 58
rect 26 56 46 58
rect 48 56 50 58
rect 22 55 50 56
rect 22 50 26 55
rect 10 46 26 50
rect 10 33 14 46
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 10 22 22 26
rect 18 18 22 22
rect 18 17 45 18
rect 18 15 41 17
rect 43 15 45 17
rect 18 14 45 15
<< labels >>
rlabel alu0 12 36 12 36 6 zn
rlabel alu0 31 16 31 16 6 zn
rlabel alu0 36 57 36 57 6 zn
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 40 20 40 6 a
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 24 28 24 6 c
rlabel alu1 36 24 36 24 6 c
rlabel alu1 28 36 28 36 6 a
rlabel alu1 36 48 36 48 6 b
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 28 44 28 6 c
rlabel alu1 44 44 44 44 6 b
<< end >>
