magic
tech scmos
timestamp 1199543100
<< ab >>
rect 0 0 120 100
<< nwell >>
rect -5 48 125 105
<< pwell >>
rect -5 -5 125 48
<< poly >>
rect 35 94 37 98
rect 47 94 49 98
rect 57 94 59 98
rect 11 84 13 88
rect 23 85 25 89
rect 11 43 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 93 94 95 98
rect 105 94 107 98
rect 81 76 83 80
rect 21 51 25 53
rect 33 51 37 53
rect 21 43 23 51
rect 33 43 35 51
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 35 43
rect 27 39 29 41
rect 31 39 35 41
rect 47 43 49 55
rect 57 43 59 55
rect 81 53 83 56
rect 81 51 89 53
rect 81 49 85 51
rect 87 49 89 51
rect 81 47 89 49
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 27 37 35 39
rect 11 34 13 37
rect 21 34 23 37
rect 33 34 35 37
rect 45 37 53 39
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 45 34 47 37
rect 57 34 59 37
rect 81 35 83 47
rect 93 43 95 55
rect 105 43 107 55
rect 87 41 107 43
rect 87 39 89 41
rect 91 39 107 41
rect 87 37 107 39
rect 93 34 95 37
rect 105 34 107 37
rect 33 18 35 22
rect 45 18 47 22
rect 11 12 13 16
rect 21 13 23 17
rect 57 18 59 22
rect 81 21 83 25
rect 93 11 95 15
rect 105 11 107 15
<< ndif >>
rect 3 16 11 34
rect 13 17 21 34
rect 23 22 33 34
rect 35 22 45 34
rect 47 22 57 34
rect 59 22 67 34
rect 73 31 81 35
rect 73 29 75 31
rect 77 29 81 31
rect 73 25 81 29
rect 83 34 88 35
rect 83 31 93 34
rect 83 29 87 31
rect 89 29 93 31
rect 83 25 93 29
rect 23 21 31 22
rect 23 19 27 21
rect 29 19 31 21
rect 23 17 31 19
rect 37 21 43 22
rect 37 19 39 21
rect 41 19 43 21
rect 37 17 43 19
rect 13 16 18 17
rect 3 11 9 16
rect 49 11 55 22
rect 61 21 67 22
rect 85 21 93 25
rect 61 19 63 21
rect 65 19 67 21
rect 61 17 67 19
rect 85 19 87 21
rect 89 19 93 21
rect 85 15 93 19
rect 95 31 105 34
rect 95 29 99 31
rect 101 29 105 31
rect 95 21 105 29
rect 95 19 99 21
rect 101 19 105 21
rect 95 15 105 19
rect 107 31 115 34
rect 107 29 111 31
rect 113 29 115 31
rect 107 21 115 29
rect 107 19 111 21
rect 113 19 115 21
rect 107 15 115 19
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 85 21 89
rect 30 85 35 94
rect 15 84 23 85
rect 3 81 11 84
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 56 23 84
rect 25 81 35 85
rect 25 79 29 81
rect 31 79 35 81
rect 25 56 35 79
rect 37 71 47 94
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 13 55 18 56
rect 42 55 47 56
rect 49 55 57 94
rect 59 81 67 94
rect 85 91 93 94
rect 85 89 87 91
rect 89 89 93 91
rect 59 79 63 81
rect 65 79 67 81
rect 85 81 93 89
rect 59 55 67 79
rect 85 79 87 81
rect 89 79 93 81
rect 85 76 93 79
rect 73 61 81 76
rect 73 59 75 61
rect 77 59 81 61
rect 73 56 81 59
rect 83 56 93 76
rect 88 55 93 56
rect 95 81 105 94
rect 95 79 99 81
rect 101 79 105 81
rect 95 71 105 79
rect 95 69 99 71
rect 101 69 105 71
rect 95 61 105 69
rect 95 59 99 61
rect 101 59 105 61
rect 95 55 105 59
rect 107 91 115 94
rect 107 89 111 91
rect 113 89 115 91
rect 107 81 115 89
rect 107 79 111 81
rect 113 79 115 81
rect 107 71 115 79
rect 107 69 111 71
rect 113 69 115 71
rect 107 61 115 69
rect 107 59 111 61
rect 113 59 115 61
rect 107 55 115 59
<< alu1 >>
rect -2 93 122 100
rect -2 91 75 93
rect 77 91 122 93
rect -2 89 17 91
rect 19 89 87 91
rect 89 89 111 91
rect 113 89 122 91
rect -2 88 122 89
rect 3 81 67 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 79 63 81
rect 65 79 67 81
rect 3 78 67 79
rect 86 81 90 88
rect 86 79 87 81
rect 89 79 90 81
rect 86 77 90 79
rect 98 81 102 83
rect 98 79 99 81
rect 101 79 102 81
rect 8 41 12 73
rect 8 39 9 41
rect 11 39 12 41
rect 8 17 12 39
rect 18 41 22 73
rect 18 39 19 41
rect 21 39 22 41
rect 18 27 22 39
rect 28 41 32 73
rect 28 39 29 41
rect 31 39 32 41
rect 28 37 32 39
rect 38 71 88 72
rect 38 69 41 71
rect 43 69 88 71
rect 38 68 88 69
rect 38 32 42 68
rect 28 28 42 32
rect 48 41 52 63
rect 48 39 49 41
rect 51 39 52 41
rect 28 22 32 28
rect 48 27 52 39
rect 58 41 62 63
rect 58 39 59 41
rect 61 39 62 41
rect 58 27 62 39
rect 74 61 78 63
rect 74 59 75 61
rect 77 59 78 61
rect 74 42 78 59
rect 84 51 88 68
rect 84 49 85 51
rect 87 49 88 51
rect 84 47 88 49
rect 98 71 102 79
rect 98 69 99 71
rect 101 69 102 71
rect 98 61 102 69
rect 98 59 99 61
rect 101 59 102 61
rect 74 41 93 42
rect 74 39 89 41
rect 91 39 93 41
rect 74 38 93 39
rect 74 31 78 38
rect 74 29 75 31
rect 77 29 78 31
rect 74 27 78 29
rect 86 31 90 33
rect 86 29 87 31
rect 89 29 90 31
rect 25 21 32 22
rect 25 19 27 21
rect 29 19 32 21
rect 25 18 32 19
rect 37 21 67 22
rect 37 19 39 21
rect 41 19 63 21
rect 65 19 67 21
rect 37 18 67 19
rect 86 21 90 29
rect 86 19 87 21
rect 89 19 90 21
rect 86 12 90 19
rect 98 31 102 59
rect 110 81 114 88
rect 110 79 111 81
rect 113 79 114 81
rect 110 71 114 79
rect 110 69 111 71
rect 113 69 114 71
rect 110 61 114 69
rect 110 59 111 61
rect 113 59 114 61
rect 110 57 114 59
rect 98 29 99 31
rect 101 29 102 31
rect 98 21 102 29
rect 98 19 99 21
rect 101 19 102 21
rect 98 17 102 19
rect 110 31 114 33
rect 110 29 111 31
rect 113 29 114 31
rect 110 21 114 29
rect 110 19 111 21
rect 113 19 114 21
rect 110 12 114 19
rect -2 11 122 12
rect -2 9 5 11
rect 7 9 51 11
rect 53 9 122 11
rect -2 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 122 9
rect -2 5 63 7
rect 65 5 75 7
rect 77 5 87 7
rect 89 5 99 7
rect 101 5 111 7
rect 113 5 122 7
rect -2 0 122 5
<< ptie >>
rect 21 9 43 11
rect 21 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 43 9
rect 61 7 115 9
rect 21 5 43 7
rect 61 5 63 7
rect 65 5 75 7
rect 77 5 87 7
rect 89 5 99 7
rect 101 5 111 7
rect 113 5 115 7
rect 61 3 115 5
<< ntie >>
rect 73 93 79 95
rect 73 91 75 93
rect 77 91 79 93
rect 73 84 79 91
<< nmos >>
rect 11 16 13 34
rect 21 17 23 34
rect 33 22 35 34
rect 45 22 47 34
rect 57 22 59 34
rect 81 25 83 35
rect 93 15 95 34
rect 105 15 107 34
<< pmos >>
rect 11 55 13 84
rect 23 56 25 85
rect 35 56 37 94
rect 47 55 49 94
rect 57 55 59 94
rect 81 56 83 76
rect 93 55 95 94
rect 105 55 107 94
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 85 49 87 51
rect 49 39 51 41
rect 59 39 61 41
rect 89 39 91 41
<< ndifct1 >>
rect 75 29 77 31
rect 87 29 89 31
rect 27 19 29 21
rect 39 19 41 21
rect 63 19 65 21
rect 87 19 89 21
rect 99 29 101 31
rect 99 19 101 21
rect 111 29 113 31
rect 111 19 113 21
rect 5 9 7 11
rect 51 9 53 11
<< ntiect1 >>
rect 75 91 77 93
<< ptiect1 >>
rect 23 7 25 9
rect 31 7 33 9
rect 39 7 41 9
rect 63 5 65 7
rect 75 5 77 7
rect 87 5 89 7
rect 99 5 101 7
rect 111 5 113 7
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 29 79 31 81
rect 41 69 43 71
rect 87 89 89 91
rect 63 79 65 81
rect 87 79 89 81
rect 75 59 77 61
rect 99 79 101 81
rect 99 69 101 71
rect 99 59 101 61
rect 111 89 113 91
rect 111 79 113 81
rect 111 69 113 71
rect 111 59 113 61
<< labels >>
rlabel alu1 10 45 10 45 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 30 55 30 55 6 i4
rlabel alu1 60 6 60 6 6 vss
rlabel alu1 60 45 60 45 6 i3
rlabel alu1 60 94 60 94 6 vdd
rlabel alu1 100 50 100 50 6 nq
<< end >>
