magic
tech scmos
timestamp 1199203670
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 32 68 34 73
rect 39 68 41 73
rect 49 68 51 73
rect 59 68 61 73
rect 9 61 11 65
rect 22 63 24 68
rect 9 40 11 50
rect 22 47 24 50
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 19 41 25 43
rect 49 47 51 55
rect 49 45 55 47
rect 49 43 51 45
rect 53 43 55 45
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 9 26 11 34
rect 21 26 23 41
rect 32 39 34 42
rect 39 39 41 42
rect 49 41 55 43
rect 49 39 51 41
rect 29 37 35 39
rect 39 37 51 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 32 30 34 33
rect 42 30 44 37
rect 59 35 61 55
rect 65 43 71 45
rect 65 41 67 43
rect 69 41 71 43
rect 65 39 71 41
rect 57 33 64 35
rect 57 31 59 33
rect 61 31 64 33
rect 9 15 11 20
rect 57 29 64 31
rect 62 25 64 29
rect 69 25 71 39
rect 21 11 23 16
rect 32 15 34 20
rect 42 15 44 20
rect 62 10 64 15
rect 69 10 71 15
<< ndif >>
rect 25 26 32 30
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 11 20 21 26
rect 13 18 15 20
rect 17 18 21 20
rect 13 16 21 18
rect 23 20 32 26
rect 34 28 42 30
rect 34 26 37 28
rect 39 26 42 28
rect 34 20 42 26
rect 44 26 49 30
rect 44 24 51 26
rect 44 22 47 24
rect 49 22 51 24
rect 44 20 51 22
rect 23 18 26 20
rect 28 18 30 20
rect 23 16 30 18
rect 55 19 62 25
rect 55 17 57 19
rect 59 17 62 19
rect 55 15 62 17
rect 64 15 69 25
rect 71 23 78 25
rect 71 21 74 23
rect 76 21 78 23
rect 71 19 78 21
rect 71 15 76 19
<< pdif >>
rect 27 63 32 68
rect 13 61 22 63
rect 4 56 9 61
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 11 59 15 61
rect 17 59 22 61
rect 11 50 22 59
rect 24 54 32 63
rect 24 52 27 54
rect 29 52 32 54
rect 24 50 32 52
rect 27 42 32 50
rect 34 42 39 68
rect 41 65 49 68
rect 41 63 44 65
rect 46 63 49 65
rect 41 55 49 63
rect 51 60 59 68
rect 51 58 54 60
rect 56 58 59 60
rect 51 55 59 58
rect 61 63 67 68
rect 61 61 68 63
rect 61 59 64 61
rect 66 59 68 61
rect 61 55 68 59
rect 41 42 47 55
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 2 54 7 56
rect 2 52 4 54
rect 6 52 7 54
rect 2 50 7 52
rect 2 30 6 50
rect 49 45 70 46
rect 49 43 51 45
rect 53 43 70 45
rect 49 42 67 43
rect 66 41 67 42
rect 69 41 70 43
rect 29 37 62 38
rect 29 35 31 37
rect 33 35 62 37
rect 29 34 62 35
rect 2 26 15 30
rect 58 33 62 34
rect 66 33 70 41
rect 58 31 59 33
rect 61 31 62 33
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 17 7 22
rect 58 25 62 31
rect -2 1 82 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 9 20 11 26
rect 21 16 23 26
rect 32 20 34 30
rect 42 20 44 30
rect 62 15 64 25
rect 69 15 71 25
<< pmos >>
rect 9 50 11 61
rect 22 50 24 63
rect 32 42 34 68
rect 39 42 41 68
rect 49 55 51 68
rect 59 55 61 68
<< polyct0 >>
rect 21 43 23 45
rect 11 36 13 38
<< polyct1 >>
rect 51 43 53 45
rect 31 35 33 37
rect 67 41 69 43
rect 59 31 61 33
<< ndifct0 >>
rect 15 18 17 20
rect 37 26 39 28
rect 47 22 49 24
rect 26 18 28 20
rect 57 17 59 19
rect 74 21 76 23
<< ndifct1 >>
rect 4 22 6 24
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 15 59 17 61
rect 27 52 29 54
rect 44 63 46 65
rect 54 58 56 60
rect 64 59 66 61
<< pdifct1 >>
rect 4 52 6 54
<< alu0 >>
rect 13 61 19 68
rect 43 65 47 68
rect 43 63 44 65
rect 46 63 47 65
rect 43 61 47 63
rect 13 59 15 61
rect 17 59 19 61
rect 13 58 19 59
rect 53 60 57 62
rect 53 58 54 60
rect 56 58 57 60
rect 62 61 68 68
rect 62 59 64 61
rect 66 59 68 61
rect 62 58 68 59
rect 10 54 31 55
rect 53 54 57 58
rect 10 52 27 54
rect 29 52 31 54
rect 10 51 31 52
rect 10 38 14 51
rect 34 50 78 54
rect 34 46 38 50
rect 19 45 38 46
rect 19 43 21 45
rect 23 43 38 45
rect 19 42 38 43
rect 10 36 11 38
rect 13 36 22 38
rect 10 34 22 36
rect 18 29 22 34
rect 18 28 41 29
rect 18 26 37 28
rect 39 26 41 28
rect 18 25 41 26
rect 46 24 50 26
rect 74 25 78 50
rect 46 22 47 24
rect 49 22 50 24
rect 46 21 50 22
rect 73 23 78 25
rect 73 21 74 23
rect 76 21 78 23
rect 13 20 19 21
rect 13 18 15 20
rect 17 18 19 20
rect 13 12 19 18
rect 24 20 50 21
rect 24 18 26 20
rect 28 18 50 20
rect 24 17 50 18
rect 56 19 60 21
rect 73 19 78 21
rect 56 17 57 19
rect 59 17 60 19
rect 56 12 60 17
<< labels >>
rlabel alu0 12 44 12 44 6 n5
rlabel alu0 28 44 28 44 6 n2
rlabel alu0 20 53 20 53 6 n5
rlabel alu0 48 21 48 21 6 n4
rlabel alu0 37 19 37 19 6 n4
rlabel alu0 29 27 29 27 6 n5
rlabel alu0 55 56 55 56 6 n2
rlabel alu0 76 36 76 36 6 n2
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 36 36 36 36 6 b
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 44 36 44 36 6 b
rlabel alu1 52 36 52 36 6 b
rlabel polyct1 52 44 52 44 6 a
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 28 60 28 6 b
rlabel alu1 68 36 68 36 6 a
rlabel alu1 60 44 60 44 6 a
<< end >>
