magic
tech scmos
timestamp 1199202074
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 30 11 33
rect 19 30 21 33
rect 9 11 11 16
rect 19 11 21 16
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 16 9 19
rect 11 20 19 30
rect 11 18 14 20
rect 16 18 19 20
rect 11 16 19 18
rect 21 28 28 30
rect 21 26 24 28
rect 26 26 28 28
rect 21 21 28 26
rect 21 19 24 21
rect 26 19 28 21
rect 21 16 28 19
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 19 70
rect 11 66 14 68
rect 16 66 19 68
rect 11 42 19 66
rect 21 55 26 70
rect 21 53 28 55
rect 21 51 24 53
rect 26 51 28 53
rect 21 49 28 51
rect 21 42 26 49
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 62 7 63
rect 2 58 15 62
rect 2 53 6 58
rect 2 51 4 53
rect 2 46 6 51
rect 2 44 4 46
rect 2 30 6 44
rect 26 39 30 47
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 18 37 30 39
rect 18 35 21 37
rect 23 35 30 37
rect 18 33 30 35
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 21 35 23 37
<< ndifct0 >>
rect 14 18 16 20
rect 24 26 26 28
rect 24 19 26 21
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 14 66 16 68
rect 24 51 26 53
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 12 66 14 68
rect 16 66 18 68
rect 12 65 18 66
rect 6 42 7 58
rect 10 53 28 54
rect 10 51 24 53
rect 26 51 28 53
rect 10 50 28 51
rect 10 37 14 50
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 10 28 28 29
rect 10 26 24 28
rect 26 26 28 28
rect 10 25 28 26
rect 23 21 28 25
rect 12 20 18 21
rect 12 18 14 20
rect 16 18 18 20
rect 12 12 18 18
rect 23 19 24 21
rect 26 19 28 21
rect 23 17 28 19
<< labels >>
rlabel alu0 12 39 12 39 6 an
rlabel alu0 25 23 25 23 6 an
rlabel alu0 19 52 19 52 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 12 60 12 60 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 40 28 40 6 a
<< end >>
