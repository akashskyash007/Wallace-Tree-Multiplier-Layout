magic
tech scmos
timestamp 1199201789
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 10 70 12 74
rect 17 70 19 74
rect 27 70 29 74
rect 37 70 39 74
rect 10 39 12 42
rect 2 37 12 39
rect 2 35 4 37
rect 6 35 12 37
rect 2 33 12 35
rect 17 39 19 42
rect 27 39 29 42
rect 37 39 39 42
rect 17 37 23 39
rect 17 35 19 37
rect 21 35 23 37
rect 17 33 23 35
rect 27 37 33 39
rect 27 35 29 37
rect 31 35 33 37
rect 27 33 33 35
rect 37 37 46 39
rect 37 35 42 37
rect 44 35 46 37
rect 37 33 46 35
rect 10 30 12 33
rect 20 30 22 33
rect 10 19 12 24
rect 20 20 22 24
rect 30 23 32 33
rect 37 23 39 33
rect 30 9 32 14
rect 37 9 39 14
<< ndif >>
rect 2 24 10 30
rect 12 28 20 30
rect 12 26 15 28
rect 17 26 20 28
rect 12 24 20 26
rect 22 24 28 30
rect 2 14 8 24
rect 24 23 28 24
rect 24 18 30 23
rect 2 12 4 14
rect 6 12 8 14
rect 2 10 8 12
rect 22 14 30 18
rect 32 14 37 23
rect 39 21 46 23
rect 39 19 42 21
rect 44 19 46 21
rect 39 17 46 19
rect 39 14 44 17
rect 22 12 24 14
rect 26 12 28 14
rect 22 10 28 12
<< pdif >>
rect 5 55 10 70
rect 3 53 10 55
rect 3 51 5 53
rect 7 51 10 53
rect 3 46 10 51
rect 3 44 5 46
rect 7 44 10 46
rect 3 42 10 44
rect 12 42 17 70
rect 19 61 27 70
rect 19 59 22 61
rect 24 59 27 61
rect 19 42 27 59
rect 29 68 37 70
rect 29 66 32 68
rect 34 66 37 68
rect 29 42 37 66
rect 39 63 44 70
rect 39 61 46 63
rect 39 59 42 61
rect 44 59 46 61
rect 39 57 46 59
rect 39 42 44 57
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 2 55 6 63
rect 2 53 8 55
rect 2 51 5 53
rect 7 51 8 53
rect 2 47 8 51
rect 18 49 30 55
rect 34 49 46 55
rect 2 46 14 47
rect 2 44 5 46
rect 7 44 14 46
rect 2 43 14 44
rect 2 37 6 39
rect 2 35 4 37
rect 2 22 6 35
rect 10 26 14 43
rect 18 37 22 49
rect 18 35 19 37
rect 21 35 22 37
rect 18 33 22 35
rect 26 37 34 39
rect 26 35 29 37
rect 31 35 34 37
rect 26 33 34 35
rect 40 37 46 49
rect 40 35 42 37
rect 44 35 46 37
rect 40 34 46 35
rect 30 30 34 33
rect 20 22 24 29
rect 30 26 39 30
rect 2 18 15 22
rect 20 21 46 22
rect 20 19 42 21
rect 44 19 46 21
rect 20 18 46 19
rect -2 1 50 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 10 24 12 30
rect 20 24 22 30
rect 30 14 32 23
rect 37 14 39 23
<< pmos >>
rect 10 42 12 70
rect 17 42 19 70
rect 27 42 29 70
rect 37 42 39 70
<< polyct1 >>
rect 4 35 6 37
rect 19 35 21 37
rect 29 35 31 37
rect 42 35 44 37
<< ndifct0 >>
rect 15 26 17 28
rect 4 12 6 14
rect 24 12 26 14
<< ndifct1 >>
rect 42 19 44 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 22 59 24 61
rect 32 66 34 68
rect 42 59 44 61
<< pdifct1 >>
rect 5 51 7 53
rect 5 44 7 46
<< alu0 >>
rect 30 66 32 68
rect 34 66 36 68
rect 30 65 36 66
rect 20 61 46 62
rect 20 59 22 61
rect 24 59 42 61
rect 44 59 46 61
rect 20 58 46 59
rect 6 33 7 39
rect 14 29 24 30
rect 14 28 20 29
rect 14 26 15 28
rect 17 26 20 28
rect 10 25 20 26
rect 2 14 8 15
rect 2 12 4 14
rect 6 12 8 14
rect 22 14 28 15
rect 22 12 24 14
rect 26 12 28 14
<< labels >>
rlabel alu0 33 60 33 60 6 n1
rlabel alu1 4 32 4 32 6 c
rlabel alu1 4 56 4 56 6 z
rlabel alu1 12 20 12 20 6 c
rlabel alu1 12 36 12 36 6 z
rlabel alu1 20 44 20 44 6 b
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 36 28 36 6 a1
rlabel alu1 28 52 28 52 6 b
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 36 52 36 52 6 a2
rlabel alu1 44 48 44 48 6 a2
<< end >>
