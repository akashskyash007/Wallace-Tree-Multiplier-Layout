magic
tech scmos
timestamp 1199203060
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 18 70 20 74
rect 25 70 27 74
rect 32 70 34 74
rect 39 70 41 74
rect 18 45 20 48
rect 9 43 20 45
rect 9 41 11 43
rect 13 41 15 43
rect 9 39 15 41
rect 25 39 27 48
rect 9 25 11 39
rect 19 37 27 39
rect 19 35 21 37
rect 23 36 27 37
rect 23 35 25 36
rect 19 33 25 35
rect 19 25 21 33
rect 32 32 34 48
rect 39 45 41 48
rect 39 43 47 45
rect 39 41 43 43
rect 45 41 47 43
rect 39 39 47 41
rect 29 30 35 32
rect 29 28 31 30
rect 33 28 35 30
rect 29 26 35 28
rect 29 23 31 26
rect 39 23 41 39
rect 9 15 11 19
rect 19 15 21 19
rect 29 12 31 17
rect 39 12 41 17
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 23 19 25
rect 11 21 14 23
rect 16 21 19 23
rect 11 19 19 21
rect 21 23 27 25
rect 21 19 29 23
rect 23 17 29 19
rect 31 21 39 23
rect 31 19 34 21
rect 36 19 39 21
rect 31 17 39 19
rect 41 17 50 23
rect 23 13 27 17
rect 21 11 27 13
rect 21 9 23 11
rect 25 9 27 11
rect 21 7 27 9
rect 44 11 50 17
rect 44 9 46 11
rect 48 9 50 11
rect 44 7 50 9
<< pdif >>
rect 13 63 18 70
rect 11 61 18 63
rect 11 59 13 61
rect 15 59 18 61
rect 11 57 18 59
rect 13 48 18 57
rect 20 48 25 70
rect 27 48 32 70
rect 34 48 39 70
rect 41 68 48 70
rect 41 66 44 68
rect 46 66 48 68
rect 41 60 48 66
rect 41 58 44 60
rect 46 58 48 60
rect 41 48 48 58
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 61 17 63
rect 2 59 13 61
rect 15 59 17 61
rect 2 58 17 59
rect 2 34 6 58
rect 10 50 23 54
rect 10 43 14 50
rect 34 46 38 63
rect 10 41 11 43
rect 13 41 14 43
rect 10 39 14 41
rect 22 42 38 46
rect 42 43 46 47
rect 42 41 43 43
rect 45 41 46 43
rect 42 38 46 41
rect 2 30 17 34
rect 33 34 46 38
rect 13 23 17 30
rect 25 28 31 30
rect 33 28 47 30
rect 25 26 47 28
rect 13 21 14 23
rect 16 22 17 23
rect 16 21 38 22
rect 13 19 34 21
rect 36 19 38 21
rect 13 18 38 19
rect 42 17 47 26
rect -2 11 58 12
rect -2 9 23 11
rect 25 9 46 11
rect 48 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 17 31 23
rect 39 17 41 23
<< pmos >>
rect 18 48 20 70
rect 25 48 27 70
rect 32 48 34 70
rect 39 48 41 70
<< polyct0 >>
rect 21 35 23 37
<< polyct1 >>
rect 11 41 13 43
rect 43 41 45 43
rect 31 28 33 30
<< ndifct0 >>
rect 4 21 6 23
<< ndifct1 >>
rect 14 21 16 23
rect 34 19 36 21
rect 23 9 25 11
rect 46 9 48 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 44 66 46 68
rect 44 58 46 60
<< pdifct1 >>
rect 13 59 15 61
<< alu0 >>
rect 43 66 44 68
rect 46 66 47 68
rect 43 60 47 66
rect 43 58 44 60
rect 46 58 47 60
rect 43 56 47 58
rect 20 42 22 46
rect 20 37 24 42
rect 20 35 21 37
rect 23 35 24 37
rect 20 33 24 35
rect 29 30 35 31
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 12 7 21
<< labels >>
rlabel alu1 4 48 4 48 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 44 12 44 6 d
rlabel alu1 20 52 20 52 6 d
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 b
rlabel alu1 36 36 36 36 6 a
rlabel alu1 36 28 36 28 6 b
rlabel alu1 28 44 28 44 6 c
rlabel alu1 36 56 36 56 6 c
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 24 44 24 6 b
rlabel alu1 44 44 44 44 6 a
<< end >>
