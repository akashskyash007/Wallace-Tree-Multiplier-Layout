magic
tech scmos
timestamp 1199202576
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 49 66 51 71
rect 59 66 61 71
rect 69 66 71 71
rect 79 58 81 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 79 39 81 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 33 39
rect 19 35 28 37
rect 30 35 33 37
rect 19 33 33 35
rect 12 30 14 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 37 51 39
rect 38 35 40 37
rect 42 35 47 37
rect 49 35 51 37
rect 38 33 51 35
rect 55 37 62 39
rect 55 35 58 37
rect 60 35 62 37
rect 55 33 62 35
rect 66 37 81 39
rect 66 35 77 37
rect 79 35 81 37
rect 66 33 81 35
rect 38 30 40 33
rect 48 30 50 33
rect 55 30 57 33
rect 66 30 68 33
rect 12 6 14 10
rect 19 6 21 10
rect 31 6 33 10
rect 38 6 40 10
rect 48 6 50 10
rect 55 6 57 10
rect 66 6 68 10
<< ndif >>
rect 5 28 12 30
rect 5 26 7 28
rect 9 26 12 28
rect 5 21 12 26
rect 5 19 7 21
rect 9 19 12 21
rect 5 17 12 19
rect 7 10 12 17
rect 14 10 19 30
rect 21 14 31 30
rect 21 12 25 14
rect 27 12 31 14
rect 21 10 31 12
rect 33 10 38 30
rect 40 28 48 30
rect 40 26 43 28
rect 45 26 48 28
rect 40 21 48 26
rect 40 19 43 21
rect 45 19 48 21
rect 40 10 48 19
rect 50 10 55 30
rect 57 21 66 30
rect 57 19 61 21
rect 63 19 66 21
rect 57 14 66 19
rect 57 12 61 14
rect 63 12 66 14
rect 57 10 66 12
rect 68 28 75 30
rect 68 26 71 28
rect 73 26 75 28
rect 68 21 75 26
rect 68 19 71 21
rect 73 19 75 21
rect 68 17 75 19
rect 68 10 73 17
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 42 9 62
rect 11 61 19 66
rect 11 59 14 61
rect 16 59 19 61
rect 11 53 19 59
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 42 29 62
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 42 49 62
rect 51 61 59 66
rect 51 59 54 61
rect 56 59 59 61
rect 51 54 59 59
rect 51 52 54 54
rect 56 52 59 54
rect 51 42 59 52
rect 61 64 69 66
rect 61 62 64 64
rect 66 62 69 64
rect 61 56 69 62
rect 61 54 64 56
rect 66 54 69 56
rect 61 42 69 54
rect 71 58 76 66
rect 71 53 79 58
rect 71 51 74 53
rect 76 51 79 53
rect 71 46 79 51
rect 71 44 74 46
rect 76 44 79 46
rect 71 42 79 44
rect 81 56 89 58
rect 81 54 84 56
rect 86 54 89 56
rect 81 48 89 54
rect 81 46 84 48
rect 86 46 89 48
rect 81 42 89 46
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 68 98 79
rect 33 61 38 63
rect 2 54 15 55
rect 33 59 34 61
rect 36 59 38 61
rect 53 61 57 63
rect 33 54 38 59
rect 53 59 54 61
rect 56 59 57 61
rect 53 54 57 59
rect 2 53 54 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 52 54 53
rect 56 52 57 54
rect 36 51 57 52
rect 2 50 57 51
rect 2 29 6 50
rect 17 39 23 46
rect 10 37 23 39
rect 10 35 11 37
rect 13 35 23 37
rect 10 33 23 35
rect 35 37 51 38
rect 35 35 40 37
rect 42 35 47 37
rect 49 35 51 37
rect 35 34 51 35
rect 17 30 23 33
rect 35 30 39 34
rect 74 37 86 39
rect 74 35 77 37
rect 79 35 86 37
rect 74 33 86 35
rect 2 28 11 29
rect 2 26 7 28
rect 9 26 11 28
rect 17 26 39 30
rect 2 25 11 26
rect 7 22 11 25
rect 7 21 47 22
rect 9 19 43 21
rect 45 19 47 21
rect 7 18 47 19
rect 82 17 86 33
rect -2 1 98 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 31 10 33 30
rect 38 10 40 30
rect 48 10 50 30
rect 55 10 57 30
rect 66 10 68 30
<< pmos >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
rect 49 42 51 66
rect 59 42 61 66
rect 69 42 71 66
rect 79 42 81 58
<< polyct0 >>
rect 28 35 30 37
rect 58 35 60 37
<< polyct1 >>
rect 11 35 13 37
rect 40 35 42 37
rect 47 35 49 37
rect 77 35 79 37
<< ndifct0 >>
rect 25 12 27 14
rect 43 26 45 28
rect 61 19 63 21
rect 61 12 63 14
rect 71 26 73 28
rect 71 19 73 21
<< ndifct1 >>
rect 7 26 9 28
rect 7 19 9 21
rect 43 19 45 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 62 6 64
rect 14 59 16 61
rect 24 62 26 64
rect 44 62 46 64
rect 64 62 66 64
rect 64 54 66 56
rect 74 51 76 53
rect 74 44 76 46
rect 84 54 86 56
rect 84 46 86 48
<< pdifct1 >>
rect 14 51 16 53
rect 34 59 36 61
rect 34 51 36 53
rect 54 59 56 61
rect 54 52 56 54
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 23 64 27 68
rect 3 60 7 62
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 23 62 24 64
rect 26 62 27 64
rect 43 64 47 68
rect 23 60 27 62
rect 13 55 17 59
rect 15 54 17 55
rect 43 62 44 64
rect 46 62 47 64
rect 63 64 67 68
rect 43 60 47 62
rect 63 62 64 64
rect 66 62 67 64
rect 63 56 67 62
rect 63 54 64 56
rect 66 54 67 56
rect 83 56 87 68
rect 63 52 67 54
rect 73 53 77 55
rect 73 51 74 53
rect 76 51 77 53
rect 73 46 77 51
rect 27 44 74 46
rect 76 44 77 46
rect 83 54 84 56
rect 86 54 87 56
rect 83 48 87 54
rect 83 46 84 48
rect 86 46 87 48
rect 83 44 87 46
rect 27 42 77 44
rect 27 37 31 42
rect 27 35 28 37
rect 30 35 31 37
rect 27 33 31 35
rect 57 37 61 42
rect 57 35 58 37
rect 60 35 61 37
rect 57 30 61 35
rect 42 28 47 30
rect 42 26 43 28
rect 45 26 47 28
rect 57 28 74 30
rect 57 26 71 28
rect 73 26 74 28
rect 5 18 7 25
rect 42 22 47 26
rect 59 21 65 22
rect 59 19 61 21
rect 63 19 65 21
rect 23 14 29 15
rect 23 12 25 14
rect 27 12 29 14
rect 59 14 65 19
rect 70 21 74 26
rect 70 19 71 21
rect 73 19 74 21
rect 70 17 74 19
rect 59 12 61 14
rect 63 12 65 14
<< labels >>
rlabel alu0 29 39 29 39 6 an
rlabel polyct0 59 36 59 36 6 an
rlabel alu0 72 23 72 23 6 an
rlabel alu0 75 48 75 48 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 36 20 36 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 4 40 4 40 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel ndifct1 44 20 44 20 6 z
rlabel alu1 44 36 44 36 6 b
rlabel alu1 36 28 36 28 6 b
rlabel alu1 28 28 28 28 6 b
rlabel alu1 36 56 36 56 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel alu1 52 52 52 52 6 z
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 76 36 76 36 6 a
rlabel alu1 84 28 84 28 6 a
<< end >>
