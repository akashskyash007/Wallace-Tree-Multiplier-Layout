magic
tech scmos
timestamp 1199542410
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -2 48 102 104
<< pwell >>
rect -2 -4 102 48
<< poly >>
rect 23 95 25 98
rect 35 95 37 98
rect 11 75 13 78
rect 51 85 53 88
rect 63 85 65 88
rect 75 85 77 88
rect 87 85 89 88
rect 11 53 13 55
rect 11 51 19 53
rect 11 49 15 51
rect 17 49 19 51
rect 11 47 19 49
rect 23 43 25 55
rect 35 43 37 55
rect 9 41 37 43
rect 9 39 11 41
rect 13 39 37 41
rect 9 37 37 39
rect 11 31 19 33
rect 11 29 15 31
rect 17 29 19 31
rect 11 27 19 29
rect 11 25 13 27
rect 23 25 25 37
rect 35 25 37 37
rect 51 33 53 65
rect 63 63 65 65
rect 59 61 65 63
rect 59 43 61 61
rect 75 53 77 65
rect 67 51 77 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 47 31 53 33
rect 47 29 49 31
rect 51 29 53 31
rect 47 27 53 29
rect 51 25 53 27
rect 59 25 61 37
rect 67 25 69 47
rect 77 41 83 43
rect 77 39 79 41
rect 81 39 83 41
rect 87 39 89 65
rect 75 37 89 39
rect 75 25 77 37
rect 11 12 13 15
rect 23 2 25 5
rect 35 2 37 5
rect 51 2 53 5
rect 59 2 61 5
rect 67 2 69 5
rect 75 2 77 5
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 15 11 23 15
rect 15 9 17 11
rect 19 9 23 11
rect 15 5 23 9
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 5 35 19
rect 37 11 51 25
rect 37 9 43 11
rect 45 9 51 11
rect 37 5 51 9
rect 53 5 59 25
rect 61 5 67 25
rect 69 5 75 25
rect 77 21 93 25
rect 77 19 89 21
rect 91 19 93 21
rect 77 15 93 19
rect 77 5 85 15
<< pdif >>
rect 15 91 23 95
rect 15 89 17 91
rect 19 89 23 91
rect 15 75 23 89
rect 3 71 11 75
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 55 23 75
rect 25 71 35 95
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 91 49 95
rect 37 89 43 91
rect 45 89 49 91
rect 37 85 49 89
rect 67 91 73 93
rect 67 89 69 91
rect 71 89 73 91
rect 67 85 73 89
rect 91 91 97 93
rect 91 89 93 91
rect 95 89 97 91
rect 91 85 97 89
rect 37 65 51 85
rect 53 81 63 85
rect 53 79 57 81
rect 59 79 63 81
rect 53 65 63 79
rect 65 65 75 85
rect 77 81 87 85
rect 77 79 81 81
rect 83 79 87 81
rect 77 65 87 79
rect 89 65 97 85
rect 37 55 45 65
<< alu1 >>
rect -2 95 102 100
rect -2 93 5 95
rect 7 93 102 95
rect -2 91 102 93
rect -2 89 17 91
rect 19 89 43 91
rect 45 89 69 91
rect 71 89 93 91
rect 95 89 102 91
rect -2 88 102 89
rect 56 81 60 82
rect 80 81 84 82
rect 20 79 57 81
rect 59 79 81 81
rect 83 79 92 81
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 62 7 68
rect 4 61 8 62
rect 4 59 5 61
rect 7 59 8 61
rect 4 58 8 59
rect 5 42 7 58
rect 20 52 22 79
rect 56 78 60 79
rect 80 78 84 79
rect 14 51 22 52
rect 14 49 15 51
rect 17 49 22 51
rect 14 48 22 49
rect 5 41 14 42
rect 5 39 11 41
rect 13 39 14 41
rect 5 38 14 39
rect 5 22 7 38
rect 20 32 22 48
rect 14 31 22 32
rect 14 29 15 31
rect 17 29 22 31
rect 14 28 22 29
rect 28 71 32 72
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 4 21 8 22
rect 4 19 5 21
rect 7 19 8 21
rect 4 18 8 19
rect 28 21 32 59
rect 28 19 29 21
rect 31 19 32 21
rect 28 18 32 19
rect 48 31 52 72
rect 48 29 49 31
rect 51 29 52 31
rect 48 18 52 29
rect 58 41 62 72
rect 58 39 59 41
rect 61 39 62 41
rect 58 18 62 39
rect 68 51 72 72
rect 68 49 69 51
rect 71 49 72 51
rect 68 18 72 49
rect 78 41 82 72
rect 78 39 79 41
rect 81 39 82 41
rect 78 18 82 39
rect 90 22 92 79
rect 88 21 92 22
rect 88 19 89 21
rect 91 19 92 21
rect 88 18 92 19
rect -2 11 102 12
rect -2 9 17 11
rect 19 9 43 11
rect 45 9 102 11
rect -2 0 102 9
<< ntie >>
rect 3 95 9 97
rect 3 93 5 95
rect 7 93 9 95
rect 3 85 9 93
<< nmos >>
rect 11 15 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 51 5 53 25
rect 59 5 61 25
rect 67 5 69 25
rect 75 5 77 25
<< pmos >>
rect 11 55 13 75
rect 23 55 25 95
rect 35 55 37 95
rect 51 65 53 85
rect 63 65 65 85
rect 75 65 77 85
rect 87 65 89 85
<< polyct1 >>
rect 15 49 17 51
rect 11 39 13 41
rect 15 29 17 31
rect 69 49 71 51
rect 59 39 61 41
rect 49 29 51 31
rect 79 39 81 41
<< ndifct1 >>
rect 5 19 7 21
rect 17 9 19 11
rect 29 19 31 21
rect 43 9 45 11
rect 89 19 91 21
<< ntiect1 >>
rect 5 93 7 95
<< pdifct1 >>
rect 17 89 19 91
rect 5 69 7 71
rect 5 59 7 61
rect 29 69 31 71
rect 29 59 31 61
rect 43 89 45 91
rect 69 89 71 91
rect 93 89 95 91
rect 57 79 59 81
rect 81 79 83 81
<< labels >>
rlabel alu1 30 45 30 45 6 nq
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 50 45 50 45 6 i0
rlabel alu1 70 45 70 45 6 i2
rlabel alu1 60 45 60 45 6 i1
rlabel alu1 50 94 50 94 6 vdd
rlabel alu1 80 45 80 45 6 i3
<< end >>
