magic
tech scmos
timestamp 1199203026
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 13 70 15 74
rect 21 70 23 74
rect 29 70 31 74
rect 39 70 41 74
rect 46 70 48 74
rect 53 70 55 74
rect 63 70 65 74
rect 70 70 72 74
rect 77 70 79 74
rect 87 61 89 66
rect 94 61 96 65
rect 101 61 103 65
rect 13 39 15 42
rect 21 39 23 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 29 37 41 39
rect 29 35 37 37
rect 39 35 41 37
rect 29 33 41 35
rect 9 30 11 33
rect 21 30 23 33
rect 31 30 33 33
rect 46 23 48 42
rect 53 39 55 42
rect 63 39 65 42
rect 53 37 65 39
rect 59 35 61 37
rect 63 35 65 37
rect 59 33 65 35
rect 70 23 72 42
rect 77 39 79 42
rect 87 39 89 42
rect 77 37 89 39
rect 77 29 83 37
rect 77 27 79 29
rect 81 27 83 29
rect 77 25 83 27
rect 94 23 96 42
rect 101 39 103 42
rect 101 37 107 39
rect 101 35 103 37
rect 105 35 107 37
rect 101 33 107 35
rect 46 21 52 23
rect 46 19 48 21
rect 50 19 52 21
rect 46 17 52 19
rect 66 21 72 23
rect 66 19 68 21
rect 70 19 72 21
rect 66 17 72 19
rect 89 21 96 23
rect 89 19 91 21
rect 93 19 96 21
rect 89 17 96 19
rect 9 6 11 11
rect 21 6 23 11
rect 31 6 33 11
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 11 9 17
rect 11 11 21 30
rect 23 21 31 30
rect 23 19 26 21
rect 28 19 31 21
rect 23 11 31 19
rect 33 22 41 30
rect 33 20 36 22
rect 38 20 41 22
rect 33 15 41 20
rect 33 13 36 15
rect 38 13 41 15
rect 33 11 41 13
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 5 68 13 70
rect 5 66 8 68
rect 10 66 13 68
rect 5 61 13 66
rect 5 59 8 61
rect 10 59 13 61
rect 5 42 13 59
rect 15 42 21 70
rect 23 42 29 70
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 42 46 70
rect 48 42 53 70
rect 55 68 63 70
rect 55 66 58 68
rect 60 66 63 68
rect 55 61 63 66
rect 55 59 58 61
rect 60 59 63 61
rect 55 42 63 59
rect 65 42 70 70
rect 72 42 77 70
rect 79 61 84 70
rect 79 53 87 61
rect 79 51 82 53
rect 84 51 87 53
rect 79 46 87 51
rect 79 44 82 46
rect 84 44 87 46
rect 79 42 87 44
rect 89 42 94 61
rect 96 42 101 61
rect 103 59 110 61
rect 103 57 106 59
rect 108 57 110 59
rect 103 52 110 57
rect 103 50 106 52
rect 108 50 110 52
rect 103 42 110 50
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 68 114 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 2 53 87 54
rect 2 51 34 53
rect 36 51 82 53
rect 84 51 87 53
rect 2 50 87 51
rect 2 29 6 50
rect 81 46 87 50
rect 10 42 63 46
rect 81 44 82 46
rect 84 44 95 46
rect 81 42 95 44
rect 10 37 14 42
rect 59 38 63 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 19 37 31 38
rect 19 35 21 37
rect 23 35 31 37
rect 19 34 31 35
rect 35 37 55 38
rect 35 35 37 37
rect 39 35 55 37
rect 35 34 55 35
rect 59 37 107 38
rect 59 35 61 37
rect 63 35 103 37
rect 105 35 107 37
rect 59 34 107 35
rect 25 30 31 34
rect 51 30 55 34
rect 2 28 8 29
rect 2 26 4 28
rect 6 26 8 28
rect 25 26 47 30
rect 51 29 87 30
rect 51 27 79 29
rect 81 27 87 29
rect 51 26 87 27
rect 2 22 8 26
rect 2 21 31 22
rect 2 19 4 21
rect 6 19 26 21
rect 28 19 31 21
rect 2 18 31 19
rect 43 22 47 26
rect 43 21 95 22
rect 43 19 48 21
rect 50 19 68 21
rect 70 19 91 21
rect 93 19 95 21
rect 43 18 95 19
rect -2 11 114 12
rect -2 9 15 11
rect 17 9 114 11
rect -2 1 114 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 9 11 11 30
rect 21 11 23 30
rect 31 11 33 30
<< pmos >>
rect 13 42 15 70
rect 21 42 23 70
rect 29 42 31 70
rect 39 42 41 70
rect 46 42 48 70
rect 53 42 55 70
rect 63 42 65 70
rect 70 42 72 70
rect 77 42 79 70
rect 87 42 89 61
rect 94 42 96 61
rect 101 42 103 61
<< polyct1 >>
rect 11 35 13 37
rect 21 35 23 37
rect 37 35 39 37
rect 61 35 63 37
rect 79 27 81 29
rect 103 35 105 37
rect 48 19 50 21
rect 68 19 70 21
rect 91 19 93 21
<< ndifct0 >>
rect 36 20 38 22
rect 36 13 38 15
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
rect 26 19 28 21
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 8 66 10 68
rect 8 59 10 61
rect 58 66 60 68
rect 58 59 60 61
rect 106 57 108 59
rect 106 50 108 52
<< pdifct1 >>
rect 34 59 36 61
rect 34 51 36 53
rect 82 51 84 53
rect 82 44 84 46
<< alu0 >>
rect 6 66 8 68
rect 10 66 12 68
rect 6 61 12 66
rect 56 66 58 68
rect 60 66 62 68
rect 6 59 8 61
rect 10 59 12 61
rect 6 58 12 59
rect 56 61 62 66
rect 56 59 58 61
rect 60 59 62 61
rect 56 58 62 59
rect 104 59 110 68
rect 104 57 106 59
rect 108 57 110 59
rect 104 52 110 57
rect 104 50 106 52
rect 108 50 110 52
rect 104 49 110 50
rect 34 22 40 23
rect 34 20 36 22
rect 38 20 40 22
rect 34 15 40 20
rect 34 13 36 15
rect 38 13 40 15
rect 34 12 40 13
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 36 28 36 28 6 b
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 32 28 32 6 b
rlabel alu1 20 44 20 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 28 44 28 44 6 a
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 56 6 56 6 6 vss
rlabel alu1 44 28 44 28 6 b
rlabel alu1 60 28 60 28 6 c
rlabel alu1 60 20 60 20 6 b
rlabel alu1 52 20 52 20 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 44 36 44 36 6 c
rlabel alu1 60 44 60 44 6 a
rlabel alu1 52 44 52 44 6 a
rlabel alu1 52 36 52 36 6 c
rlabel alu1 60 52 60 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 56 74 56 74 6 vdd
rlabel alu1 68 28 68 28 6 c
rlabel alu1 68 20 68 20 6 b
rlabel alu1 84 28 84 28 6 c
rlabel alu1 84 20 84 20 6 b
rlabel alu1 76 28 76 28 6 c
rlabel alu1 76 20 76 20 6 b
rlabel alu1 68 36 68 36 6 a
rlabel alu1 84 36 84 36 6 a
rlabel alu1 76 36 76 36 6 a
rlabel alu1 84 48 84 48 6 z
rlabel alu1 76 52 76 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel polyct1 92 20 92 20 6 b
rlabel alu1 92 44 92 44 6 z
rlabel alu1 92 36 92 36 6 a
rlabel alu1 100 36 100 36 6 a
<< end >>
