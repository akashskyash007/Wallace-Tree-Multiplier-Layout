magic
tech scmos
timestamp 1199202151
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 12 65 14 70
rect 22 65 24 70
rect 29 65 31 70
rect 39 65 41 70
rect 49 65 51 70
rect 61 65 63 70
rect 12 35 14 38
rect 22 35 24 38
rect 9 33 24 35
rect 9 31 11 33
rect 13 31 24 33
rect 29 32 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 61 35 63 38
rect 9 29 24 31
rect 28 29 31 32
rect 37 33 43 35
rect 37 31 39 33
rect 41 31 43 33
rect 37 29 43 31
rect 47 33 53 35
rect 47 31 49 33
rect 51 31 53 33
rect 47 29 53 31
rect 57 33 63 35
rect 57 31 59 33
rect 61 31 63 33
rect 57 29 63 31
rect 9 24 11 29
rect 21 26 23 29
rect 28 26 30 29
rect 38 26 40 29
rect 48 26 50 29
rect 59 26 61 29
rect 9 7 11 12
rect 21 9 23 14
rect 28 5 30 14
rect 38 9 40 14
rect 48 5 50 14
rect 59 9 61 14
rect 28 3 50 5
<< ndif >>
rect 13 24 21 26
rect 4 18 9 24
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 14 21 24
rect 23 14 28 26
rect 30 24 38 26
rect 30 22 33 24
rect 35 22 38 24
rect 30 14 38 22
rect 40 18 48 26
rect 40 16 43 18
rect 45 16 48 18
rect 40 14 48 16
rect 50 18 59 26
rect 50 16 53 18
rect 55 16 59 18
rect 50 14 59 16
rect 61 24 68 26
rect 61 22 64 24
rect 66 22 68 24
rect 61 20 68 22
rect 61 14 66 20
rect 11 12 19 14
rect 13 7 19 12
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
<< pdif >>
rect 7 59 12 65
rect 5 57 12 59
rect 5 55 7 57
rect 9 55 12 57
rect 5 50 12 55
rect 5 48 7 50
rect 9 48 12 50
rect 5 46 12 48
rect 7 38 12 46
rect 14 63 22 65
rect 14 61 17 63
rect 19 61 22 63
rect 14 56 22 61
rect 14 54 17 56
rect 19 54 22 56
rect 14 38 22 54
rect 24 38 29 65
rect 31 49 39 65
rect 31 47 34 49
rect 36 47 39 49
rect 31 42 39 47
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 58 49 65
rect 41 56 44 58
rect 46 56 49 58
rect 41 38 49 56
rect 51 63 61 65
rect 51 61 55 63
rect 57 61 61 63
rect 51 38 61 61
rect 63 51 68 65
rect 63 49 70 51
rect 63 47 66 49
rect 68 47 70 49
rect 63 42 70 47
rect 63 40 66 42
rect 68 40 70 42
rect 63 38 70 40
<< alu1 >>
rect -2 64 74 72
rect 33 49 38 51
rect 33 47 34 49
rect 36 47 38 49
rect 2 35 6 43
rect 33 42 38 47
rect 18 40 34 42
rect 36 40 38 42
rect 18 38 38 40
rect 42 41 46 51
rect 50 45 62 51
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 18 26 22 38
rect 42 37 54 41
rect 48 33 54 37
rect 48 31 49 33
rect 51 31 54 33
rect 48 29 54 31
rect 58 33 62 45
rect 58 31 59 33
rect 61 31 62 33
rect 58 29 62 31
rect 18 24 37 26
rect 18 22 33 24
rect 35 22 37 24
rect 18 21 37 22
rect -2 7 74 8
rect -2 5 15 7
rect 17 5 74 7
rect -2 0 74 5
<< nmos >>
rect 9 12 11 24
rect 21 14 23 26
rect 28 14 30 26
rect 38 14 40 26
rect 48 14 50 26
rect 59 14 61 26
<< pmos >>
rect 12 38 14 65
rect 22 38 24 65
rect 29 38 31 65
rect 39 38 41 65
rect 49 38 51 65
rect 61 38 63 65
<< polyct0 >>
rect 39 31 41 33
<< polyct1 >>
rect 11 31 13 33
rect 49 31 51 33
rect 59 31 61 33
<< ndifct0 >>
rect 4 14 6 16
rect 43 16 45 18
rect 53 16 55 18
rect 64 22 66 24
<< ndifct1 >>
rect 33 22 35 24
rect 15 5 17 7
<< pdifct0 >>
rect 7 55 9 57
rect 7 48 9 50
rect 17 61 19 63
rect 17 54 19 56
rect 44 56 46 58
rect 55 61 57 63
rect 66 47 68 49
rect 66 40 68 42
<< pdifct1 >>
rect 34 47 36 49
rect 34 40 36 42
<< alu0 >>
rect 15 63 21 64
rect 15 61 17 63
rect 19 61 21 63
rect 6 57 10 59
rect 6 55 7 57
rect 9 55 10 57
rect 6 50 10 55
rect 15 56 21 61
rect 54 63 58 64
rect 54 61 55 63
rect 57 61 58 63
rect 54 59 58 61
rect 15 54 17 56
rect 19 54 21 56
rect 15 53 21 54
rect 24 58 48 59
rect 24 56 44 58
rect 46 56 48 58
rect 24 55 48 56
rect 24 50 28 55
rect 6 48 7 50
rect 9 48 28 50
rect 6 46 28 48
rect 37 33 45 34
rect 37 31 39 33
rect 41 31 45 33
rect 37 30 45 31
rect 41 26 45 30
rect 65 49 70 51
rect 65 47 66 49
rect 68 47 70 49
rect 65 42 70 47
rect 65 40 66 42
rect 68 40 70 42
rect 65 38 70 40
rect 66 26 70 38
rect 41 24 70 26
rect 41 22 64 24
rect 66 22 70 24
rect 62 21 70 22
rect 41 18 47 19
rect 41 17 43 18
rect 2 16 43 17
rect 45 16 47 18
rect 2 14 4 16
rect 6 14 47 16
rect 2 13 47 14
rect 51 18 57 19
rect 51 16 53 18
rect 55 16 57 18
rect 51 8 57 16
<< labels >>
rlabel alu0 8 52 8 52 6 n1
rlabel alu0 24 15 24 15 6 n3
rlabel alu0 44 16 44 16 6 n3
rlabel alu0 36 57 36 57 6 n1
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 4 36 4 36 6 a
rlabel alu1 20 28 20 28 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 52 32 52 32 6 b
rlabel alu1 36 48 36 48 6 z
rlabel alu1 52 48 52 48 6 c
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 40 60 40 6 c
<< end >>
