magic
tech scmos
timestamp 1199203617
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 6 68 30 70
rect 6 59 8 68
rect 18 60 20 64
rect 28 60 30 68
rect 38 68 60 70
rect 38 60 40 68
rect 48 60 50 64
rect 58 60 60 68
rect 2 57 8 59
rect 2 55 4 57
rect 6 55 8 57
rect 2 53 8 55
rect 18 35 20 38
rect 8 33 20 35
rect 28 33 30 38
rect 38 34 40 38
rect 48 34 50 38
rect 58 35 60 38
rect 8 31 10 33
rect 12 31 14 33
rect 28 31 34 33
rect 8 29 14 31
rect 12 26 14 29
rect 22 25 24 29
rect 32 25 34 31
rect 48 32 54 34
rect 48 30 50 32
rect 52 30 54 32
rect 42 28 54 30
rect 58 33 64 35
rect 58 31 60 33
rect 62 31 64 33
rect 58 29 64 31
rect 42 25 44 28
rect 61 25 63 29
rect 12 10 14 15
rect 22 6 24 14
rect 32 10 34 14
rect 42 10 44 14
rect 61 6 63 14
rect 22 4 63 6
<< ndif >>
rect 2 19 12 26
rect 2 17 4 19
rect 6 17 12 19
rect 2 15 12 17
rect 14 25 19 26
rect 14 22 22 25
rect 14 20 17 22
rect 19 20 22 22
rect 14 15 22 20
rect 17 14 22 15
rect 24 23 32 25
rect 24 21 27 23
rect 29 21 32 23
rect 24 14 32 21
rect 34 23 42 25
rect 34 21 37 23
rect 39 21 42 23
rect 34 14 42 21
rect 44 18 61 25
rect 44 16 56 18
rect 58 16 61 18
rect 44 14 61 16
rect 63 23 70 25
rect 63 21 66 23
rect 68 21 70 23
rect 63 19 70 21
rect 63 14 68 19
<< pdif >>
rect 11 58 18 60
rect 11 56 13 58
rect 15 56 18 58
rect 11 38 18 56
rect 20 42 28 60
rect 20 40 23 42
rect 25 40 28 42
rect 20 38 28 40
rect 30 42 38 60
rect 30 40 33 42
rect 35 40 38 42
rect 30 38 38 40
rect 40 42 48 60
rect 40 40 43 42
rect 45 40 48 42
rect 40 38 48 40
rect 50 58 58 60
rect 50 56 53 58
rect 55 56 58 58
rect 50 38 58 56
rect 60 52 65 60
rect 60 50 67 52
rect 60 48 63 50
rect 65 48 67 50
rect 60 46 67 48
rect 60 38 65 46
<< alu1 >>
rect -2 64 74 72
rect 2 35 6 43
rect 30 42 38 43
rect 30 40 33 42
rect 35 40 38 42
rect 2 33 14 35
rect 2 31 10 33
rect 12 31 14 33
rect 2 29 14 31
rect 30 37 38 40
rect 30 34 34 37
rect 50 37 62 43
rect 58 35 62 37
rect 25 30 34 34
rect 25 23 31 30
rect 58 33 63 35
rect 58 31 60 33
rect 62 31 63 33
rect 58 29 63 31
rect 25 21 27 23
rect 29 21 31 23
rect 25 20 31 21
rect -2 7 74 8
rect -2 5 5 7
rect 7 5 74 7
rect -2 0 74 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< nmos >>
rect 12 15 14 26
rect 22 14 24 25
rect 32 14 34 25
rect 42 14 44 25
rect 61 14 63 25
<< pmos >>
rect 18 38 20 60
rect 28 38 30 60
rect 38 38 40 60
rect 48 38 50 60
rect 58 38 60 60
<< polyct0 >>
rect 4 55 6 57
rect 50 30 52 32
<< polyct1 >>
rect 10 31 12 33
rect 60 31 62 33
<< ndifct0 >>
rect 4 17 6 19
rect 17 20 19 22
rect 37 21 39 23
rect 56 16 58 18
rect 66 21 68 23
<< ndifct1 >>
rect 27 21 29 23
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 13 56 15 58
rect 23 40 25 42
rect 43 40 45 42
rect 53 56 55 58
rect 63 48 65 50
<< pdifct1 >>
rect 33 40 35 42
<< alu0 >>
rect 3 57 7 59
rect 3 55 4 57
rect 6 55 7 57
rect 11 58 17 64
rect 11 56 13 58
rect 15 56 17 58
rect 11 55 17 56
rect 51 58 57 64
rect 51 56 53 58
rect 55 56 57 58
rect 51 55 57 56
rect 3 51 7 55
rect 3 50 70 51
rect 3 48 63 50
rect 65 48 70 50
rect 3 47 70 48
rect 17 42 27 43
rect 17 40 23 42
rect 25 40 27 42
rect 17 39 27 40
rect 17 24 21 39
rect 42 42 46 44
rect 42 40 43 42
rect 45 40 46 42
rect 42 34 46 40
rect 16 22 21 24
rect 3 19 7 21
rect 3 17 4 19
rect 6 17 7 19
rect 16 20 17 22
rect 19 20 21 22
rect 38 30 46 34
rect 49 32 53 34
rect 49 30 50 32
rect 52 30 53 32
rect 38 24 42 30
rect 49 27 53 30
rect 35 23 42 24
rect 35 21 37 23
rect 39 21 42 23
rect 35 20 42 21
rect 47 23 53 27
rect 66 25 70 47
rect 65 23 70 25
rect 16 18 21 20
rect 3 8 7 17
rect 17 17 21 18
rect 47 17 51 23
rect 65 21 66 23
rect 68 21 70 23
rect 17 13 51 17
rect 55 18 59 20
rect 65 19 70 21
rect 55 16 56 18
rect 58 16 59 18
rect 55 8 59 16
<< labels >>
rlabel alu0 5 53 5 53 6 bn
rlabel alu0 19 28 19 28 6 an
rlabel alu0 22 41 22 41 6 an
rlabel ndifct0 38 22 38 22 6 ai
rlabel alu0 44 37 44 37 6 ai
rlabel alu0 51 28 51 28 6 an
rlabel alu0 68 35 68 35 6 bn
rlabel alu0 36 49 36 49 6 bn
rlabel alu1 12 32 12 32 6 a
rlabel alu1 4 36 4 36 6 a
rlabel alu1 28 28 28 28 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 52 40 52 40 6 b
rlabel alu1 36 40 36 40 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 36 60 36 6 b
<< end >>
