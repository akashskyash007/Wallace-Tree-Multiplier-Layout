magic
tech scmos
timestamp 1199541665
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -2 48 52 104
<< pwell >>
rect -2 -4 52 48
<< poly >>
rect 17 95 19 98
rect 25 95 27 98
rect 37 75 39 78
rect 17 43 19 55
rect 13 41 21 43
rect 13 39 17 41
rect 19 39 21 41
rect 13 37 21 39
rect 25 41 27 55
rect 37 53 39 55
rect 31 51 39 53
rect 31 49 33 51
rect 35 49 39 51
rect 31 47 39 49
rect 41 41 47 43
rect 25 39 43 41
rect 45 39 47 41
rect 13 25 15 37
rect 25 25 27 39
rect 41 37 47 39
rect 31 31 39 33
rect 31 29 33 31
rect 35 29 39 31
rect 31 27 39 29
rect 37 25 39 27
rect 13 12 15 15
rect 25 12 27 15
rect 37 12 39 15
<< ndif >>
rect 5 15 13 25
rect 15 21 25 25
rect 15 19 19 21
rect 21 19 25 21
rect 15 15 25 19
rect 27 15 37 25
rect 39 21 47 25
rect 39 19 43 21
rect 45 19 47 21
rect 39 15 47 19
rect 5 11 11 15
rect 5 9 7 11
rect 9 9 11 11
rect 5 7 11 9
rect 29 11 35 15
rect 29 9 31 11
rect 33 9 35 11
rect 29 7 35 9
<< pdif >>
rect 13 85 17 95
rect 5 81 17 85
rect 5 79 7 81
rect 9 79 17 81
rect 5 71 17 79
rect 5 69 7 71
rect 9 69 17 71
rect 5 61 17 69
rect 5 59 7 61
rect 9 59 17 61
rect 5 55 17 59
rect 19 55 25 95
rect 27 91 35 95
rect 27 89 31 91
rect 33 89 35 91
rect 27 75 35 89
rect 27 55 37 75
rect 39 71 47 75
rect 39 69 43 71
rect 45 69 47 71
rect 39 61 47 69
rect 39 59 43 61
rect 45 59 47 61
rect 39 55 47 59
<< alu1 >>
rect -2 95 52 100
rect -2 93 43 95
rect 45 93 52 95
rect -2 91 52 93
rect -2 89 31 91
rect 33 89 52 91
rect -2 88 52 89
rect 6 81 12 82
rect 6 79 7 81
rect 9 79 12 81
rect 6 78 12 79
rect 8 72 12 78
rect 6 71 12 72
rect 6 69 7 71
rect 9 69 12 71
rect 6 68 12 69
rect 8 62 12 68
rect 6 61 12 62
rect 6 59 7 61
rect 9 59 12 61
rect 6 58 12 59
rect 8 52 12 58
rect 4 48 12 52
rect 4 32 8 48
rect 18 42 22 82
rect 16 41 22 42
rect 16 39 17 41
rect 19 39 22 41
rect 16 38 22 39
rect 4 28 12 32
rect 18 28 22 38
rect 28 52 32 82
rect 42 71 46 72
rect 42 69 43 71
rect 45 69 46 71
rect 42 68 46 69
rect 43 62 45 68
rect 42 61 46 62
rect 42 59 43 61
rect 45 59 46 61
rect 42 58 46 59
rect 28 51 36 52
rect 28 49 33 51
rect 35 49 36 51
rect 28 48 36 49
rect 28 32 32 48
rect 43 42 45 58
rect 42 41 46 42
rect 42 39 43 41
rect 45 39 46 41
rect 42 38 46 39
rect 28 31 36 32
rect 28 29 33 31
rect 35 29 36 31
rect 28 28 36 29
rect 8 22 12 28
rect 8 21 22 22
rect 8 19 19 21
rect 21 19 22 21
rect 8 18 22 19
rect 28 18 32 28
rect 43 22 45 38
rect 42 21 46 22
rect 42 19 43 21
rect 45 19 46 21
rect 42 18 46 19
rect -2 11 52 12
rect -2 9 7 11
rect 9 9 31 11
rect 33 9 52 11
rect -2 0 52 9
<< ntie >>
rect 41 95 47 97
rect 41 93 43 95
rect 45 93 47 95
rect 41 85 47 93
<< nmos >>
rect 13 15 15 25
rect 25 15 27 25
rect 37 15 39 25
<< pmos >>
rect 17 55 19 95
rect 25 55 27 95
rect 37 55 39 75
<< polyct1 >>
rect 17 39 19 41
rect 33 49 35 51
rect 43 39 45 41
rect 33 29 35 31
<< ndifct1 >>
rect 19 19 21 21
rect 43 19 45 21
rect 7 9 9 11
rect 31 9 33 11
<< ntiect1 >>
rect 43 93 45 95
<< pdifct1 >>
rect 7 79 9 81
rect 7 69 9 71
rect 7 59 9 61
rect 31 89 33 91
rect 43 69 45 71
rect 43 59 45 61
<< labels >>
rlabel alu1 10 25 10 25 6 q
rlabel alu1 20 55 20 55 6 i0
rlabel alu1 10 65 10 65 6 q
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 50 30 50 6 i1
rlabel alu1 25 94 25 94 6 vdd
<< end >>
