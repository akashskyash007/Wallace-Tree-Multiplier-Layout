magic
tech scmos
timestamp 1199202658
<< ab >>
rect 0 0 88 80
<< nwell >>
rect -5 36 93 88
<< pwell >>
rect -5 -8 93 36
<< poly >>
rect 9 66 11 71
rect 19 66 21 71
rect 29 66 31 71
rect 39 66 41 71
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 39 39 41 42
rect 39 37 47 39
rect 39 35 43 37
rect 45 35 47 37
rect 57 37 63 39
rect 57 35 59 37
rect 61 35 63 37
rect 72 37 79 39
rect 72 35 75 37
rect 77 35 79 37
rect 19 33 31 35
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 33 50 35
rect 36 30 38 33
rect 48 30 50 33
rect 55 33 67 35
rect 55 30 57 33
rect 65 30 67 33
rect 72 33 79 35
rect 72 30 74 33
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
rect 48 6 50 10
rect 55 6 57 10
rect 65 6 67 10
rect 72 6 74 10
<< ndif >>
rect 3 14 12 30
rect 3 12 6 14
rect 8 12 12 14
rect 3 10 12 12
rect 14 10 19 30
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 10 29 19
rect 31 10 36 30
rect 38 14 48 30
rect 38 12 42 14
rect 44 12 48 14
rect 38 10 48 12
rect 50 10 55 30
rect 57 21 65 30
rect 57 19 60 21
rect 62 19 65 21
rect 57 10 65 19
rect 67 10 72 30
rect 74 21 82 30
rect 74 19 77 21
rect 79 19 82 21
rect 74 14 82 19
rect 74 12 77 14
rect 79 12 82 14
rect 74 10 82 12
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 42 9 62
rect 11 60 19 66
rect 11 58 14 60
rect 16 58 19 60
rect 11 53 19 58
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 42 29 62
rect 31 61 39 66
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 56 49 62
rect 41 54 44 56
rect 46 54 49 56
rect 41 42 49 54
<< alu1 >>
rect -2 81 90 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 90 81
rect -2 68 90 79
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 2 53 38 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 51 38 53
rect 2 50 38 51
rect 2 22 6 50
rect 25 42 63 46
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 41 37 47 38
rect 41 35 43 37
rect 45 35 47 37
rect 41 30 47 35
rect 57 37 63 42
rect 57 35 59 37
rect 61 35 63 37
rect 57 34 63 35
rect 73 37 79 38
rect 73 35 75 37
rect 77 35 79 37
rect 73 30 79 35
rect 10 26 79 30
rect 2 21 64 22
rect 2 19 24 21
rect 26 19 60 21
rect 62 19 64 21
rect 2 18 64 19
rect -2 1 90 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 90 1
rect -2 -2 90 -1
<< ptie >>
rect 0 1 88 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 88 1
rect 0 -3 88 -1
<< ntie >>
rect 0 81 88 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 88 81
rect 0 77 88 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 48 10 50 30
rect 55 10 57 30
rect 65 10 67 30
rect 72 10 74 30
<< pmos >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 43 35 45 37
rect 59 35 61 37
rect 75 35 77 37
<< ndifct0 >>
rect 6 12 8 14
rect 42 12 44 14
rect 77 19 79 21
rect 77 12 79 14
<< ndifct1 >>
rect 24 19 26 21
rect 60 19 62 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
<< pdifct0 >>
rect 4 62 6 64
rect 14 58 16 60
rect 24 62 26 64
rect 44 62 46 64
rect 44 54 46 56
<< pdifct1 >>
rect 14 51 16 53
rect 34 59 36 61
rect 34 51 36 53
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 23 64 27 68
rect 23 62 24 64
rect 26 62 27 64
rect 43 64 47 68
rect 3 60 7 62
rect 13 60 17 62
rect 23 60 27 62
rect 13 58 14 60
rect 16 58 17 60
rect 13 54 17 58
rect 43 62 44 64
rect 46 62 47 64
rect 43 56 47 62
rect 43 54 44 56
rect 46 54 47 56
rect 43 52 47 54
rect 75 21 81 22
rect 75 19 77 21
rect 79 19 81 21
rect 4 14 10 15
rect 4 12 6 14
rect 8 12 10 14
rect 40 14 46 15
rect 40 12 42 14
rect 44 12 46 14
rect 75 14 81 19
rect 75 12 77 14
rect 79 12 81 14
<< labels >>
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel polyct1 28 36 28 36 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 44 6 44 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 20 44 20 6 z
rlabel alu1 44 32 44 32 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 60 36 60 6 z
rlabel alu1 44 74 44 74 6 vdd
rlabel alu1 52 20 52 20 6 z
rlabel alu1 52 28 52 28 6 a
rlabel alu1 60 20 60 20 6 z
rlabel alu1 60 28 60 28 6 a
rlabel alu1 68 28 68 28 6 a
rlabel alu1 52 44 52 44 6 b
rlabel polyct1 60 36 60 36 6 b
rlabel alu1 60 40 60 40 6 b
rlabel alu1 76 32 76 32 6 a
<< end >>
