magic
tech scmos
timestamp 1199202154
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 12 69 14 74
rect 22 69 24 74
rect 29 69 31 74
rect 39 69 41 74
rect 49 69 51 74
rect 61 69 63 74
rect 12 39 14 42
rect 22 39 24 42
rect 9 37 24 39
rect 9 35 11 37
rect 13 35 24 37
rect 29 36 31 42
rect 39 39 41 42
rect 49 39 51 42
rect 61 39 63 42
rect 9 33 24 35
rect 28 33 31 36
rect 37 37 43 39
rect 37 35 39 37
rect 41 35 43 37
rect 37 33 43 35
rect 47 37 53 39
rect 47 35 49 37
rect 51 35 53 37
rect 47 33 53 35
rect 57 37 63 39
rect 57 35 59 37
rect 61 35 63 37
rect 57 33 63 35
rect 9 28 11 33
rect 21 30 23 33
rect 28 30 30 33
rect 38 30 40 33
rect 48 30 50 33
rect 59 30 61 33
rect 9 11 11 16
rect 21 13 23 18
rect 28 9 30 18
rect 38 13 40 18
rect 48 9 50 18
rect 59 13 61 18
rect 28 7 50 9
<< ndif >>
rect 13 28 21 30
rect 4 22 9 28
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 18 21 28
rect 23 18 28 30
rect 30 28 38 30
rect 30 26 33 28
rect 35 26 38 28
rect 30 18 38 26
rect 40 22 48 30
rect 40 20 43 22
rect 45 20 48 22
rect 40 18 48 20
rect 50 22 59 30
rect 50 20 53 22
rect 55 20 59 22
rect 50 18 59 20
rect 61 28 68 30
rect 61 26 64 28
rect 66 26 68 28
rect 61 24 68 26
rect 61 18 66 24
rect 11 16 19 18
rect 13 11 19 16
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
<< pdif >>
rect 7 63 12 69
rect 5 61 12 63
rect 5 59 7 61
rect 9 59 12 61
rect 5 54 12 59
rect 5 52 7 54
rect 9 52 12 54
rect 5 50 12 52
rect 7 42 12 50
rect 14 67 22 69
rect 14 65 17 67
rect 19 65 22 67
rect 14 60 22 65
rect 14 58 17 60
rect 19 58 22 60
rect 14 42 22 58
rect 24 42 29 69
rect 31 53 39 69
rect 31 51 34 53
rect 36 51 39 53
rect 31 46 39 51
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 62 49 69
rect 41 60 44 62
rect 46 60 49 62
rect 41 42 49 60
rect 51 67 61 69
rect 51 65 55 67
rect 57 65 61 67
rect 51 42 61 65
rect 63 55 68 69
rect 63 53 70 55
rect 63 51 66 53
rect 68 51 70 53
rect 63 46 70 51
rect 63 44 66 46
rect 68 44 70 46
rect 63 42 70 44
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 33 53 38 55
rect 33 51 34 53
rect 36 51 38 53
rect 2 39 6 47
rect 33 46 38 51
rect 18 44 34 46
rect 36 44 38 46
rect 18 42 38 44
rect 42 45 46 55
rect 50 49 62 55
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 18 30 22 42
rect 42 41 54 45
rect 48 37 54 41
rect 48 35 49 37
rect 51 35 54 37
rect 48 33 54 35
rect 58 37 62 49
rect 58 35 59 37
rect 61 35 62 37
rect 58 33 62 35
rect 18 28 37 30
rect 18 26 33 28
rect 35 26 37 28
rect 18 25 37 26
rect -2 11 74 12
rect -2 9 15 11
rect 17 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 9 16 11 28
rect 21 18 23 30
rect 28 18 30 30
rect 38 18 40 30
rect 48 18 50 30
rect 59 18 61 30
<< pmos >>
rect 12 42 14 69
rect 22 42 24 69
rect 29 42 31 69
rect 39 42 41 69
rect 49 42 51 69
rect 61 42 63 69
<< polyct0 >>
rect 39 35 41 37
<< polyct1 >>
rect 11 35 13 37
rect 49 35 51 37
rect 59 35 61 37
<< ndifct0 >>
rect 4 18 6 20
rect 43 20 45 22
rect 53 20 55 22
rect 64 26 66 28
<< ndifct1 >>
rect 33 26 35 28
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 7 59 9 61
rect 7 52 9 54
rect 17 65 19 67
rect 17 58 19 60
rect 44 60 46 62
rect 55 65 57 67
rect 66 51 68 53
rect 66 44 68 46
<< pdifct1 >>
rect 34 51 36 53
rect 34 44 36 46
<< alu0 >>
rect 15 67 21 68
rect 15 65 17 67
rect 19 65 21 67
rect 6 61 10 63
rect 6 59 7 61
rect 9 59 10 61
rect 6 54 10 59
rect 15 60 21 65
rect 54 67 58 68
rect 54 65 55 67
rect 57 65 58 67
rect 54 63 58 65
rect 15 58 17 60
rect 19 58 21 60
rect 15 57 21 58
rect 24 62 48 63
rect 24 60 44 62
rect 46 60 48 62
rect 24 59 48 60
rect 24 54 28 59
rect 6 52 7 54
rect 9 52 28 54
rect 6 50 28 52
rect 37 37 45 38
rect 37 35 39 37
rect 41 35 45 37
rect 37 34 45 35
rect 41 30 45 34
rect 65 53 70 55
rect 65 51 66 53
rect 68 51 70 53
rect 65 46 70 51
rect 65 44 66 46
rect 68 44 70 46
rect 65 42 70 44
rect 66 30 70 42
rect 41 28 70 30
rect 41 26 64 28
rect 66 26 70 28
rect 62 25 70 26
rect 41 22 47 23
rect 41 21 43 22
rect 2 20 43 21
rect 45 20 47 22
rect 2 18 4 20
rect 6 18 47 20
rect 2 17 47 18
rect 51 22 57 23
rect 51 20 53 22
rect 55 20 57 22
rect 51 12 57 20
<< labels >>
rlabel alu0 8 56 8 56 6 n1
rlabel alu0 24 19 24 19 6 n3
rlabel alu0 36 61 36 61 6 n1
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 4 40 4 40 6 a
rlabel alu1 20 32 20 32 6 z
rlabel alu1 28 28 28 28 6 z
rlabel alu1 28 44 28 44 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 52 36 52 36 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 52 52 52 52 6 c
rlabel alu1 44 48 44 48 6 b
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 44 60 44 6 c
<< end >>
