magic
tech scmos
timestamp 1199202394
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 22 39
rect 9 35 18 37
rect 20 35 22 37
rect 9 33 22 35
rect 10 30 12 33
rect 20 30 22 33
rect 10 15 12 19
rect 20 15 22 19
<< ndif >>
rect 2 21 10 30
rect 2 19 4 21
rect 6 19 10 21
rect 12 28 20 30
rect 12 26 15 28
rect 17 26 20 28
rect 12 19 20 26
rect 22 24 29 30
rect 22 22 25 24
rect 27 22 29 24
rect 22 19 29 22
rect 2 17 8 19
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 68 28 70
rect 21 66 24 68
rect 26 66 28 68
rect 21 61 28 66
rect 21 59 24 61
rect 26 59 28 61
rect 21 42 28 59
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 52 14 54
rect 16 52 23 54
rect 2 50 23 52
rect 2 29 6 50
rect 17 39 23 46
rect 17 37 30 39
rect 17 35 18 37
rect 20 35 30 37
rect 17 33 30 35
rect 2 28 19 29
rect 2 26 15 28
rect 17 26 19 28
rect 2 25 19 26
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 10 19 12 30
rect 20 19 22 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
<< polyct1 >>
rect 18 35 20 37
<< ndifct0 >>
rect 4 19 6 21
rect 25 22 27 24
<< ndifct1 >>
rect 15 26 17 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 14 59 16 61
rect 24 66 26 68
rect 24 59 26 61
<< pdifct1 >>
rect 14 52 16 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 22 66 24 68
rect 26 66 28 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 61 28 66
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 24 24 28 26
rect 24 22 25 24
rect 27 22 28 24
rect 2 21 8 22
rect 2 19 4 21
rect 6 19 8 21
rect 2 12 8 19
rect 24 12 28 22
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 20 40 20 40 6 a
rlabel alu1 20 52 20 52 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 28 36 28 36 6 a
<< end >>
