magic
tech scmos
timestamp 1199203197
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 39 65 41 70
rect 46 65 48 70
rect 29 58 31 63
rect 9 50 11 55
rect 29 43 31 50
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 9 35 11 38
rect 29 37 35 39
rect 9 33 18 35
rect 9 31 14 33
rect 16 31 18 33
rect 9 29 18 31
rect 9 26 11 29
rect 29 26 31 37
rect 39 35 41 50
rect 46 43 48 50
rect 46 41 57 43
rect 51 39 53 41
rect 55 39 57 41
rect 51 37 57 39
rect 39 33 47 35
rect 39 31 43 33
rect 45 31 47 33
rect 39 29 47 31
rect 39 26 41 29
rect 9 15 11 20
rect 51 19 53 37
rect 29 14 31 19
rect 39 14 41 19
rect 51 7 53 12
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 11 24 18 26
rect 11 22 14 24
rect 16 22 18 24
rect 11 20 18 22
rect 22 24 29 26
rect 22 22 24 24
rect 26 22 29 24
rect 22 19 29 22
rect 31 23 39 26
rect 31 21 34 23
rect 36 21 39 23
rect 31 19 39 21
rect 41 19 49 26
rect 43 12 51 19
rect 53 16 60 19
rect 53 14 56 16
rect 58 14 60 16
rect 53 12 60 14
rect 43 7 49 12
rect 43 5 45 7
rect 47 5 49 7
rect 43 3 49 5
<< pdif >>
rect 13 58 27 60
rect 34 58 39 65
rect 13 56 15 58
rect 17 56 29 58
rect 13 50 29 56
rect 31 56 39 58
rect 31 54 34 56
rect 36 54 39 56
rect 31 50 39 54
rect 41 50 46 65
rect 48 63 56 65
rect 48 61 51 63
rect 53 61 56 63
rect 48 56 56 61
rect 48 54 51 56
rect 53 54 56 56
rect 48 50 56 54
rect 4 44 9 50
rect 2 42 9 44
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 48 15 50
rect 17 48 27 50
rect 11 38 27 48
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 66 67
rect -2 64 66 65
rect 2 42 15 43
rect 2 40 4 42
rect 6 40 15 42
rect 2 38 15 40
rect 2 26 6 38
rect 42 46 46 51
rect 34 43 46 46
rect 30 42 46 43
rect 30 41 38 42
rect 30 39 31 41
rect 33 39 38 41
rect 30 37 38 39
rect 50 41 62 43
rect 50 39 53 41
rect 55 39 62 41
rect 50 37 62 39
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 20 7 22
rect 2 13 6 20
rect 42 33 46 35
rect 42 31 43 33
rect 45 31 46 33
rect 42 27 46 31
rect 58 29 62 37
rect 42 21 54 27
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 13 7
rect 15 5 45 7
rect 47 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 17 9
rect 3 5 5 7
rect 7 5 13 7
rect 15 5 17 7
rect 3 3 17 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 57 9 65
<< nmos >>
rect 9 20 11 26
rect 29 19 31 26
rect 39 19 41 26
rect 51 12 53 19
<< pmos >>
rect 29 50 31 58
rect 39 50 41 65
rect 46 50 48 65
rect 9 38 11 50
<< polyct0 >>
rect 14 31 16 33
<< polyct1 >>
rect 31 39 33 41
rect 53 39 55 41
rect 43 31 45 33
<< ndifct0 >>
rect 14 22 16 24
rect 24 22 26 24
rect 34 21 36 23
rect 56 14 58 16
<< ndifct1 >>
rect 4 22 6 24
rect 45 5 47 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
rect 13 5 15 7
<< pdifct0 >>
rect 15 56 17 58
rect 34 54 36 56
rect 51 61 53 63
rect 51 54 53 56
rect 15 48 17 50
<< pdifct1 >>
rect 4 40 6 42
<< alu0 >>
rect 13 58 19 64
rect 13 56 15 58
rect 17 56 19 58
rect 50 63 54 64
rect 50 61 51 63
rect 53 61 54 63
rect 13 50 19 56
rect 13 48 15 50
rect 17 48 19 50
rect 13 47 19 48
rect 23 56 38 57
rect 23 54 34 56
rect 36 54 38 56
rect 23 53 38 54
rect 50 56 54 61
rect 50 54 51 56
rect 53 54 54 56
rect 23 34 27 53
rect 50 52 54 54
rect 12 33 27 34
rect 12 31 14 33
rect 16 31 27 33
rect 12 30 27 31
rect 13 24 17 26
rect 13 22 14 24
rect 16 22 17 24
rect 13 8 17 22
rect 23 24 27 30
rect 23 22 24 24
rect 26 22 27 24
rect 23 20 27 22
rect 33 23 37 25
rect 33 21 34 23
rect 36 21 37 23
rect 33 17 37 21
rect 33 16 60 17
rect 33 14 56 16
rect 58 14 60 16
rect 33 13 60 14
<< labels >>
rlabel alu0 35 19 35 19 6 n1
rlabel alu0 19 32 19 32 6 zn
rlabel alu0 25 38 25 38 6 zn
rlabel alu0 30 55 30 55 6 zn
rlabel alu0 46 15 46 15 6 n1
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 36 40 36 40 6 b
rlabel alu1 44 48 44 48 6 b
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 24 52 24 6 a2
rlabel alu1 60 36 60 36 6 a1
rlabel alu1 52 40 52 40 6 a1
<< end >>
