magic
tech scmos
timestamp 1199202161
<< ab >>
rect 0 0 128 80
<< nwell >>
rect -5 36 133 88
<< pwell >>
rect -5 -8 133 36
<< poly >>
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 71 70 73 74
rect 78 70 80 74
rect 88 70 90 74
rect 95 70 97 74
rect 107 70 109 74
rect 117 70 119 74
rect 9 58 11 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 21 39
rect 9 35 11 37
rect 13 35 21 37
rect 9 33 21 35
rect 25 37 31 39
rect 25 35 27 37
rect 29 35 31 37
rect 25 33 31 35
rect 9 30 11 33
rect 19 27 21 33
rect 29 30 31 33
rect 39 39 41 42
rect 49 39 51 42
rect 39 37 51 39
rect 39 35 41 37
rect 43 35 51 37
rect 39 33 51 35
rect 39 30 41 33
rect 49 30 51 33
rect 59 39 61 42
rect 71 39 73 42
rect 59 37 73 39
rect 59 35 63 37
rect 65 35 73 37
rect 59 33 73 35
rect 59 30 61 33
rect 71 30 73 33
rect 78 39 80 42
rect 88 39 90 42
rect 78 37 90 39
rect 78 35 86 37
rect 88 35 90 37
rect 78 33 90 35
rect 78 30 80 33
rect 88 30 90 33
rect 95 39 97 42
rect 107 39 109 42
rect 117 39 119 42
rect 95 37 103 39
rect 95 35 99 37
rect 101 35 103 37
rect 95 33 103 35
rect 107 37 119 39
rect 107 35 115 37
rect 117 35 119 37
rect 107 33 119 35
rect 95 30 97 33
rect 107 30 109 33
rect 117 30 119 33
rect 9 15 11 19
rect 19 11 21 16
rect 29 11 31 16
rect 39 11 41 16
rect 49 11 51 16
rect 59 11 61 16
rect 88 15 90 19
rect 95 15 97 19
rect 71 8 73 13
rect 78 8 80 13
rect 107 11 109 16
rect 117 11 119 16
<< ndif >>
rect 2 23 9 30
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 27 16 30
rect 23 27 29 30
rect 11 25 19 27
rect 11 23 14 25
rect 16 23 19 25
rect 11 19 19 23
rect 14 16 19 19
rect 21 20 29 27
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 31 20 39 30
rect 31 18 34 20
rect 36 18 39 20
rect 31 16 39 18
rect 41 28 49 30
rect 41 26 44 28
rect 46 26 49 28
rect 41 16 49 26
rect 51 20 59 30
rect 51 18 54 20
rect 56 18 59 20
rect 51 16 59 18
rect 61 16 71 30
rect 63 13 71 16
rect 73 13 78 30
rect 80 28 88 30
rect 80 26 83 28
rect 85 26 88 28
rect 80 19 88 26
rect 90 19 95 30
rect 97 19 107 30
rect 80 13 85 19
rect 99 16 107 19
rect 109 20 117 30
rect 109 18 112 20
rect 114 18 117 20
rect 109 16 117 18
rect 119 27 126 30
rect 119 25 122 27
rect 124 25 126 27
rect 119 20 126 25
rect 119 18 122 20
rect 124 18 126 20
rect 119 16 126 18
rect 63 11 69 13
rect 63 9 65 11
rect 67 9 69 11
rect 63 7 69 9
rect 99 11 105 16
rect 99 9 101 11
rect 103 9 105 11
rect 99 7 105 9
<< pdif >>
rect 14 58 19 70
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 42 9 54
rect 11 53 19 58
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 42 39 59
rect 41 46 49 70
rect 41 44 44 46
rect 46 44 49 46
rect 41 42 49 44
rect 51 61 59 70
rect 51 59 54 61
rect 56 59 59 61
rect 51 42 59 59
rect 61 68 71 70
rect 61 66 65 68
rect 67 66 71 68
rect 61 42 71 66
rect 73 42 78 70
rect 80 46 88 70
rect 80 44 83 46
rect 85 44 88 46
rect 80 42 88 44
rect 90 42 95 70
rect 97 68 107 70
rect 97 66 101 68
rect 103 66 107 68
rect 97 42 107 66
rect 109 61 117 70
rect 109 59 112 61
rect 114 59 117 61
rect 109 54 117 59
rect 109 52 112 54
rect 114 52 117 54
rect 109 42 117 52
rect 119 68 126 70
rect 119 66 122 68
rect 124 66 126 68
rect 119 60 126 66
rect 119 58 122 60
rect 124 58 126 60
rect 119 42 126 58
<< alu1 >>
rect -2 81 130 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 130 81
rect -2 68 130 79
rect 2 39 6 47
rect 26 50 103 54
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 26 37 30 50
rect 41 44 44 46
rect 46 44 55 46
rect 41 42 55 44
rect 26 35 27 37
rect 29 35 30 37
rect 26 33 30 35
rect 50 30 55 42
rect 73 44 83 46
rect 85 44 87 46
rect 73 42 87 44
rect 97 42 103 50
rect 73 30 78 42
rect 84 37 95 38
rect 84 35 86 37
rect 88 35 95 37
rect 84 34 95 35
rect 89 30 95 34
rect 114 37 118 39
rect 114 35 115 37
rect 117 35 118 37
rect 114 30 118 35
rect 41 28 78 30
rect 41 26 44 28
rect 46 26 78 28
rect 89 26 118 30
rect -2 11 130 12
rect -2 9 65 11
rect 67 9 101 11
rect 103 9 130 11
rect -2 1 130 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 130 1
rect -2 -2 130 -1
<< ptie >>
rect 0 1 128 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 128 1
rect 0 -3 128 -1
<< ntie >>
rect 0 81 128 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 128 81
rect 0 77 128 79
<< nmos >>
rect 9 19 11 30
rect 19 16 21 27
rect 29 16 31 30
rect 39 16 41 30
rect 49 16 51 30
rect 59 16 61 30
rect 71 13 73 30
rect 78 13 80 30
rect 88 19 90 30
rect 95 19 97 30
rect 107 16 109 30
rect 117 16 119 30
<< pmos >>
rect 9 42 11 58
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 71 42 73 70
rect 78 42 80 70
rect 88 42 90 70
rect 95 42 97 70
rect 107 42 109 70
rect 117 42 119 70
<< polyct0 >>
rect 41 35 43 37
rect 63 35 65 37
rect 99 35 101 37
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 86 35 88 37
rect 115 35 117 37
<< ndifct0 >>
rect 4 21 6 23
rect 14 23 16 25
rect 24 18 26 20
rect 34 18 36 20
rect 54 18 56 20
rect 83 26 85 28
rect 112 18 114 20
rect 122 25 124 27
rect 122 18 124 20
<< ndifct1 >>
rect 44 26 46 28
rect 65 9 67 11
rect 101 9 103 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
<< pdifct0 >>
rect 4 54 6 56
rect 14 51 16 53
rect 14 44 16 46
rect 24 66 26 68
rect 24 59 26 61
rect 34 59 36 61
rect 54 59 56 61
rect 65 66 67 68
rect 101 66 103 68
rect 112 59 114 61
rect 112 52 114 54
rect 122 66 124 68
rect 122 58 124 60
<< pdifct1 >>
rect 44 44 46 46
rect 83 44 85 46
<< alu0 >>
rect 3 56 7 68
rect 23 66 24 68
rect 26 66 27 68
rect 23 61 27 66
rect 63 66 65 68
rect 67 66 69 68
rect 63 65 69 66
rect 99 66 101 68
rect 103 66 105 68
rect 99 65 105 66
rect 121 66 122 68
rect 124 66 125 68
rect 23 59 24 61
rect 26 59 27 61
rect 23 57 27 59
rect 32 61 116 62
rect 32 59 34 61
rect 36 59 54 61
rect 56 59 112 61
rect 114 59 116 61
rect 32 58 116 59
rect 3 54 4 56
rect 6 54 7 56
rect 3 52 7 54
rect 13 53 17 55
rect 111 54 116 58
rect 121 60 125 66
rect 121 58 122 60
rect 124 58 125 60
rect 121 56 125 58
rect 13 51 14 53
rect 16 51 17 53
rect 13 46 17 51
rect 111 52 112 54
rect 114 52 116 54
rect 111 50 116 52
rect 13 44 14 46
rect 16 44 22 46
rect 13 42 22 44
rect 18 29 22 42
rect 42 46 48 47
rect 34 37 45 38
rect 34 35 41 37
rect 43 35 45 37
rect 34 34 45 35
rect 34 29 38 34
rect 62 37 66 50
rect 81 46 87 47
rect 62 35 63 37
rect 65 35 66 37
rect 62 33 66 35
rect 98 37 102 42
rect 98 35 99 37
rect 101 35 102 37
rect 98 33 102 35
rect 13 25 38 29
rect 78 28 86 30
rect 78 26 83 28
rect 85 26 86 28
rect 121 27 125 29
rect 42 25 48 26
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 13 23 14 25
rect 16 23 17 25
rect 73 24 86 26
rect 121 25 122 27
rect 124 25 125 27
rect 13 21 17 23
rect 3 12 7 21
rect 23 20 27 22
rect 23 18 24 20
rect 26 18 27 20
rect 23 12 27 18
rect 32 20 116 21
rect 32 18 34 20
rect 36 18 54 20
rect 56 18 112 20
rect 114 18 116 20
rect 32 17 116 18
rect 121 20 125 25
rect 121 18 122 20
rect 124 18 125 20
rect 121 12 125 18
<< labels >>
rlabel alu0 15 48 15 48 6 cn
rlabel alu0 39 36 39 36 6 cn
rlabel alu0 25 27 25 27 6 cn
rlabel alu0 74 19 74 19 6 n3
rlabel alu0 113 56 113 56 6 n1
rlabel alu0 74 60 74 60 6 n1
rlabel alu1 4 40 4 40 6 c
rlabel polyct1 12 36 12 36 6 c
rlabel alu1 44 28 44 28 6 z
rlabel alu1 28 40 28 40 6 a
rlabel alu1 44 44 44 44 6 z
rlabel alu1 36 52 36 52 6 a
rlabel alu1 44 52 44 52 6 a
rlabel alu1 64 6 64 6 6 vss
rlabel alu1 60 28 60 28 6 z
rlabel alu1 68 28 68 28 6 z
rlabel alu1 52 36 52 36 6 z
rlabel alu1 60 52 60 52 6 a
rlabel alu1 68 52 68 52 6 a
rlabel alu1 52 52 52 52 6 a
rlabel alu1 64 74 64 74 6 vdd
rlabel alu1 100 28 100 28 6 b
rlabel alu1 92 32 92 32 6 b
rlabel alu1 76 36 76 36 6 z
rlabel alu1 84 44 84 44 6 z
rlabel alu1 100 48 100 48 6 a
rlabel alu1 84 52 84 52 6 a
rlabel alu1 92 52 92 52 6 a
rlabel alu1 76 52 76 52 6 a
rlabel alu1 108 28 108 28 6 b
rlabel polyct1 116 36 116 36 6 b
<< end >>
