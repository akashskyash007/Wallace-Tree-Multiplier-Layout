magic
tech scmos
timestamp 1199543171
<< ab >>
rect 0 0 130 100
<< nwell >>
rect -5 48 135 105
<< pwell >>
rect -5 -5 135 48
<< poly >>
rect 23 94 25 98
rect 35 94 37 98
rect 11 79 13 83
rect 47 85 49 89
rect 59 85 61 89
rect 71 85 73 89
rect 83 85 85 89
rect 97 85 99 89
rect 107 85 109 89
rect 117 85 119 89
rect 11 43 13 55
rect 23 53 25 56
rect 35 53 37 56
rect 17 51 37 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 47 43 49 63
rect 59 43 61 63
rect 71 43 73 63
rect 83 43 85 61
rect 11 41 43 43
rect 11 29 13 41
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 67 41 73 43
rect 67 39 69 41
rect 71 39 73 41
rect 67 37 73 39
rect 77 41 85 43
rect 77 39 79 41
rect 81 39 85 41
rect 97 53 99 56
rect 107 53 109 56
rect 97 51 103 53
rect 97 49 99 51
rect 101 49 103 51
rect 97 47 103 49
rect 107 51 113 53
rect 107 49 109 51
rect 111 49 113 51
rect 107 47 113 49
rect 97 39 99 47
rect 107 39 109 47
rect 77 37 85 39
rect 93 37 99 39
rect 105 37 109 39
rect 117 43 119 55
rect 117 41 123 43
rect 117 39 119 41
rect 121 39 123 41
rect 117 37 123 39
rect 17 35 23 37
rect 17 33 19 35
rect 21 33 23 35
rect 49 33 51 37
rect 59 33 61 37
rect 69 33 71 37
rect 17 31 37 33
rect 23 28 25 31
rect 35 28 37 31
rect 11 11 13 15
rect 81 29 83 37
rect 93 25 95 37
rect 105 25 107 37
rect 117 25 119 37
rect 49 13 51 17
rect 59 13 61 17
rect 69 13 71 17
rect 81 13 83 17
rect 93 13 95 17
rect 105 13 107 17
rect 117 13 119 17
rect 23 4 25 8
rect 35 4 37 8
<< ndif >>
rect 3 25 11 29
rect 3 23 5 25
rect 7 23 11 25
rect 3 15 11 23
rect 13 28 18 29
rect 41 28 49 33
rect 13 25 23 28
rect 13 23 17 25
rect 19 23 23 25
rect 13 15 23 23
rect 15 13 17 15
rect 19 13 23 15
rect 15 8 23 13
rect 25 21 35 28
rect 25 19 29 21
rect 31 19 35 21
rect 25 8 35 19
rect 37 17 49 28
rect 51 17 59 33
rect 61 17 69 33
rect 71 29 76 33
rect 71 21 81 29
rect 71 19 75 21
rect 77 19 81 21
rect 71 17 81 19
rect 83 25 90 29
rect 83 21 93 25
rect 83 19 87 21
rect 89 19 93 21
rect 83 17 93 19
rect 95 17 105 25
rect 107 21 117 25
rect 107 19 111 21
rect 113 19 117 21
rect 107 17 117 19
rect 119 21 127 25
rect 119 19 123 21
rect 125 19 127 21
rect 119 17 127 19
rect 37 11 47 17
rect 97 11 103 17
rect 37 9 43 11
rect 45 9 47 11
rect 37 8 47 9
rect 41 7 47 8
rect 97 9 99 11
rect 101 9 103 11
rect 97 7 103 9
<< pdif >>
rect 15 91 23 94
rect 15 89 17 91
rect 19 89 23 91
rect 15 81 23 89
rect 15 79 17 81
rect 19 79 23 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 71 23 79
rect 13 69 17 71
rect 19 69 23 71
rect 13 61 23 69
rect 13 59 17 61
rect 19 59 23 61
rect 13 56 23 59
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 56 35 59
rect 37 85 44 94
rect 63 91 69 93
rect 63 89 65 91
rect 67 89 69 91
rect 63 85 69 89
rect 37 81 47 85
rect 37 79 41 81
rect 43 79 47 81
rect 37 63 47 79
rect 49 81 59 85
rect 49 79 53 81
rect 55 79 59 81
rect 49 63 59 79
rect 61 63 71 85
rect 73 81 83 85
rect 73 79 77 81
rect 79 79 83 81
rect 73 63 83 79
rect 37 56 44 63
rect 13 55 18 56
rect 76 61 83 63
rect 85 71 97 85
rect 85 69 89 71
rect 91 69 97 71
rect 85 61 97 69
rect 87 59 89 61
rect 91 59 97 61
rect 87 56 97 59
rect 99 56 107 85
rect 109 56 117 85
rect 112 55 117 56
rect 119 81 127 85
rect 119 79 123 81
rect 125 79 127 81
rect 119 55 127 79
<< alu1 >>
rect -2 95 132 100
rect -2 93 5 95
rect 7 93 77 95
rect 79 93 89 95
rect 91 93 101 95
rect 103 93 113 95
rect 115 93 132 95
rect -2 91 132 93
rect -2 89 17 91
rect 19 89 65 91
rect 67 89 132 91
rect -2 88 132 89
rect 16 81 20 88
rect 16 79 17 81
rect 19 79 20 81
rect 4 71 8 73
rect 4 69 5 71
rect 7 69 8 71
rect 4 61 8 69
rect 4 59 5 61
rect 7 59 8 61
rect 4 52 8 59
rect 16 71 20 79
rect 16 69 17 71
rect 19 69 20 71
rect 16 61 20 69
rect 16 59 17 61
rect 19 59 20 61
rect 16 57 20 59
rect 28 81 32 83
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 40 81 44 88
rect 40 79 41 81
rect 43 79 44 81
rect 40 77 44 79
rect 51 81 127 82
rect 51 79 53 81
rect 55 79 77 81
rect 79 79 123 81
rect 125 79 127 81
rect 51 78 127 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 4 51 23 52
rect 4 49 19 51
rect 21 49 23 51
rect 4 48 23 49
rect 4 36 8 48
rect 4 35 23 36
rect 4 33 19 35
rect 21 33 23 35
rect 4 32 23 33
rect 4 25 8 32
rect 4 23 5 25
rect 7 23 8 25
rect 4 21 8 23
rect 16 25 20 27
rect 16 23 17 25
rect 19 23 20 25
rect 16 15 20 23
rect 28 21 32 59
rect 28 19 29 21
rect 31 19 32 21
rect 28 17 32 19
rect 38 41 42 43
rect 38 39 39 41
rect 41 39 42 41
rect 38 22 42 39
rect 48 41 52 73
rect 48 39 49 41
rect 51 39 52 41
rect 48 27 52 39
rect 58 41 62 73
rect 58 39 59 41
rect 61 39 62 41
rect 58 27 62 39
rect 68 41 72 73
rect 68 39 69 41
rect 71 39 72 41
rect 68 37 72 39
rect 78 41 82 73
rect 78 39 79 41
rect 81 39 82 41
rect 78 37 82 39
rect 88 71 92 73
rect 88 69 89 71
rect 91 69 92 71
rect 88 61 92 69
rect 88 59 89 61
rect 91 59 92 61
rect 88 32 92 59
rect 74 28 92 32
rect 98 51 102 73
rect 98 49 99 51
rect 101 49 102 51
rect 74 22 78 28
rect 98 27 102 49
rect 108 51 112 73
rect 108 49 109 51
rect 111 49 112 51
rect 108 27 112 49
rect 118 41 122 73
rect 118 39 119 41
rect 121 39 122 41
rect 118 27 122 39
rect 38 21 78 22
rect 38 19 75 21
rect 77 19 78 21
rect 38 18 78 19
rect 85 21 115 22
rect 85 19 87 21
rect 89 19 111 21
rect 113 19 115 21
rect 85 18 115 19
rect 122 21 126 23
rect 122 19 123 21
rect 125 19 126 21
rect 74 17 78 18
rect 16 13 17 15
rect 19 13 20 15
rect 16 12 20 13
rect 122 12 126 19
rect -2 11 132 12
rect -2 9 43 11
rect 45 9 99 11
rect 101 9 132 11
rect -2 7 55 9
rect 57 7 65 9
rect 67 7 75 9
rect 77 7 86 9
rect 88 7 113 9
rect 115 7 121 9
rect 123 7 132 9
rect -2 0 132 7
<< ptie >>
rect 53 9 90 11
rect 53 7 55 9
rect 57 7 65 9
rect 67 7 75 9
rect 77 7 86 9
rect 88 7 90 9
rect 111 9 125 11
rect 111 7 113 9
rect 115 7 121 9
rect 123 7 125 9
rect 53 5 90 7
rect 111 5 125 7
<< ntie >>
rect 3 95 9 97
rect 3 93 5 95
rect 7 93 9 95
rect 75 95 117 97
rect 3 86 9 93
rect 75 93 77 95
rect 79 93 89 95
rect 91 93 101 95
rect 103 93 113 95
rect 115 93 117 95
rect 75 91 117 93
<< nmos >>
rect 11 15 13 29
rect 23 8 25 28
rect 35 8 37 28
rect 49 17 51 33
rect 59 17 61 33
rect 69 17 71 33
rect 81 17 83 29
rect 93 17 95 25
rect 105 17 107 25
rect 117 17 119 25
<< pmos >>
rect 11 55 13 79
rect 23 56 25 94
rect 35 56 37 94
rect 47 63 49 85
rect 59 63 61 85
rect 71 63 73 85
rect 83 61 85 85
rect 97 56 99 85
rect 107 56 109 85
rect 117 55 119 85
<< polyct1 >>
rect 19 49 21 51
rect 39 39 41 41
rect 49 39 51 41
rect 59 39 61 41
rect 69 39 71 41
rect 79 39 81 41
rect 99 49 101 51
rect 109 49 111 51
rect 119 39 121 41
rect 19 33 21 35
<< ndifct1 >>
rect 5 23 7 25
rect 17 23 19 25
rect 17 13 19 15
rect 29 19 31 21
rect 75 19 77 21
rect 87 19 89 21
rect 111 19 113 21
rect 123 19 125 21
rect 43 9 45 11
rect 99 9 101 11
<< ntiect1 >>
rect 5 93 7 95
rect 77 93 79 95
rect 89 93 91 95
rect 101 93 103 95
rect 113 93 115 95
<< ptiect1 >>
rect 55 7 57 9
rect 65 7 67 9
rect 75 7 77 9
rect 86 7 88 9
rect 113 7 115 9
rect 121 7 123 9
<< pdifct1 >>
rect 17 89 19 91
rect 17 79 19 81
rect 5 69 7 71
rect 5 59 7 61
rect 17 69 19 71
rect 17 59 19 61
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
rect 65 89 67 91
rect 41 79 43 81
rect 53 79 55 81
rect 77 79 79 81
rect 89 69 91 71
rect 89 59 91 61
rect 123 79 125 81
<< labels >>
rlabel alu1 50 50 50 50 6 i0
rlabel alu1 60 50 60 50 6 i1
rlabel alu1 30 50 30 50 6 nq
rlabel alu1 65 6 65 6 6 vss
rlabel alu1 80 55 80 55 6 i6
rlabel alu1 70 55 70 55 6 i2
rlabel alu1 65 94 65 94 6 vdd
rlabel polyct1 110 50 110 50 6 i4
rlabel alu1 120 50 120 50 6 i5
rlabel polyct1 100 50 100 50 6 i3
<< end >>
