magic
tech scmos
timestamp 1199201937
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 31 70 33 74
rect 41 70 43 74
rect 31 47 33 50
rect 41 47 43 50
rect 31 45 37 47
rect 9 39 11 45
rect 19 39 21 45
rect 31 43 33 45
rect 35 43 37 45
rect 31 41 37 43
rect 41 45 47 47
rect 41 43 43 45
rect 45 43 47 45
rect 41 41 47 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 13 30 15 33
rect 20 30 22 33
rect 32 30 34 41
rect 41 36 43 41
rect 39 33 43 36
rect 39 30 41 33
rect 13 6 15 10
rect 20 6 22 10
rect 32 8 34 13
rect 39 8 41 13
<< ndif >>
rect 8 22 13 30
rect 6 20 13 22
rect 6 18 8 20
rect 10 18 13 20
rect 6 16 13 18
rect 8 10 13 16
rect 15 10 20 30
rect 22 13 32 30
rect 34 13 39 30
rect 41 22 46 30
rect 41 20 48 22
rect 41 18 44 20
rect 46 18 48 20
rect 41 16 48 18
rect 41 13 46 16
rect 22 11 30 13
rect 22 10 26 11
rect 24 9 26 10
rect 28 9 30 11
rect 24 7 30 9
<< pdif >>
rect 23 69 31 70
rect 2 67 9 69
rect 2 65 4 67
rect 6 65 9 67
rect 2 60 9 65
rect 2 58 4 60
rect 6 58 9 60
rect 2 45 9 58
rect 11 61 19 69
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 45 19 52
rect 21 68 31 69
rect 21 66 25 68
rect 27 66 31 68
rect 21 50 31 66
rect 33 61 41 70
rect 33 59 36 61
rect 38 59 41 61
rect 33 50 41 59
rect 43 68 50 70
rect 43 66 46 68
rect 48 66 50 68
rect 43 61 50 66
rect 43 59 46 61
rect 48 59 50 61
rect 43 50 50 59
rect 21 45 29 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 2 52 14 54
rect 16 52 17 54
rect 2 50 17 52
rect 2 21 6 50
rect 10 37 14 39
rect 33 50 46 54
rect 31 45 38 46
rect 31 43 33 45
rect 35 43 38 45
rect 31 42 38 43
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 10 25 22 29
rect 2 20 12 21
rect 2 18 8 20
rect 10 18 12 20
rect 2 17 12 18
rect 18 17 22 25
rect 34 31 38 42
rect 42 45 46 50
rect 42 43 43 45
rect 45 43 46 45
rect 42 41 46 43
rect 34 25 46 31
rect -2 11 58 12
rect -2 9 26 11
rect 28 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 13 10 15 30
rect 20 10 22 30
rect 32 13 34 30
rect 39 13 41 30
<< pmos >>
rect 9 45 11 69
rect 19 45 21 69
rect 31 50 33 70
rect 41 50 43 70
<< polyct0 >>
rect 21 35 23 37
<< polyct1 >>
rect 33 43 35 45
rect 43 43 45 45
rect 11 35 13 37
<< ndifct0 >>
rect 44 18 46 20
<< ndifct1 >>
rect 8 18 10 20
rect 26 9 28 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 65 6 67
rect 4 58 6 60
rect 25 66 27 68
rect 36 59 38 61
rect 46 66 48 68
rect 46 59 48 61
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
<< alu0 >>
rect 2 67 8 68
rect 2 65 4 67
rect 6 65 8 67
rect 23 66 25 68
rect 27 66 29 68
rect 23 65 29 66
rect 44 66 46 68
rect 48 66 50 68
rect 2 60 8 65
rect 2 58 4 60
rect 6 58 8 60
rect 2 57 8 58
rect 23 61 40 62
rect 23 59 36 61
rect 38 59 40 61
rect 23 58 40 59
rect 44 61 50 66
rect 44 59 46 61
rect 48 59 50 61
rect 44 58 50 59
rect 23 38 27 58
rect 19 37 30 38
rect 19 35 21 37
rect 23 35 30 37
rect 19 34 30 35
rect 26 21 30 34
rect 26 20 48 21
rect 26 18 44 20
rect 46 18 48 20
rect 26 17 48 18
<< labels >>
rlabel alu0 24 36 24 36 6 an
rlabel alu0 31 60 31 60 6 an
rlabel alu0 37 19 37 19 6 an
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 20 20 20 6 b
rlabel alu1 12 32 12 32 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 32 36 32 6 a2
rlabel alu1 36 52 36 52 6 a1
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a2
rlabel polyct1 44 44 44 44 6 a1
<< end >>
