magic
tech scmos
timestamp 1199203395
<< ab >>
rect 0 0 24 72
<< nwell >>
rect -5 32 29 77
<< pwell >>
rect -5 -5 29 32
<< poly >>
rect 12 57 14 61
rect 12 36 14 39
rect 4 34 14 36
rect 4 32 6 34
rect 8 32 14 34
rect 4 30 14 32
rect 12 26 14 30
rect 12 2 14 6
<< ndif >>
rect 3 24 12 26
rect 3 22 5 24
rect 7 22 12 24
rect 3 17 12 22
rect 3 15 5 17
rect 7 15 12 17
rect 3 6 12 15
rect 14 17 22 26
rect 14 15 18 17
rect 20 15 22 17
rect 14 10 22 15
rect 14 8 18 10
rect 20 8 22 10
rect 14 6 22 8
<< pdif >>
rect 3 67 10 69
rect 3 65 6 67
rect 8 65 10 67
rect 3 59 10 65
rect 3 57 6 59
rect 8 57 10 59
rect 3 51 12 57
rect 3 49 6 51
rect 8 49 12 51
rect 3 43 12 49
rect 3 41 6 43
rect 8 41 12 43
rect 3 39 12 41
rect 14 51 22 57
rect 14 49 18 51
rect 20 49 22 51
rect 14 43 22 49
rect 14 41 18 43
rect 20 41 22 43
rect 14 39 22 41
<< alu1 >>
rect -2 67 26 72
rect -2 65 6 67
rect 8 65 17 67
rect 19 65 26 67
rect -2 64 26 65
rect 17 51 22 59
rect 17 49 18 51
rect 20 49 22 51
rect 17 43 22 49
rect 17 41 18 43
rect 20 41 22 43
rect 17 27 22 41
rect 2 24 22 27
rect 2 22 5 24
rect 7 22 22 24
rect 2 21 22 22
rect 2 17 8 21
rect 2 15 5 17
rect 7 15 8 17
rect 2 13 8 15
rect -2 0 26 8
<< ntie >>
rect 15 67 21 69
rect 15 65 17 67
rect 19 65 21 67
rect 15 63 21 65
<< nmos >>
rect 12 6 14 26
<< pmos >>
rect 12 39 14 57
<< polyct0 >>
rect 6 32 8 34
<< ndifct0 >>
rect 18 15 20 17
rect 18 8 20 10
<< ndifct1 >>
rect 5 22 7 24
rect 5 15 7 17
<< ntiect1 >>
rect 17 65 19 67
<< pdifct0 >>
rect 6 57 8 59
rect 6 49 8 51
rect 6 41 8 43
<< pdifct1 >>
rect 6 65 8 67
rect 18 49 20 51
rect 18 41 20 43
<< alu0 >>
rect 4 59 10 64
rect 4 57 6 59
rect 8 57 10 59
rect 4 51 10 57
rect 4 49 6 51
rect 8 49 10 51
rect 4 43 10 49
rect 4 41 6 43
rect 8 41 10 43
rect 4 34 10 41
rect 4 32 6 34
rect 8 32 10 34
rect 4 31 10 32
rect 16 17 22 18
rect 16 15 18 17
rect 20 15 22 17
rect 16 10 22 15
rect 16 8 18 10
rect 20 8 22 10
<< labels >>
rlabel alu1 4 20 4 20 6 z
rlabel alu1 12 4 12 4 6 vss
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 68 12 68 6 vdd
rlabel alu1 20 40 20 40 6 z
<< end >>
