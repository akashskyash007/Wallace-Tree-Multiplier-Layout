magic
tech scmos
timestamp 1199542102
<< ab >>
rect 0 0 40 100
<< nwell >>
rect -5 48 45 105
<< pwell >>
rect -5 -5 45 48
<< poly >>
rect 13 94 15 98
rect 25 94 27 98
rect 13 33 15 55
rect 25 33 27 67
rect 7 31 27 33
rect 7 29 9 31
rect 11 29 27 31
rect 7 27 27 29
rect 13 24 15 27
rect 25 24 27 27
rect 13 2 15 6
rect 25 2 27 6
<< ndif >>
rect 5 11 13 24
rect 5 9 7 11
rect 9 9 13 11
rect 5 6 13 9
rect 15 21 25 24
rect 15 19 19 21
rect 21 19 25 21
rect 15 6 25 19
rect 27 21 35 24
rect 27 19 31 21
rect 33 19 35 21
rect 27 11 35 19
rect 27 9 31 11
rect 33 9 35 11
rect 27 6 35 9
<< pdif >>
rect 5 91 13 94
rect 5 89 7 91
rect 9 89 13 91
rect 5 55 13 89
rect 15 81 25 94
rect 15 79 19 81
rect 21 79 25 81
rect 15 71 25 79
rect 15 69 19 71
rect 21 69 25 71
rect 15 67 25 69
rect 27 91 35 94
rect 27 89 31 91
rect 33 89 35 91
rect 27 81 35 89
rect 27 79 31 81
rect 33 79 35 81
rect 27 71 35 79
rect 27 69 31 71
rect 33 69 35 71
rect 27 67 35 69
rect 15 61 23 67
rect 15 59 19 61
rect 21 59 23 61
rect 15 55 23 59
<< alu1 >>
rect -2 91 42 100
rect -2 89 7 91
rect 9 89 31 91
rect 33 89 42 91
rect -2 88 42 89
rect 8 31 12 83
rect 8 29 9 31
rect 11 29 12 31
rect 8 17 12 29
rect 18 81 22 83
rect 18 79 19 81
rect 21 79 22 81
rect 18 71 22 79
rect 18 69 19 71
rect 21 69 22 71
rect 18 61 22 69
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 71 34 79
rect 30 69 31 71
rect 33 69 34 71
rect 30 67 34 69
rect 18 59 19 61
rect 21 59 22 61
rect 18 21 22 59
rect 18 19 19 21
rect 21 19 22 21
rect 18 17 22 19
rect 30 21 34 23
rect 30 19 31 21
rect 33 19 34 21
rect 30 12 34 19
rect -2 11 42 12
rect -2 9 7 11
rect 9 9 31 11
rect 33 9 42 11
rect -2 0 42 9
<< nmos >>
rect 13 6 15 24
rect 25 6 27 24
<< pmos >>
rect 13 55 15 94
rect 25 67 27 94
<< polyct1 >>
rect 9 29 11 31
<< ndifct1 >>
rect 7 9 9 11
rect 19 19 21 21
rect 31 19 33 21
rect 31 9 33 11
<< pdifct1 >>
rect 7 89 9 91
rect 19 79 21 81
rect 19 69 21 71
rect 31 89 33 91
rect 31 79 33 81
rect 31 69 33 71
rect 19 59 21 61
<< labels >>
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 10 50 10 50 6 i
rlabel alu1 20 50 20 50 6 nq
rlabel alu1 20 94 20 94 6 vdd
<< end >>
