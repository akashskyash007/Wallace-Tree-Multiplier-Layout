magic
tech scmos
timestamp 1199203311
<< ab >>
rect 0 0 88 80
<< nwell >>
rect -5 36 93 88
<< pwell >>
rect -5 -8 93 36
<< poly >>
rect 9 70 11 74
rect 21 70 23 74
rect 28 70 30 74
rect 35 70 37 74
rect 42 70 44 74
rect 52 70 54 74
rect 59 70 61 74
rect 66 70 68 74
rect 73 70 75 74
rect 21 43 23 46
rect 9 33 11 42
rect 18 41 24 43
rect 18 39 20 41
rect 22 39 24 41
rect 18 37 24 39
rect 9 31 15 33
rect 9 29 11 31
rect 13 29 15 31
rect 9 27 15 29
rect 9 24 11 27
rect 21 22 23 37
rect 28 31 30 46
rect 35 37 37 46
rect 42 43 44 46
rect 52 43 54 46
rect 42 41 55 43
rect 49 37 55 41
rect 35 35 41 37
rect 39 31 41 35
rect 49 35 51 37
rect 53 35 55 37
rect 49 33 55 35
rect 27 29 33 31
rect 27 27 29 29
rect 31 27 33 29
rect 27 25 33 27
rect 39 29 45 31
rect 39 27 41 29
rect 43 27 45 29
rect 39 25 45 27
rect 31 22 33 25
rect 43 22 45 25
rect 53 22 55 33
rect 59 27 61 46
rect 66 37 68 46
rect 73 43 75 46
rect 73 41 82 43
rect 76 39 78 41
rect 80 39 82 41
rect 76 37 82 39
rect 65 35 71 37
rect 65 33 67 35
rect 69 33 71 35
rect 65 31 71 33
rect 59 25 67 27
rect 65 23 67 25
rect 65 21 71 23
rect 65 19 67 21
rect 69 19 71 21
rect 65 17 71 19
rect 9 6 11 10
rect 21 10 23 15
rect 31 10 33 15
rect 43 10 45 15
rect 53 10 55 15
<< ndif >>
rect 2 21 9 24
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 10 9 17
rect 11 22 19 24
rect 11 15 21 22
rect 23 20 31 22
rect 23 18 26 20
rect 28 18 31 20
rect 23 15 31 18
rect 33 15 43 22
rect 45 20 53 22
rect 45 18 48 20
rect 50 18 53 20
rect 45 15 53 18
rect 55 15 63 22
rect 11 11 19 15
rect 11 10 15 11
rect 13 9 15 10
rect 17 9 19 11
rect 35 11 41 15
rect 13 7 19 9
rect 35 9 37 11
rect 39 9 41 11
rect 57 11 63 15
rect 35 7 41 9
rect 57 9 59 11
rect 61 9 63 11
rect 57 7 63 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 21 70
rect 11 66 15 68
rect 17 66 21 68
rect 11 46 21 66
rect 23 46 28 70
rect 30 46 35 70
rect 37 46 42 70
rect 44 61 52 70
rect 44 59 47 61
rect 49 59 52 61
rect 44 46 52 59
rect 54 46 59 70
rect 61 46 66 70
rect 68 46 73 70
rect 75 68 82 70
rect 75 66 78 68
rect 80 66 82 68
rect 75 61 82 66
rect 75 59 78 61
rect 80 59 82 61
rect 75 46 82 59
rect 11 42 16 46
<< alu1 >>
rect -2 81 90 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 90 81
rect -2 68 90 79
rect 2 53 6 63
rect 2 51 4 53
rect 2 46 6 51
rect 2 44 4 46
rect 2 23 6 44
rect 58 54 62 63
rect 18 50 79 54
rect 18 41 23 50
rect 18 39 20 41
rect 22 39 23 41
rect 18 37 23 39
rect 29 42 70 46
rect 29 31 33 42
rect 41 37 55 38
rect 41 35 51 37
rect 53 35 55 37
rect 41 34 55 35
rect 66 35 70 42
rect 66 33 67 35
rect 69 33 70 35
rect 74 41 79 50
rect 74 39 78 41
rect 74 33 79 39
rect 66 31 70 33
rect 2 21 14 23
rect 2 19 4 21
rect 6 19 14 21
rect 2 17 14 19
rect 26 29 33 31
rect 26 27 29 29
rect 31 27 33 29
rect 26 25 33 27
rect 39 29 61 30
rect 39 27 41 29
rect 43 27 61 29
rect 39 26 61 27
rect 57 22 61 26
rect 57 21 71 22
rect 57 19 67 21
rect 69 19 71 21
rect 57 18 71 19
rect -2 11 90 12
rect -2 9 15 11
rect 17 9 37 11
rect 39 9 59 11
rect 61 9 90 11
rect -2 1 90 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 90 1
rect -2 -2 90 -1
<< ptie >>
rect 0 1 88 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 88 1
rect 0 -3 88 -1
<< ntie >>
rect 0 81 88 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 88 81
rect 0 77 88 79
<< nmos >>
rect 9 10 11 24
rect 21 15 23 22
rect 31 15 33 22
rect 43 15 45 22
rect 53 15 55 22
<< pmos >>
rect 9 42 11 70
rect 21 46 23 70
rect 28 46 30 70
rect 35 46 37 70
rect 42 46 44 70
rect 52 46 54 70
rect 59 46 61 70
rect 66 46 68 70
rect 73 46 75 70
<< polyct0 >>
rect 11 29 13 31
rect 79 39 80 41
<< polyct1 >>
rect 20 39 22 41
rect 51 35 53 37
rect 29 27 31 29
rect 41 27 43 29
rect 78 39 79 41
rect 67 33 69 35
rect 67 19 69 21
<< ndifct0 >>
rect 26 18 28 20
rect 48 18 50 20
<< ndifct1 >>
rect 4 19 6 21
rect 15 9 17 11
rect 37 9 39 11
rect 59 9 61 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
<< pdifct0 >>
rect 15 66 17 68
rect 47 59 49 61
rect 78 66 80 68
rect 78 59 80 61
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 13 66 15 68
rect 17 66 19 68
rect 13 65 19 66
rect 76 66 78 68
rect 80 66 82 68
rect 10 61 51 62
rect 10 59 47 61
rect 49 59 51 61
rect 10 58 51 59
rect 6 42 7 55
rect 10 31 14 58
rect 76 61 82 66
rect 76 59 78 61
rect 80 59 82 61
rect 76 58 82 59
rect 79 41 82 43
rect 80 39 82 41
rect 79 37 82 39
rect 10 29 11 31
rect 13 29 22 31
rect 10 27 22 29
rect 18 21 22 27
rect 18 20 52 21
rect 18 18 26 20
rect 28 18 48 20
rect 50 18 52 20
rect 18 17 52 18
<< labels >>
rlabel alu0 12 44 12 44 6 zn
rlabel alu0 35 19 35 19 6 zn
rlabel alu0 30 60 30 60 6 zn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 28 28 28 6 b
rlabel alu1 20 44 20 44 6 a
rlabel alu1 28 52 28 52 6 a
rlabel alu1 44 6 44 6 6 vss
rlabel alu1 44 28 44 28 6 c
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 36 44 36 6 d
rlabel alu1 44 44 44 44 6 b
rlabel alu1 44 52 44 52 6 a
rlabel alu1 36 52 36 52 6 a
rlabel alu1 44 74 44 74 6 vdd
rlabel alu1 52 28 52 28 6 c
rlabel alu1 60 20 60 20 6 c
rlabel polyct1 68 20 68 20 6 c
rlabel polyct1 52 36 52 36 6 d
rlabel alu1 52 44 52 44 6 b
rlabel alu1 60 44 60 44 6 b
rlabel alu1 68 36 68 36 6 b
rlabel alu1 68 52 68 52 6 a
rlabel alu1 52 52 52 52 6 a
rlabel alu1 60 56 60 56 6 a
rlabel alu1 76 44 76 44 6 a
<< end >>
