magic
tech scmos
timestamp 1199201702
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 9 61 11 65
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 41 39
rect 49 37 51 43
rect 59 40 61 43
rect 58 38 64 40
rect 9 30 11 37
rect 19 30 21 37
rect 29 35 33 37
rect 35 35 37 37
rect 29 33 37 35
rect 48 35 54 37
rect 48 33 50 35
rect 52 33 54 35
rect 29 30 31 33
rect 41 31 54 33
rect 58 36 60 38
rect 62 36 64 38
rect 58 34 64 36
rect 9 15 11 19
rect 41 22 43 31
rect 58 27 60 34
rect 68 29 74 31
rect 68 27 70 29
rect 72 27 74 29
rect 48 25 60 27
rect 48 22 50 25
rect 58 22 60 25
rect 65 25 74 27
rect 65 22 67 25
rect 19 6 21 10
rect 29 6 31 10
rect 41 6 43 11
rect 48 6 50 11
rect 58 6 60 11
rect 65 6 67 11
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 4 19 9 24
rect 11 23 19 30
rect 11 21 14 23
rect 16 21 19 23
rect 11 19 19 21
rect 13 10 19 19
rect 21 28 29 30
rect 21 26 24 28
rect 26 26 29 28
rect 21 21 29 26
rect 21 19 24 21
rect 26 19 29 21
rect 21 10 29 19
rect 31 22 39 30
rect 31 20 34 22
rect 36 20 41 22
rect 31 14 41 20
rect 31 12 34 14
rect 36 12 41 14
rect 31 11 41 12
rect 43 11 48 22
rect 50 20 58 22
rect 50 18 53 20
rect 55 18 58 20
rect 50 11 58 18
rect 60 11 65 22
rect 67 15 75 22
rect 67 13 70 15
rect 72 13 75 15
rect 67 11 75 13
rect 31 10 39 11
<< pdif >>
rect 14 61 19 70
rect 2 59 9 61
rect 2 57 4 59
rect 6 57 9 59
rect 2 52 9 57
rect 2 50 4 52
rect 6 50 9 52
rect 2 42 9 50
rect 11 59 19 61
rect 11 57 14 59
rect 16 57 19 59
rect 11 52 19 57
rect 11 50 14 52
rect 16 50 19 52
rect 11 42 19 50
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 42 39 52
rect 41 68 49 70
rect 41 66 44 68
rect 46 66 49 68
rect 41 61 49 66
rect 41 59 44 61
rect 46 59 49 61
rect 41 43 49 59
rect 51 61 59 70
rect 51 59 54 61
rect 56 59 59 61
rect 51 54 59 59
rect 51 52 54 54
rect 56 52 59 54
rect 51 43 59 52
rect 61 63 67 70
rect 61 61 69 63
rect 61 59 64 61
rect 66 59 69 61
rect 61 54 69 59
rect 61 52 64 54
rect 66 52 69 54
rect 61 43 69 52
rect 41 42 47 43
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 12 59 18 60
rect 12 57 14 59
rect 16 57 18 59
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 12 54 18 57
rect 33 54 38 59
rect 12 52 34 54
rect 36 52 38 54
rect 12 50 14 52
rect 16 50 38 52
rect 12 49 22 50
rect 18 39 22 49
rect 2 38 22 39
rect 2 34 27 38
rect 2 28 7 34
rect 2 26 4 28
rect 6 26 7 28
rect 2 24 7 26
rect 23 28 27 34
rect 23 26 24 28
rect 26 26 27 28
rect 23 21 27 26
rect 23 19 24 21
rect 26 19 27 21
rect 23 17 27 19
rect 49 35 54 39
rect 49 33 50 35
rect 52 33 54 35
rect 58 38 63 47
rect 58 36 60 38
rect 62 36 71 38
rect 58 34 71 36
rect 49 30 54 33
rect 49 29 74 30
rect 49 27 70 29
rect 72 27 74 29
rect 49 26 74 27
rect -2 1 82 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 9 19 11 30
rect 19 10 21 30
rect 29 10 31 30
rect 41 11 43 22
rect 48 11 50 22
rect 58 11 60 22
rect 65 11 67 22
<< pmos >>
rect 9 42 11 61
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 43 51 70
rect 59 43 61 70
<< polyct0 >>
rect 33 35 35 37
<< polyct1 >>
rect 50 33 52 35
rect 60 36 62 38
rect 70 27 72 29
<< ndifct0 >>
rect 14 21 16 23
rect 34 20 36 22
rect 34 12 36 14
rect 53 18 55 20
rect 70 13 72 15
<< ndifct1 >>
rect 4 26 6 28
rect 24 26 26 28
rect 24 19 26 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 57 6 59
rect 4 50 6 52
rect 24 66 26 68
rect 24 59 26 61
rect 44 66 46 68
rect 44 59 46 61
rect 54 59 56 61
rect 54 52 56 54
rect 64 59 66 61
rect 64 52 66 54
<< pdifct1 >>
rect 14 57 16 59
rect 14 50 16 52
rect 34 59 36 61
rect 34 52 36 54
<< alu0 >>
rect 3 59 7 68
rect 22 66 24 68
rect 26 66 28 68
rect 22 61 28 66
rect 42 66 44 68
rect 46 66 48 68
rect 3 57 4 59
rect 6 57 7 59
rect 3 52 7 57
rect 3 50 4 52
rect 6 50 7 52
rect 3 48 7 50
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 42 61 48 66
rect 42 59 44 61
rect 46 59 48 61
rect 42 58 48 59
rect 53 61 57 63
rect 53 59 54 61
rect 56 59 57 61
rect 53 54 57 59
rect 41 52 54 54
rect 56 52 57 54
rect 41 50 57 52
rect 63 61 67 68
rect 63 59 64 61
rect 66 59 67 61
rect 63 54 67 59
rect 63 52 64 54
rect 66 52 67 54
rect 63 50 67 52
rect 41 38 45 50
rect 31 37 45 38
rect 31 35 33 37
rect 35 35 45 37
rect 31 34 45 35
rect 13 23 17 25
rect 13 21 14 23
rect 16 21 17 23
rect 13 12 17 21
rect 33 22 37 24
rect 33 20 34 22
rect 36 20 37 22
rect 33 14 37 20
rect 41 21 45 34
rect 41 20 57 21
rect 41 18 53 20
rect 55 18 57 20
rect 41 17 57 18
rect 33 12 34 14
rect 36 12 37 14
rect 69 15 73 17
rect 69 13 70 15
rect 72 13 73 15
rect 69 12 73 13
<< labels >>
rlabel alu0 49 19 49 19 6 zn
rlabel alu0 38 36 38 36 6 zn
rlabel alu0 55 56 55 56 6 zn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 36 12 36 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 52 32 52 32 6 a
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 28 60 28 6 a
rlabel alu1 68 36 68 36 6 b
rlabel alu1 68 28 68 28 6 a
rlabel alu1 60 44 60 44 6 b
<< end >>
