magic
tech scmos
timestamp 1199202320
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 57 11 61
rect 19 57 21 61
rect 29 59 31 64
rect 39 59 41 64
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 33 41 35
rect 9 26 11 33
rect 19 26 21 33
rect 29 31 31 33
rect 33 31 41 33
rect 29 29 41 31
rect 29 26 31 29
rect 39 26 41 29
rect 9 2 11 6
rect 19 2 21 6
rect 29 2 31 6
rect 39 2 41 6
<< ndif >>
rect 2 17 9 26
rect 2 15 4 17
rect 6 15 9 17
rect 2 10 9 15
rect 2 8 4 10
rect 6 8 9 10
rect 2 6 9 8
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 11 15 14 17
rect 16 15 19 17
rect 11 6 19 15
rect 21 17 29 26
rect 21 15 24 17
rect 26 15 29 17
rect 21 10 29 15
rect 21 8 24 10
rect 26 8 29 10
rect 21 6 29 8
rect 31 24 39 26
rect 31 22 34 24
rect 36 22 39 24
rect 31 17 39 22
rect 31 15 34 17
rect 36 15 39 17
rect 31 6 39 15
rect 41 17 49 26
rect 41 15 45 17
rect 47 15 49 17
rect 41 10 49 15
rect 41 8 45 10
rect 47 8 49 10
rect 41 6 49 8
<< pdif >>
rect 24 57 29 59
rect 2 55 9 57
rect 2 53 4 55
rect 6 53 9 55
rect 2 48 9 53
rect 2 46 4 48
rect 6 46 9 48
rect 2 38 9 46
rect 11 49 19 57
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 55 29 57
rect 21 53 24 55
rect 26 53 29 55
rect 21 48 29 53
rect 21 46 24 48
rect 26 46 29 48
rect 21 38 29 46
rect 31 49 39 59
rect 31 47 34 49
rect 36 47 39 49
rect 31 42 39 47
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 56 49 59
rect 41 54 44 56
rect 46 54 49 56
rect 41 49 49 54
rect 41 47 44 49
rect 46 47 49 49
rect 41 38 49 47
<< alu1 >>
rect -2 67 58 72
rect -2 65 5 67
rect 7 65 19 67
rect 21 65 58 67
rect -2 64 58 65
rect 33 49 38 51
rect 33 47 34 49
rect 36 47 38 49
rect 33 42 38 47
rect 9 40 14 42
rect 16 40 34 42
rect 36 40 38 42
rect 9 38 38 40
rect 18 26 22 38
rect 42 34 47 43
rect 29 33 47 34
rect 29 31 31 33
rect 33 31 47 33
rect 29 30 47 31
rect 9 24 39 26
rect 9 22 14 24
rect 16 22 34 24
rect 36 22 39 24
rect 12 17 17 22
rect 12 15 14 17
rect 16 15 17 17
rect 12 13 17 15
rect 33 17 39 22
rect 33 15 34 17
rect 36 15 39 17
rect 33 13 39 15
rect -2 0 58 8
<< ntie >>
rect 3 67 23 69
rect 3 65 5 67
rect 7 65 19 67
rect 21 65 23 67
rect 3 63 23 65
<< nmos >>
rect 9 6 11 26
rect 19 6 21 26
rect 29 6 31 26
rect 39 6 41 26
<< pmos >>
rect 9 38 11 57
rect 19 38 21 57
rect 29 38 31 59
rect 39 38 41 59
<< polyct1 >>
rect 31 31 33 33
<< ndifct0 >>
rect 4 15 6 17
rect 4 8 6 10
rect 24 15 26 17
rect 24 8 26 10
rect 45 15 47 17
rect 45 8 47 10
<< ndifct1 >>
rect 14 22 16 24
rect 14 15 16 17
rect 34 22 36 24
rect 34 15 36 17
<< ntiect1 >>
rect 5 65 7 67
rect 19 65 21 67
<< pdifct0 >>
rect 4 53 6 55
rect 4 46 6 48
rect 14 47 16 49
rect 24 53 26 55
rect 24 46 26 48
rect 44 54 46 56
rect 44 47 46 49
<< pdifct1 >>
rect 14 40 16 42
rect 34 47 36 49
rect 34 40 36 42
<< alu0 >>
rect 2 55 8 64
rect 2 53 4 55
rect 6 53 8 55
rect 2 48 8 53
rect 22 55 28 64
rect 22 53 24 55
rect 26 53 28 55
rect 2 46 4 48
rect 6 46 8 48
rect 2 45 8 46
rect 13 49 17 51
rect 13 47 14 49
rect 16 47 17 49
rect 13 42 17 47
rect 22 48 28 53
rect 42 56 48 64
rect 42 54 44 56
rect 46 54 48 56
rect 22 46 24 48
rect 26 46 28 48
rect 22 45 28 46
rect 42 49 48 54
rect 42 47 44 49
rect 46 47 48 49
rect 42 46 48 47
rect 2 17 8 18
rect 2 15 4 17
rect 6 15 8 17
rect 2 10 8 15
rect 22 17 28 18
rect 22 15 24 17
rect 26 15 28 17
rect 2 8 4 10
rect 6 8 8 10
rect 22 10 28 15
rect 43 17 49 18
rect 43 15 45 17
rect 47 15 49 17
rect 22 8 24 10
rect 26 8 28 10
rect 43 10 49 15
rect 43 8 45 10
rect 47 8 49 10
<< labels >>
rlabel alu1 12 24 12 24 6 z
rlabel alu1 20 32 20 32 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 36 32 36 32 6 a
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 36 44 36 6 a
<< end >>
