magic
tech scmos
timestamp 1199973105
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -5 40 101 97
<< pwell >>
rect -5 -9 101 40
<< poly >>
rect 2 81 11 83
rect 2 79 7 81
rect 9 79 11 81
rect 2 77 11 79
rect 9 74 11 77
rect 21 81 30 83
rect 21 79 26 81
rect 28 79 30 81
rect 21 77 30 79
rect 34 77 43 83
rect 21 74 23 77
rect 41 74 43 77
rect 53 77 62 83
rect 66 81 75 83
rect 66 79 68 81
rect 70 79 75 81
rect 66 77 75 79
rect 53 74 55 77
rect 73 74 75 77
rect 85 77 94 83
rect 85 74 87 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 73 43 75 46
rect 85 43 87 46
rect 2 37 14 43
rect 18 41 30 43
rect 18 39 20 41
rect 22 39 30 41
rect 18 37 30 39
rect 34 41 46 43
rect 34 39 39 41
rect 41 39 46 41
rect 34 37 46 39
rect 50 37 62 43
rect 66 37 78 43
rect 82 41 94 43
rect 82 39 87 41
rect 89 39 94 41
rect 82 37 94 39
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 73 34 75 37
rect 85 34 87 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 73 11 75 14
rect 53 9 62 11
rect 53 7 55 9
rect 57 7 62 9
rect 53 5 62 7
rect 66 5 75 11
rect 85 11 87 14
rect 85 5 94 11
<< ndif >>
rect 2 14 9 34
rect 11 25 21 34
rect 11 23 15 25
rect 17 23 21 25
rect 11 18 21 23
rect 11 16 15 18
rect 17 16 21 18
rect 11 14 21 16
rect 23 32 30 34
rect 23 30 26 32
rect 28 30 30 32
rect 23 25 30 30
rect 23 23 26 25
rect 28 23 30 25
rect 23 14 30 23
rect 34 29 41 34
rect 34 27 36 29
rect 38 27 41 29
rect 34 22 41 27
rect 34 20 36 22
rect 38 20 41 22
rect 34 14 41 20
rect 43 32 53 34
rect 43 30 47 32
rect 49 30 53 32
rect 43 14 53 30
rect 55 29 62 34
rect 55 27 58 29
rect 60 27 62 29
rect 55 14 62 27
rect 66 21 73 34
rect 66 19 68 21
rect 70 19 73 21
rect 66 14 73 19
rect 75 21 85 34
rect 75 19 79 21
rect 81 19 85 21
rect 75 14 85 19
rect 87 28 94 34
rect 87 26 90 28
rect 92 26 94 28
rect 87 21 94 26
rect 87 19 90 21
rect 92 19 94 21
rect 87 14 94 19
rect 13 2 19 14
rect 45 2 51 14
rect 77 12 79 14
rect 81 12 83 14
rect 77 2 83 12
<< pdif >>
rect 13 74 19 86
rect 45 74 51 86
rect 77 74 83 86
rect 2 46 9 74
rect 11 72 21 74
rect 11 70 15 72
rect 17 70 21 72
rect 11 65 21 70
rect 11 63 15 65
rect 17 63 21 65
rect 11 46 21 63
rect 23 57 30 74
rect 23 55 26 57
rect 28 55 30 57
rect 23 50 30 55
rect 23 48 26 50
rect 28 48 30 50
rect 23 46 30 48
rect 34 69 41 74
rect 34 67 36 69
rect 38 67 41 69
rect 34 46 41 67
rect 43 46 53 74
rect 55 69 62 74
rect 55 67 58 69
rect 60 67 62 69
rect 55 53 62 67
rect 55 51 58 53
rect 60 51 62 53
rect 55 46 62 51
rect 66 69 73 74
rect 66 67 68 69
rect 70 67 73 69
rect 66 53 73 67
rect 66 51 68 53
rect 70 51 73 53
rect 66 46 73 51
rect 75 58 85 74
rect 75 56 79 58
rect 81 56 85 58
rect 75 50 85 56
rect 75 48 79 50
rect 81 48 85 50
rect 75 46 85 48
rect 87 72 94 74
rect 87 70 90 72
rect 92 70 94 72
rect 87 65 94 70
rect 87 63 90 65
rect 92 63 94 65
rect 87 46 94 63
<< alu1 >>
rect -2 89 98 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 73 87 87 89
rect 89 87 91 89
rect 93 87 98 89
rect -2 86 98 87
rect 6 81 10 86
rect 6 79 7 81
rect 9 79 10 81
rect 6 77 10 79
rect 14 81 18 86
rect 14 79 15 81
rect 17 79 18 81
rect 14 72 18 79
rect 89 81 93 86
rect 89 79 90 81
rect 92 79 93 81
rect 14 70 15 72
rect 17 70 18 72
rect 89 72 93 79
rect 89 70 90 72
rect 92 70 93 72
rect 14 65 18 70
rect 14 63 15 65
rect 17 63 18 65
rect 14 61 18 63
rect 89 65 93 70
rect 89 63 90 65
rect 92 63 93 65
rect 14 33 18 55
rect 89 61 93 63
rect 46 53 72 54
rect 46 51 58 53
rect 60 51 68 53
rect 70 51 72 53
rect 46 50 72 51
rect 14 25 18 27
rect 14 23 15 25
rect 17 23 18 25
rect 14 18 18 23
rect 46 32 50 50
rect 46 30 47 32
rect 49 30 50 32
rect 86 41 90 55
rect 86 39 87 41
rect 89 39 90 41
rect 86 33 90 39
rect 46 25 50 30
rect 78 21 82 23
rect 78 19 79 21
rect 81 19 82 21
rect 14 16 15 18
rect 17 16 18 18
rect 14 9 18 16
rect 14 7 15 9
rect 17 7 18 9
rect 14 2 18 7
rect 78 14 82 19
rect 78 12 79 14
rect 81 12 82 14
rect 78 9 82 12
rect 78 7 79 9
rect 81 7 82 9
rect 78 2 82 7
rect -2 1 98 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 73 -1 87 1
rect 89 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< alu2 >>
rect -2 89 98 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 71 89
rect 73 87 87 89
rect 89 87 98 89
rect -2 81 98 87
rect -2 79 15 81
rect 17 79 90 81
rect 92 79 98 81
rect -2 76 98 79
rect -2 9 98 12
rect -2 7 15 9
rect 17 7 79 9
rect 81 7 98 9
rect -2 1 98 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 71 1
rect 73 -1 87 1
rect 89 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 71 3
rect 57 -1 59 1
rect 61 -1 67 1
rect 69 -1 71 1
rect 57 -3 71 -1
rect 89 1 96 3
rect 89 -1 91 1
rect 93 -1 96 1
rect 89 -3 96 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 71 91
rect 57 87 59 89
rect 61 87 67 89
rect 69 87 71 89
rect 57 85 71 87
rect 89 89 96 91
rect 89 87 91 89
rect 93 87 96 89
rect 89 85 96 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
rect 73 14 75 34
rect 85 14 87 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
rect 73 46 75 74
rect 85 46 87 74
<< polyct0 >>
rect 26 79 28 81
rect 68 79 70 81
rect 20 39 22 41
rect 39 39 41 41
rect 55 7 57 9
<< polyct1 >>
rect 7 79 9 81
rect 87 39 89 41
<< ndifct0 >>
rect 26 30 28 32
rect 26 23 28 25
rect 36 27 38 29
rect 36 20 38 22
rect 58 27 60 29
rect 68 19 70 21
rect 90 26 92 28
rect 90 19 92 21
<< ndifct1 >>
rect 15 23 17 25
rect 15 16 17 18
rect 47 30 49 32
rect 79 19 81 21
rect 79 12 81 14
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
rect 67 87 69 89
rect 91 87 93 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 91 -1 93 1
<< pdifct0 >>
rect 26 55 28 57
rect 26 48 28 50
rect 36 67 38 69
rect 58 67 60 69
rect 68 67 70 69
rect 79 56 81 58
rect 79 48 81 50
<< pdifct1 >>
rect 15 70 17 72
rect 15 63 17 65
rect 58 51 60 53
rect 68 51 70 53
rect 90 70 92 72
rect 90 63 92 65
<< alu0 >>
rect 24 81 72 82
rect 24 79 26 81
rect 28 79 68 81
rect 70 79 72 81
rect 24 78 72 79
rect 18 69 40 70
rect 18 67 36 69
rect 38 67 40 69
rect 18 66 40 67
rect 56 69 72 70
rect 56 67 58 69
rect 60 67 68 69
rect 70 67 72 69
rect 56 66 72 67
rect 25 57 29 59
rect 25 55 26 57
rect 28 55 29 57
rect 25 50 29 55
rect 38 58 82 62
rect 25 48 26 50
rect 28 48 34 50
rect 25 46 34 48
rect 18 41 24 42
rect 18 39 20 41
rect 22 39 24 41
rect 18 38 24 39
rect 30 34 34 46
rect 38 41 42 58
rect 78 56 79 58
rect 81 56 82 58
rect 38 39 39 41
rect 41 39 42 41
rect 38 37 42 39
rect 78 50 82 56
rect 25 32 39 34
rect 25 30 26 32
rect 28 30 39 32
rect 25 25 29 30
rect 25 23 26 25
rect 28 23 29 25
rect 25 21 29 23
rect 35 29 39 30
rect 35 27 36 29
rect 38 27 39 29
rect 35 22 39 27
rect 78 48 79 50
rect 81 48 82 50
rect 78 30 82 48
rect 56 29 93 30
rect 56 27 58 29
rect 60 28 93 29
rect 60 27 90 28
rect 56 26 90 27
rect 92 26 93 28
rect 35 20 36 22
rect 38 21 72 22
rect 38 20 68 21
rect 35 19 68 20
rect 70 19 72 21
rect 35 18 72 19
rect 54 9 58 18
rect 54 7 55 9
rect 57 7 58 9
rect 54 5 58 7
rect 89 21 93 26
rect 89 19 90 21
rect 92 19 93 21
rect 89 17 93 19
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 71 87 73 89
rect 87 87 89 89
rect 15 79 17 81
rect 90 79 92 81
rect 15 7 17 9
rect 79 7 81 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
rect 71 -1 73 1
rect 87 -1 89 1
<< labels >>
rlabel alu1 16 44 16 44 6 b
rlabel alu1 48 36 48 36 6 z
rlabel alu1 64 52 64 52 6 z
rlabel alu1 56 52 56 52 6 z
rlabel alu1 88 44 88 44 6 a
rlabel alu2 48 6 48 6 6 vss
rlabel alu2 48 82 48 82 6 vdd
<< end >>
