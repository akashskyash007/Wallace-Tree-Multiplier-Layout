magic
tech scmos
timestamp 1199543336
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 57 95 59 98
rect 11 85 13 88
rect 19 85 21 88
rect 27 85 29 88
rect 35 85 37 88
rect 11 43 13 55
rect 19 43 21 55
rect 27 43 29 55
rect 35 53 37 55
rect 35 51 43 53
rect 41 43 43 51
rect 57 43 59 55
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 47 41 59 43
rect 47 39 49 41
rect 51 39 59 41
rect 47 37 59 39
rect 11 25 13 37
rect 19 29 21 37
rect 31 29 33 37
rect 41 29 43 37
rect 19 27 25 29
rect 31 27 37 29
rect 41 27 49 29
rect 23 25 25 27
rect 35 25 37 27
rect 47 25 49 27
rect 57 25 59 37
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 47 12 49 15
rect 57 2 59 5
<< ndif >>
rect 3 15 11 25
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 15 23 19
rect 25 15 35 25
rect 37 21 47 25
rect 37 19 41 21
rect 43 19 47 21
rect 37 15 47 19
rect 49 15 57 25
rect 3 11 9 15
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 27 11 33 15
rect 27 9 29 11
rect 31 9 33 11
rect 51 9 57 15
rect 27 7 33 9
rect 49 7 57 9
rect 49 5 51 7
rect 53 5 57 7
rect 59 21 67 25
rect 59 19 63 21
rect 65 19 67 21
rect 59 5 67 19
rect 49 3 55 5
<< pdif >>
rect 39 91 57 95
rect 39 89 43 91
rect 45 89 51 91
rect 53 89 57 91
rect 39 85 57 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 55 19 85
rect 21 55 27 85
rect 29 55 35 85
rect 37 55 57 85
rect 59 81 67 95
rect 59 79 63 81
rect 65 79 67 81
rect 59 71 67 79
rect 59 69 63 71
rect 65 69 67 71
rect 59 61 67 69
rect 59 59 63 61
rect 65 59 67 61
rect 59 55 67 59
<< alu1 >>
rect -2 95 72 100
rect -2 93 5 95
rect 7 93 17 95
rect 19 93 29 95
rect 31 93 72 95
rect -2 91 72 93
rect -2 89 43 91
rect 45 89 51 91
rect 53 89 72 91
rect -2 88 72 89
rect 4 81 8 82
rect 58 81 66 82
rect 4 79 5 81
rect 7 79 52 81
rect 4 78 8 79
rect 8 41 12 72
rect 8 39 9 41
rect 11 39 12 41
rect 8 28 12 39
rect 18 41 22 72
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 28 41 32 72
rect 28 39 29 41
rect 31 39 32 41
rect 28 28 32 39
rect 38 41 42 72
rect 50 42 52 79
rect 38 39 39 41
rect 41 39 42 41
rect 38 28 42 39
rect 48 41 52 42
rect 48 39 49 41
rect 51 39 52 41
rect 48 38 52 39
rect 16 21 20 22
rect 40 21 44 22
rect 50 21 52 38
rect 16 19 17 21
rect 19 19 41 21
rect 43 19 52 21
rect 58 79 63 81
rect 65 79 66 81
rect 58 78 66 79
rect 58 72 62 78
rect 58 71 66 72
rect 58 69 63 71
rect 65 69 66 71
rect 58 68 66 69
rect 58 62 62 68
rect 58 61 66 62
rect 58 59 63 61
rect 65 59 66 61
rect 58 58 66 59
rect 58 22 62 58
rect 58 21 66 22
rect 58 19 63 21
rect 65 19 66 21
rect 16 18 20 19
rect 40 18 44 19
rect 58 18 66 19
rect -2 11 72 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 72 11
rect -2 7 72 9
rect -2 5 51 7
rect 53 5 72 7
rect -2 0 72 5
<< ntie >>
rect 3 95 33 97
rect 3 93 5 95
rect 7 93 17 95
rect 19 93 29 95
rect 31 93 33 95
rect 3 91 33 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 15 49 25
rect 57 5 59 25
<< pmos >>
rect 11 55 13 85
rect 19 55 21 85
rect 27 55 29 85
rect 35 55 37 85
rect 57 55 59 95
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 39 39 41 41
rect 49 39 51 41
<< ndifct1 >>
rect 17 19 19 21
rect 41 19 43 21
rect 5 9 7 11
rect 29 9 31 11
rect 51 5 53 7
rect 63 19 65 21
<< ntiect1 >>
rect 5 93 7 95
rect 17 93 19 95
rect 29 93 31 95
<< pdifct1 >>
rect 43 89 45 91
rect 51 89 53 91
rect 5 79 7 81
rect 63 79 65 81
rect 63 69 65 71
rect 63 59 65 61
<< labels >>
rlabel alu1 10 50 10 50 6 i3
rlabel alu1 30 50 30 50 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 50 40 50 6 i2
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 50 60 50 6 q
<< end >>
