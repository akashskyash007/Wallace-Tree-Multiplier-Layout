magic
tech scmos
timestamp 1199202606
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 14 61 16 66
rect 24 61 26 66
rect 34 61 36 66
rect 44 61 46 65
rect 14 39 16 43
rect 24 39 26 43
rect 9 37 26 39
rect 9 35 11 37
rect 13 35 26 37
rect 9 33 26 35
rect 14 30 16 33
rect 24 30 26 33
rect 34 39 36 43
rect 44 39 46 43
rect 34 37 47 39
rect 34 35 43 37
rect 45 35 47 37
rect 34 33 47 35
rect 34 30 36 33
rect 45 30 47 33
rect 14 10 16 15
rect 24 10 26 15
rect 45 15 47 19
rect 34 6 36 11
<< ndif >>
rect 9 22 14 30
rect 7 20 14 22
rect 7 18 9 20
rect 11 18 14 20
rect 7 15 14 18
rect 16 28 24 30
rect 16 26 19 28
rect 21 26 24 28
rect 16 15 24 26
rect 26 27 34 30
rect 26 25 29 27
rect 31 25 34 27
rect 26 20 34 25
rect 26 18 29 20
rect 31 18 34 20
rect 26 15 34 18
rect 29 11 34 15
rect 36 19 45 30
rect 47 28 54 30
rect 47 26 50 28
rect 52 26 54 28
rect 47 24 54 26
rect 47 19 52 24
rect 36 17 39 19
rect 41 17 43 19
rect 36 11 43 17
<< pdif >>
rect 6 59 14 61
rect 6 57 9 59
rect 11 57 14 59
rect 6 52 14 57
rect 6 50 9 52
rect 11 50 14 52
rect 6 43 14 50
rect 16 54 24 61
rect 16 52 19 54
rect 21 52 24 54
rect 16 47 24 52
rect 16 45 19 47
rect 21 45 24 47
rect 16 43 24 45
rect 26 59 34 61
rect 26 57 29 59
rect 31 57 34 59
rect 26 52 34 57
rect 26 50 29 52
rect 31 50 34 52
rect 26 43 34 50
rect 36 54 44 61
rect 36 52 39 54
rect 41 52 44 54
rect 36 47 44 52
rect 36 45 39 47
rect 41 45 44 47
rect 36 43 44 45
rect 46 59 54 61
rect 46 57 49 59
rect 51 57 54 59
rect 46 43 54 57
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 18 54 22 56
rect 18 52 19 54
rect 21 52 22 54
rect 18 47 22 52
rect 38 54 42 56
rect 38 52 39 54
rect 41 52 42 54
rect 18 45 19 47
rect 21 46 22 47
rect 38 47 42 52
rect 38 46 39 47
rect 21 45 39 46
rect 41 45 42 47
rect 18 42 42 45
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 2 25 6 33
rect 18 28 22 42
rect 50 38 54 47
rect 41 37 54 38
rect 41 35 43 37
rect 45 35 54 37
rect 41 33 54 35
rect 18 26 19 28
rect 21 26 22 28
rect 18 24 22 26
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 14 15 16 30
rect 24 15 26 30
rect 34 11 36 30
rect 45 19 47 30
<< pmos >>
rect 14 43 16 61
rect 24 43 26 61
rect 34 43 36 61
rect 44 43 46 61
<< polyct1 >>
rect 11 35 13 37
rect 43 35 45 37
<< ndifct0 >>
rect 9 18 11 20
rect 29 25 31 27
rect 29 18 31 20
rect 50 26 52 28
rect 39 17 41 19
<< ndifct1 >>
rect 19 26 21 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 9 57 11 59
rect 9 50 11 52
rect 29 57 31 59
rect 29 50 31 52
rect 49 57 51 59
<< pdifct1 >>
rect 19 52 21 54
rect 19 45 21 47
rect 39 52 41 54
rect 39 45 41 47
<< alu0 >>
rect 8 59 12 68
rect 8 57 9 59
rect 11 57 12 59
rect 8 52 12 57
rect 27 59 33 68
rect 27 57 29 59
rect 31 57 33 59
rect 8 50 9 52
rect 11 50 12 52
rect 8 48 12 50
rect 27 52 33 57
rect 48 59 52 68
rect 48 57 49 59
rect 51 57 52 59
rect 27 50 29 52
rect 31 50 33 52
rect 27 49 33 50
rect 48 55 52 57
rect 28 28 54 29
rect 28 27 50 28
rect 28 25 29 27
rect 31 26 50 27
rect 52 26 54 28
rect 31 25 54 26
rect 28 21 33 25
rect 7 20 33 21
rect 7 18 9 20
rect 11 18 29 20
rect 31 18 33 20
rect 7 17 33 18
rect 38 19 42 21
rect 38 17 39 19
rect 41 17 42 19
rect 38 12 42 17
<< labels >>
rlabel alu0 30 23 30 23 6 n1
rlabel alu0 20 19 20 19 6 n1
rlabel alu0 41 27 41 27 6 n1
rlabel alu1 4 32 4 32 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 40 20 40 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 44 36 44 6 z
rlabel alu1 28 44 28 44 6 z
rlabel alu1 28 74 28 74 6 vdd
rlabel polyct1 44 36 44 36 6 a
rlabel alu1 52 40 52 40 6 a
<< end >>
