magic
tech scmos
timestamp 1199202863
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 12 70 14 74
rect 19 70 21 74
rect 33 58 35 63
rect 12 39 14 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 11 22 13 33
rect 19 31 21 42
rect 33 39 35 42
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 19 29 25 31
rect 33 30 35 33
rect 19 27 21 29
rect 23 27 25 29
rect 19 25 25 27
rect 21 22 23 25
rect 33 17 35 22
rect 11 8 13 14
rect 21 8 23 14
<< ndif >>
rect 27 22 33 30
rect 35 28 42 30
rect 35 26 38 28
rect 40 26 42 28
rect 35 24 42 26
rect 35 22 40 24
rect 3 14 11 22
rect 13 20 21 22
rect 13 18 16 20
rect 18 18 21 20
rect 13 14 21 18
rect 23 19 31 22
rect 23 17 27 19
rect 29 17 31 19
rect 23 14 31 17
rect 3 11 9 14
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
<< pdif >>
rect 7 63 12 70
rect 5 61 12 63
rect 5 59 7 61
rect 9 59 12 61
rect 5 54 12 59
rect 5 52 7 54
rect 9 52 12 54
rect 5 50 12 52
rect 7 42 12 50
rect 14 42 19 70
rect 21 67 31 70
rect 21 65 27 67
rect 29 65 31 67
rect 21 58 31 65
rect 21 56 33 58
rect 21 54 27 56
rect 29 54 33 56
rect 21 42 33 54
rect 35 55 40 58
rect 35 53 42 55
rect 35 51 38 53
rect 40 51 42 53
rect 35 46 42 51
rect 35 44 38 46
rect 40 44 42 46
rect 35 42 42 44
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 6 61 14 63
rect 6 59 7 61
rect 9 59 14 61
rect 6 57 14 59
rect 6 55 11 57
rect 2 54 11 55
rect 2 52 7 54
rect 9 52 11 54
rect 2 51 11 52
rect 2 22 6 51
rect 18 47 22 55
rect 10 43 22 47
rect 10 37 14 43
rect 26 39 30 47
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 18 37 34 39
rect 18 35 31 37
rect 33 35 34 37
rect 18 33 34 35
rect 2 20 23 22
rect 2 18 16 20
rect 18 18 23 20
rect 2 17 23 18
rect -2 11 50 12
rect -2 9 5 11
rect 7 9 50 11
rect -2 1 50 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 33 22 35 30
rect 11 14 13 22
rect 21 14 23 22
<< pmos >>
rect 12 42 14 70
rect 19 42 21 70
rect 33 42 35 58
<< polyct0 >>
rect 21 27 23 29
<< polyct1 >>
rect 11 35 13 37
rect 31 35 33 37
<< ndifct0 >>
rect 38 26 40 28
rect 27 17 29 19
<< ndifct1 >>
rect 16 18 18 20
rect 5 9 7 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 27 65 29 67
rect 27 54 29 56
rect 38 51 40 53
rect 38 44 40 46
<< pdifct1 >>
rect 7 59 9 61
rect 7 52 9 54
<< alu0 >>
rect 26 67 30 68
rect 26 65 27 67
rect 29 65 30 67
rect 26 56 30 65
rect 26 54 27 56
rect 29 54 30 56
rect 26 52 30 54
rect 37 53 42 55
rect 37 51 38 53
rect 40 51 42 53
rect 37 46 42 51
rect 37 44 38 46
rect 40 44 42 46
rect 37 42 42 44
rect 19 29 25 30
rect 38 29 42 42
rect 19 27 21 29
rect 23 28 42 29
rect 23 27 38 28
rect 19 26 38 27
rect 40 26 42 28
rect 19 25 42 26
rect 26 19 30 21
rect 26 17 27 19
rect 29 17 30 19
rect 26 12 30 17
<< labels >>
rlabel alu0 30 27 30 27 6 an
rlabel alu0 39 48 39 48 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 36 20 36 6 a
rlabel alu1 12 40 12 40 6 b
rlabel alu1 20 52 20 52 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 40 28 40 6 a
rlabel alu1 24 74 24 74 6 vdd
<< end >>
