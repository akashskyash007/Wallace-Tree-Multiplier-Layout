magic
tech scmos
timestamp 1199202817
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 10 62 12 67
rect 20 62 22 67
rect 30 62 32 67
rect 40 62 42 67
rect 50 62 52 67
rect 60 62 62 67
rect 70 62 72 67
rect 80 62 82 67
rect 90 62 92 67
rect 10 39 12 42
rect 20 39 22 42
rect 30 39 32 42
rect 10 37 32 39
rect 10 35 12 37
rect 14 35 19 37
rect 21 35 32 37
rect 10 33 32 35
rect 10 30 12 33
rect 20 30 22 33
rect 30 30 32 33
rect 40 39 42 42
rect 50 39 52 42
rect 60 39 62 42
rect 40 37 62 39
rect 40 35 43 37
rect 45 35 51 37
rect 53 35 62 37
rect 40 33 62 35
rect 40 30 42 33
rect 50 30 52 33
rect 60 30 62 33
rect 70 39 72 42
rect 80 39 82 42
rect 90 39 92 42
rect 70 37 103 39
rect 70 35 99 37
rect 101 35 103 37
rect 70 33 103 35
rect 70 30 72 33
rect 80 30 82 33
rect 90 30 92 33
rect 101 30 103 33
rect 90 15 92 20
rect 101 15 103 20
rect 10 6 12 10
rect 20 6 22 10
rect 30 6 32 10
rect 40 6 42 10
rect 50 6 52 10
rect 60 6 62 10
rect 70 6 72 10
rect 80 6 82 10
<< ndif >>
rect 2 21 10 30
rect 2 19 4 21
rect 6 19 10 21
rect 2 14 10 19
rect 2 12 4 14
rect 6 12 10 14
rect 2 10 10 12
rect 12 28 20 30
rect 12 26 15 28
rect 17 26 20 28
rect 12 21 20 26
rect 12 19 15 21
rect 17 19 20 21
rect 12 10 20 19
rect 22 14 30 30
rect 22 12 25 14
rect 27 12 30 14
rect 22 10 30 12
rect 32 21 40 30
rect 32 19 35 21
rect 37 19 40 21
rect 32 10 40 19
rect 42 28 50 30
rect 42 26 45 28
rect 47 26 50 28
rect 42 10 50 26
rect 52 21 60 30
rect 52 19 55 21
rect 57 19 60 21
rect 52 10 60 19
rect 62 28 70 30
rect 62 26 65 28
rect 67 26 70 28
rect 62 21 70 26
rect 62 19 65 21
rect 67 19 70 21
rect 62 10 70 19
rect 72 28 80 30
rect 72 26 75 28
rect 77 26 80 28
rect 72 10 80 26
rect 82 24 90 30
rect 82 22 85 24
rect 87 22 90 24
rect 82 20 90 22
rect 92 28 101 30
rect 92 26 95 28
rect 97 26 101 28
rect 92 20 101 26
rect 103 26 108 30
rect 103 24 110 26
rect 103 22 106 24
rect 108 22 110 24
rect 103 20 110 22
rect 82 10 87 20
<< pdif >>
rect 2 60 10 62
rect 2 58 4 60
rect 6 58 10 60
rect 2 53 10 58
rect 2 51 4 53
rect 6 51 10 53
rect 2 42 10 51
rect 12 53 20 62
rect 12 51 15 53
rect 17 51 20 53
rect 12 46 20 51
rect 12 44 15 46
rect 17 44 20 46
rect 12 42 20 44
rect 22 60 30 62
rect 22 58 25 60
rect 27 58 30 60
rect 22 53 30 58
rect 22 51 25 53
rect 27 51 30 53
rect 22 42 30 51
rect 32 53 40 62
rect 32 51 35 53
rect 37 51 40 53
rect 32 46 40 51
rect 32 44 35 46
rect 37 44 40 46
rect 32 42 40 44
rect 42 60 50 62
rect 42 58 45 60
rect 47 58 50 60
rect 42 53 50 58
rect 42 51 45 53
rect 47 51 50 53
rect 42 42 50 51
rect 52 53 60 62
rect 52 51 55 53
rect 57 51 60 53
rect 52 46 60 51
rect 52 44 55 46
rect 57 44 60 46
rect 52 42 60 44
rect 62 60 70 62
rect 62 58 65 60
rect 67 58 70 60
rect 62 53 70 58
rect 62 51 65 53
rect 67 51 70 53
rect 62 42 70 51
rect 72 53 80 62
rect 72 51 75 53
rect 77 51 80 53
rect 72 46 80 51
rect 72 44 75 46
rect 77 44 80 46
rect 72 42 80 44
rect 82 60 90 62
rect 82 58 85 60
rect 87 58 90 60
rect 82 53 90 58
rect 82 51 85 53
rect 87 51 90 53
rect 82 42 90 51
rect 92 55 97 62
rect 92 53 99 55
rect 92 51 95 53
rect 97 51 99 53
rect 92 46 99 51
rect 92 44 95 46
rect 97 44 99 46
rect 92 42 99 44
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 68 114 79
rect 14 53 18 55
rect 14 51 15 53
rect 17 51 18 53
rect 2 38 6 47
rect 14 46 18 51
rect 34 53 38 55
rect 34 51 35 53
rect 37 51 38 53
rect 34 46 38 51
rect 54 53 58 55
rect 54 51 55 53
rect 57 51 58 53
rect 54 46 58 51
rect 74 53 78 63
rect 74 51 75 53
rect 77 51 78 53
rect 74 46 78 51
rect 90 46 96 47
rect 14 44 15 46
rect 17 44 35 46
rect 37 44 55 46
rect 57 44 75 46
rect 77 44 95 46
rect 14 43 96 44
rect 14 42 94 43
rect 74 41 94 42
rect 2 37 23 38
rect 2 35 12 37
rect 14 35 19 37
rect 21 35 23 37
rect 2 34 23 35
rect 33 37 55 38
rect 33 35 43 37
rect 45 35 51 37
rect 53 35 55 37
rect 33 34 55 35
rect 2 25 6 34
rect 33 26 39 34
rect 74 28 78 41
rect 74 26 75 28
rect 77 26 78 28
rect 106 39 110 55
rect 98 37 110 39
rect 98 35 99 37
rect 101 35 110 37
rect 98 33 110 35
rect 74 24 78 26
rect -2 1 114 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 10 10 12 30
rect 20 10 22 30
rect 30 10 32 30
rect 40 10 42 30
rect 50 10 52 30
rect 60 10 62 30
rect 70 10 72 30
rect 80 10 82 30
rect 90 20 92 30
rect 101 20 103 30
<< pmos >>
rect 10 42 12 62
rect 20 42 22 62
rect 30 42 32 62
rect 40 42 42 62
rect 50 42 52 62
rect 60 42 62 62
rect 70 42 72 62
rect 80 42 82 62
rect 90 42 92 62
<< polyct1 >>
rect 12 35 14 37
rect 19 35 21 37
rect 43 35 45 37
rect 51 35 53 37
rect 99 35 101 37
<< ndifct0 >>
rect 4 19 6 21
rect 4 12 6 14
rect 15 26 17 28
rect 15 19 17 21
rect 25 12 27 14
rect 35 19 37 21
rect 45 26 47 28
rect 55 19 57 21
rect 65 26 67 28
rect 65 19 67 21
rect 85 22 87 24
rect 95 26 97 28
rect 106 22 108 24
<< ndifct1 >>
rect 75 26 77 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 4 58 6 60
rect 4 51 6 53
rect 25 58 27 60
rect 25 51 27 53
rect 45 58 47 60
rect 45 51 47 53
rect 65 58 67 60
rect 65 51 67 53
rect 85 58 87 60
rect 85 51 87 53
rect 95 51 97 53
rect 96 44 97 46
<< pdifct1 >>
rect 15 51 17 53
rect 15 44 17 46
rect 35 51 37 53
rect 35 44 37 46
rect 55 51 57 53
rect 55 44 57 46
rect 75 51 77 53
rect 75 44 77 46
rect 95 44 96 46
<< alu0 >>
rect 2 60 8 68
rect 2 58 4 60
rect 6 58 8 60
rect 2 53 8 58
rect 23 60 29 68
rect 23 58 25 60
rect 27 58 29 60
rect 2 51 4 53
rect 6 51 8 53
rect 2 50 8 51
rect 23 53 29 58
rect 43 60 49 68
rect 43 58 45 60
rect 47 58 49 60
rect 23 51 25 53
rect 27 51 29 53
rect 23 50 29 51
rect 43 53 49 58
rect 63 60 69 68
rect 63 58 65 60
rect 67 58 69 60
rect 43 51 45 53
rect 47 51 49 53
rect 43 50 49 51
rect 63 53 69 58
rect 63 51 65 53
rect 67 51 69 53
rect 63 50 69 51
rect 83 60 89 68
rect 83 58 85 60
rect 87 58 89 60
rect 83 53 89 58
rect 83 51 85 53
rect 87 51 89 53
rect 83 50 89 51
rect 94 53 98 55
rect 94 51 95 53
rect 97 51 98 53
rect 94 47 98 51
rect 96 46 98 47
rect 97 44 98 46
rect 96 43 98 44
rect 94 42 98 43
rect 94 41 95 42
rect 13 28 18 30
rect 13 26 15 28
rect 17 26 18 28
rect 43 28 69 29
rect 43 26 45 28
rect 47 26 65 28
rect 67 26 69 28
rect 13 22 18 26
rect 43 25 69 26
rect 2 21 8 22
rect 2 19 4 21
rect 6 19 8 21
rect 2 14 8 19
rect 13 21 59 22
rect 13 19 15 21
rect 17 19 35 21
rect 37 19 55 21
rect 57 19 59 21
rect 13 18 59 19
rect 64 21 69 25
rect 91 29 95 41
rect 91 28 99 29
rect 91 26 95 28
rect 97 26 99 28
rect 84 24 88 26
rect 91 25 99 26
rect 84 22 85 24
rect 87 22 88 24
rect 84 21 88 22
rect 105 24 109 26
rect 105 22 106 24
rect 108 22 109 24
rect 105 21 109 22
rect 64 19 65 21
rect 67 19 109 21
rect 64 17 109 19
rect 2 12 4 14
rect 6 12 8 14
rect 23 14 29 15
rect 23 12 25 14
rect 27 12 29 14
<< labels >>
rlabel alu0 15 24 15 24 6 n1
rlabel alu0 66 23 66 23 6 n2
rlabel ndifct0 36 20 36 20 6 n1
rlabel alu0 56 27 56 27 6 n2
rlabel alu0 107 21 107 21 6 n2
rlabel alu0 86 21 86 21 6 n2
rlabel polyct1 20 36 20 36 6 a
rlabel alu1 12 36 12 36 6 a
rlabel alu1 4 36 4 36 6 a
rlabel alu1 20 44 20 44 6 z
rlabel polyct1 52 36 52 36 6 b
rlabel polyct1 44 36 44 36 6 b
rlabel alu1 36 32 36 32 6 b
rlabel alu1 44 44 44 44 6 z
rlabel alu1 52 44 52 44 6 z
rlabel alu1 28 44 28 44 6 z
rlabel alu1 36 48 36 48 6 z
rlabel alu1 56 6 56 6 6 vss
rlabel alu1 68 44 68 44 6 z
rlabel alu1 76 44 76 44 6 z
rlabel alu1 60 44 60 44 6 z
rlabel alu1 56 74 56 74 6 vdd
rlabel polyct1 100 36 100 36 6 c
rlabel alu1 92 44 92 44 6 z
rlabel alu1 108 44 108 44 6 c
rlabel alu1 84 44 84 44 6 z
<< end >>
