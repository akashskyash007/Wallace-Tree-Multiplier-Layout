magic
tech scmos
timestamp 1199973099
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -5 40 69 97
<< pwell >>
rect -5 -9 69 40
<< poly >>
rect 2 81 11 83
rect 2 79 7 81
rect 9 79 11 81
rect 2 77 11 79
rect 9 74 11 77
rect 21 81 30 83
rect 21 79 23 81
rect 25 79 30 81
rect 21 77 30 79
rect 34 81 43 83
rect 34 79 39 81
rect 41 79 43 81
rect 34 77 43 79
rect 21 74 23 77
rect 41 74 43 77
rect 53 81 62 83
rect 53 79 55 81
rect 57 79 62 81
rect 53 77 62 79
rect 53 74 55 77
rect 9 43 11 46
rect 21 43 23 46
rect 41 43 43 46
rect 53 43 55 46
rect 2 37 14 43
rect 18 37 30 43
rect 34 37 46 43
rect 50 37 62 43
rect 9 34 11 37
rect 21 34 23 37
rect 41 34 43 37
rect 53 34 55 37
rect 9 11 11 14
rect 2 5 11 11
rect 21 11 23 14
rect 41 11 43 14
rect 21 5 30 11
rect 34 5 43 11
rect 53 11 55 14
rect 53 5 62 11
<< ndif >>
rect 2 14 9 34
rect 11 14 21 34
rect 23 14 30 34
rect 34 14 41 34
rect 43 14 53 34
rect 55 14 62 34
rect 13 9 19 14
rect 13 7 15 9
rect 17 7 19 9
rect 13 2 19 7
rect 45 9 51 14
rect 45 7 47 9
rect 49 7 51 9
rect 45 2 51 7
<< pdif >>
rect 13 81 19 86
rect 13 79 15 81
rect 17 79 19 81
rect 13 74 19 79
rect 45 81 51 86
rect 45 79 47 81
rect 49 79 51 81
rect 45 74 51 79
rect 2 46 9 74
rect 11 46 21 74
rect 23 46 30 74
rect 34 46 41 74
rect 43 46 53 74
rect 55 46 62 74
<< alu1 >>
rect -2 89 66 90
rect -2 87 3 89
rect 5 87 7 89
rect 9 87 23 89
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 41 87 55 89
rect 57 87 59 89
rect 61 87 66 89
rect -2 86 66 87
rect 5 81 59 82
rect 5 79 7 81
rect 9 79 15 81
rect 17 79 23 81
rect 25 79 39 81
rect 41 79 47 81
rect 49 79 55 81
rect 57 79 59 81
rect 5 78 59 79
rect 13 9 51 10
rect 13 7 15 9
rect 17 7 47 9
rect 49 7 51 9
rect 13 6 51 7
rect -2 1 66 2
rect -2 -1 3 1
rect 5 -1 7 1
rect 9 -1 23 1
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 41 -1 55 1
rect 57 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< alu2 >>
rect -2 89 66 90
rect -2 87 7 89
rect 9 87 23 89
rect 25 87 39 89
rect 41 87 55 89
rect 57 87 66 89
rect -2 81 66 87
rect -2 79 7 81
rect 9 79 15 81
rect 17 79 23 81
rect 25 79 39 81
rect 41 79 47 81
rect 49 79 55 81
rect 57 79 66 81
rect -2 76 66 79
rect -2 9 66 12
rect -2 7 15 9
rect 17 7 47 9
rect 49 7 66 9
rect -2 1 66 7
rect -2 -1 7 1
rect 9 -1 23 1
rect 25 -1 39 1
rect 41 -1 55 1
rect 57 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 7 3
rect 0 -1 3 1
rect 5 -1 7 1
rect 0 -3 7 -1
rect 25 1 39 3
rect 25 -1 27 1
rect 29 -1 35 1
rect 37 -1 39 1
rect 25 -3 39 -1
rect 57 1 64 3
rect 57 -1 59 1
rect 61 -1 64 1
rect 57 -3 64 -1
<< ntie >>
rect 0 89 7 91
rect 0 87 3 89
rect 5 87 7 89
rect 0 85 7 87
rect 25 89 39 91
rect 25 87 27 89
rect 29 87 35 89
rect 37 87 39 89
rect 25 85 39 87
rect 57 89 64 91
rect 57 87 59 89
rect 61 87 64 89
rect 57 85 64 87
<< nmos >>
rect 9 14 11 34
rect 21 14 23 34
rect 41 14 43 34
rect 53 14 55 34
<< pmos >>
rect 9 46 11 74
rect 21 46 23 74
rect 41 46 43 74
rect 53 46 55 74
<< polyct1 >>
rect 7 79 9 81
rect 23 79 25 81
rect 39 79 41 81
rect 55 79 57 81
<< ndifct1 >>
rect 15 7 17 9
rect 47 7 49 9
<< ntiect1 >>
rect 3 87 5 89
rect 27 87 29 89
rect 35 87 37 89
rect 59 87 61 89
<< ptiect1 >>
rect 3 -1 5 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 59 -1 61 1
<< pdifct1 >>
rect 15 79 17 81
rect 47 79 49 81
<< via1 >>
rect 7 87 9 89
rect 23 87 25 89
rect 39 87 41 89
rect 55 87 57 89
rect 7 79 9 81
rect 15 79 17 81
rect 23 79 25 81
rect 39 79 41 81
rect 47 79 49 81
rect 55 79 57 81
rect 15 7 17 9
rect 47 7 49 9
rect 7 -1 9 1
rect 23 -1 25 1
rect 39 -1 41 1
rect 55 -1 57 1
<< labels >>
rlabel alu2 32 6 32 6 6 vss
rlabel alu2 32 82 32 82 6 vdd
<< end >>
