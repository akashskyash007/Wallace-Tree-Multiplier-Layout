magic
tech scmos
timestamp 1199203410
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 9 70 11 74
rect 27 70 29 74
rect 37 70 39 74
rect 44 70 46 74
rect 57 70 59 74
rect 67 70 69 74
rect 9 39 11 42
rect 27 39 29 42
rect 9 37 29 39
rect 9 35 11 37
rect 13 35 15 37
rect 37 35 39 42
rect 44 39 46 42
rect 57 39 59 42
rect 9 33 15 35
rect 33 33 39 35
rect 43 37 49 39
rect 43 35 45 37
rect 47 35 49 37
rect 57 37 63 39
rect 57 35 59 37
rect 61 35 63 37
rect 43 33 52 35
rect 57 33 63 35
rect 67 36 69 42
rect 67 34 73 36
rect 11 26 13 33
rect 33 31 35 33
rect 37 31 39 33
rect 21 29 39 31
rect 21 26 23 29
rect 50 27 52 33
rect 60 27 62 33
rect 67 32 69 34
rect 71 32 73 34
rect 67 30 73 32
rect 67 27 69 30
rect 11 8 13 13
rect 21 8 23 13
rect 50 6 52 10
rect 60 6 62 10
rect 67 6 69 10
<< ndif >>
rect 4 17 11 26
rect 4 15 6 17
rect 8 15 11 17
rect 4 13 11 15
rect 13 24 21 26
rect 13 22 16 24
rect 18 22 21 24
rect 13 13 21 22
rect 23 24 31 26
rect 23 22 27 24
rect 29 22 31 24
rect 45 23 50 27
rect 23 20 31 22
rect 42 21 50 23
rect 23 13 28 20
rect 42 19 44 21
rect 46 19 50 21
rect 42 17 50 19
rect 45 10 50 17
rect 52 25 60 27
rect 52 23 55 25
rect 57 23 60 25
rect 52 10 60 23
rect 62 10 67 27
rect 69 14 76 27
rect 69 12 72 14
rect 74 12 76 14
rect 69 10 76 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 48 16 70
rect 22 63 27 70
rect 20 61 27 63
rect 20 59 22 61
rect 24 59 27 61
rect 20 57 27 59
rect 11 46 18 48
rect 11 44 14 46
rect 16 44 18 46
rect 11 42 18 44
rect 22 42 27 57
rect 29 46 37 70
rect 29 44 32 46
rect 34 44 37 46
rect 29 42 37 44
rect 39 42 44 70
rect 46 68 57 70
rect 46 66 50 68
rect 52 66 57 68
rect 46 42 57 66
rect 59 61 67 70
rect 59 59 62 61
rect 64 59 67 61
rect 59 54 67 59
rect 59 52 62 54
rect 64 52 67 54
rect 59 42 67 52
rect 69 68 77 70
rect 69 66 72 68
rect 74 66 77 68
rect 69 61 77 66
rect 69 59 72 61
rect 74 59 77 61
rect 69 42 77 59
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 2 39 6 47
rect 2 37 14 39
rect 2 35 11 37
rect 13 35 14 37
rect 2 33 14 35
rect 2 25 6 33
rect 26 26 30 46
rect 58 41 78 47
rect 58 37 62 41
rect 58 35 59 37
rect 61 35 62 37
rect 58 33 62 35
rect 66 29 78 31
rect 65 25 78 29
rect 34 18 38 22
rect 42 21 46 22
rect 42 19 44 21
rect 42 18 46 19
rect 65 18 71 25
rect -2 1 82 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 11 13 13 26
rect 21 13 23 26
rect 50 10 52 27
rect 60 10 62 27
rect 67 10 69 27
<< pmos >>
rect 9 42 11 70
rect 27 42 29 70
rect 37 42 39 70
rect 44 42 46 70
rect 57 42 59 70
rect 67 42 69 70
<< polyct0 >>
rect 45 35 47 37
rect 35 31 37 33
rect 69 32 71 34
<< polyct1 >>
rect 11 35 13 37
rect 59 35 61 37
<< ndifct0 >>
rect 6 15 8 17
rect 16 22 18 24
rect 27 22 29 24
rect 55 23 57 25
rect 72 12 74 14
<< ndifct1 >>
rect 44 19 46 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 22 59 24 61
rect 14 44 16 46
rect 32 44 34 46
rect 50 66 52 68
rect 62 59 64 61
rect 62 52 64 54
rect 72 66 74 68
rect 72 59 74 61
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 48 66 50 68
rect 52 66 54 68
rect 48 65 54 66
rect 70 66 72 68
rect 74 66 76 68
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 20 61 55 62
rect 20 59 22 61
rect 24 59 55 61
rect 20 58 55 59
rect 51 55 55 58
rect 61 61 66 63
rect 61 59 62 61
rect 64 59 66 61
rect 61 55 66 59
rect 70 61 76 66
rect 70 59 72 61
rect 74 59 76 61
rect 70 58 76 59
rect 51 54 66 55
rect 18 50 46 54
rect 18 47 22 50
rect 12 46 22 47
rect 12 44 14 46
rect 16 44 22 46
rect 12 43 22 44
rect 18 25 22 43
rect 14 24 22 25
rect 14 22 16 24
rect 18 22 22 24
rect 14 21 22 22
rect 26 46 36 47
rect 30 44 32 46
rect 34 44 36 46
rect 30 43 36 44
rect 42 39 46 50
rect 51 52 62 54
rect 64 52 66 54
rect 51 51 66 52
rect 42 37 48 39
rect 42 35 45 37
rect 47 35 48 37
rect 34 33 38 35
rect 42 33 48 35
rect 34 31 35 33
rect 37 31 38 33
rect 34 30 38 31
rect 51 30 55 51
rect 68 34 72 36
rect 68 32 69 34
rect 71 32 72 34
rect 68 31 72 32
rect 34 26 55 30
rect 26 24 30 26
rect 26 22 27 24
rect 29 22 30 24
rect 51 25 59 26
rect 51 23 55 25
rect 57 23 59 25
rect 51 22 59 23
rect 5 17 9 19
rect 26 18 34 22
rect 38 18 42 22
rect 46 18 48 22
rect 5 15 6 17
rect 8 15 9 17
rect 5 12 9 15
rect 70 14 76 15
rect 70 12 72 14
rect 74 12 76 14
<< labels >>
rlabel alu0 36 30 36 30 6 an
rlabel alu0 20 37 20 37 6 bn
rlabel alu0 17 45 17 45 6 bn
rlabel alu0 45 36 45 36 6 bn
rlabel alu0 37 60 37 60 6 an
rlabel alu0 53 42 53 42 6 an
rlabel alu0 63 57 63 57 6 an
rlabel alu1 4 36 4 36 6 b
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 36 28 36 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 76 28 76 28 6 a1
rlabel alu1 68 24 68 24 6 a1
rlabel alu1 68 44 68 44 6 a2
rlabel alu1 76 44 76 44 6 a2
rlabel alu1 60 40 60 40 6 a2
<< end >>
