magic
tech scmos
timestamp 1199980699
<< ab >>
rect 0 0 32 88
<< nwell >>
rect -8 40 40 97
<< pwell >>
rect -8 -9 40 40
<< poly >>
rect 5 84 14 86
rect 5 82 7 84
rect 9 82 14 84
rect 5 80 14 82
rect 18 84 27 86
rect 18 82 23 84
rect 25 82 27 84
rect 18 80 27 82
rect 9 77 11 80
rect 21 77 23 80
rect 9 48 11 51
rect 21 48 23 51
rect 2 42 11 48
rect 15 42 30 48
rect 2 32 17 38
rect 21 32 30 38
rect 9 29 11 32
rect 21 29 23 32
rect 9 8 11 11
rect 21 8 23 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 6 27 8
rect 18 4 23 6
rect 25 4 27 6
rect 18 2 27 4
<< ndif >>
rect 2 11 9 29
rect 11 11 21 29
rect 23 11 30 29
<< pdif >>
rect 2 51 9 77
rect 11 51 21 77
rect 23 51 30 77
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect -2 83 -1 85
rect 1 84 31 85
rect 1 83 7 84
rect -2 82 7 83
rect 9 82 23 84
rect 25 83 31 84
rect 33 83 34 85
rect 25 82 34 83
rect -2 81 34 82
rect -2 6 34 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 4 23 6
rect 25 5 34 6
rect 25 4 31 5
rect 1 3 31 4
rect 33 3 34 5
rect -2 -2 2 3
rect 30 -2 34 3
<< alu2 >>
rect -2 85 34 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 80 34 83
rect -2 5 34 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 34 5
rect -2 -2 34 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
<< polyct1 >>
rect 7 82 9 84
rect 23 82 25 84
rect 7 4 9 6
rect 23 4 25 6
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect -1 3 1 5
rect 31 3 33 5
<< labels >>
rlabel alu2 16 4 16 4 6 vss
rlabel alu2 16 84 16 84 6 vdd
<< end >>
