magic
tech scmos
timestamp 1199201643
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 9 35 11 38
rect 19 35 21 47
rect 29 43 31 47
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 29 37 35 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 9 26 11 29
rect 22 26 24 29
rect 29 26 31 37
rect 9 7 11 12
rect 22 8 24 13
rect 29 8 31 13
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 16 9 22
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 13 22 26
rect 24 13 29 26
rect 31 19 36 26
rect 31 17 38 19
rect 31 15 34 17
rect 36 15 38 17
rect 31 13 38 15
rect 11 12 20 13
rect 13 7 20 12
rect 13 5 15 7
rect 17 5 20 7
rect 13 3 20 5
<< pdif >>
rect 4 59 9 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 4 38 9 46
rect 11 64 19 66
rect 11 62 14 64
rect 16 62 19 64
rect 11 57 19 62
rect 11 55 14 57
rect 16 55 19 57
rect 11 47 19 55
rect 21 58 29 66
rect 21 56 24 58
rect 26 56 29 58
rect 21 51 29 56
rect 21 49 24 51
rect 26 49 29 51
rect 21 47 29 49
rect 31 64 38 66
rect 31 62 34 64
rect 36 62 38 64
rect 31 57 38 62
rect 31 55 34 57
rect 36 55 38 57
rect 31 47 38 55
rect 11 38 17 47
<< alu1 >>
rect -2 64 42 72
rect 2 57 7 59
rect 2 55 4 57
rect 6 55 7 57
rect 2 50 7 55
rect 2 48 4 50
rect 6 48 7 50
rect 2 46 7 48
rect 2 24 6 46
rect 34 42 38 51
rect 25 41 38 42
rect 25 39 31 41
rect 33 39 38 41
rect 25 38 38 39
rect 17 33 31 34
rect 17 31 21 33
rect 23 31 31 33
rect 17 30 31 31
rect 2 22 4 24
rect 2 19 6 22
rect 2 16 14 19
rect 2 14 4 16
rect 6 14 14 16
rect 26 21 31 30
rect 2 13 14 14
rect -2 7 42 8
rect -2 5 15 7
rect 17 5 42 7
rect -2 0 42 5
<< nmos >>
rect 9 12 11 26
rect 22 13 24 26
rect 29 13 31 26
<< pmos >>
rect 9 38 11 66
rect 19 47 21 66
rect 29 47 31 66
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 31 39 33 41
rect 21 31 23 33
<< ndifct0 >>
rect 34 15 36 17
<< ndifct1 >>
rect 4 22 6 24
rect 4 14 6 16
rect 15 5 17 7
<< pdifct0 >>
rect 14 62 16 64
rect 14 55 16 57
rect 24 56 26 58
rect 24 49 26 51
rect 34 62 36 64
rect 34 55 36 57
<< pdifct1 >>
rect 4 55 6 57
rect 4 48 6 50
<< alu0 >>
rect 12 62 14 64
rect 16 62 18 64
rect 12 57 18 62
rect 32 62 34 64
rect 36 62 38 64
rect 12 55 14 57
rect 16 55 18 57
rect 12 54 18 55
rect 22 58 28 59
rect 22 56 24 58
rect 26 56 28 58
rect 22 51 28 56
rect 32 57 38 62
rect 32 55 34 57
rect 36 55 38 57
rect 32 54 38 55
rect 22 50 24 51
rect 14 49 24 50
rect 26 49 28 51
rect 14 46 28 49
rect 14 42 18 46
rect 10 38 18 42
rect 10 33 14 38
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 6 19 7 26
rect 10 22 22 26
rect 18 18 22 22
rect 18 17 38 18
rect 18 15 34 17
rect 36 15 38 17
rect 18 14 38 15
<< labels >>
rlabel polyct0 12 32 12 32 6 zn
rlabel alu0 28 16 28 16 6 zn
rlabel alu0 25 52 25 52 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 20 32 20 32 6 a
rlabel alu1 28 28 28 28 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 36 48 36 48 6 b
<< end >>
