magic
tech scmos
timestamp 1199203546
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 19 66 21 70
rect 29 66 31 70
rect 36 66 38 70
rect 9 59 11 64
rect 69 54 71 59
rect 52 48 58 50
rect 52 46 54 48
rect 56 46 58 48
rect 9 40 11 43
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 19 35 21 43
rect 10 19 12 34
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 29 34 31 43
rect 36 40 38 43
rect 52 40 58 46
rect 36 38 58 40
rect 29 32 48 34
rect 19 29 25 31
rect 37 30 44 32
rect 46 30 48 32
rect 19 25 21 29
rect 17 22 21 25
rect 37 28 48 30
rect 56 31 58 38
rect 69 35 71 38
rect 65 33 71 35
rect 65 31 67 33
rect 69 31 71 33
rect 56 28 59 31
rect 65 29 71 31
rect 17 19 19 22
rect 27 19 29 24
rect 37 19 39 28
rect 57 25 59 28
rect 69 20 71 29
rect 57 14 59 18
rect 10 7 12 12
rect 17 7 19 12
rect 27 4 29 12
rect 37 8 39 12
rect 69 4 71 13
rect 27 2 71 4
<< ndif >>
rect 50 22 57 25
rect 50 20 52 22
rect 54 20 57 22
rect 2 12 10 19
rect 12 12 17 19
rect 19 17 27 19
rect 19 15 22 17
rect 24 15 27 17
rect 19 12 27 15
rect 29 17 37 19
rect 29 15 32 17
rect 34 15 37 17
rect 29 12 37 15
rect 39 16 46 19
rect 50 18 57 20
rect 59 20 67 25
rect 59 18 69 20
rect 39 14 42 16
rect 44 14 46 16
rect 61 17 69 18
rect 61 15 63 17
rect 65 15 69 17
rect 39 12 46 14
rect 61 13 69 15
rect 71 18 78 20
rect 71 16 74 18
rect 76 16 78 18
rect 71 13 78 16
rect 2 7 8 12
rect 2 5 4 7
rect 6 5 8 7
rect 2 3 8 5
<< pdif >>
rect 14 59 19 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 53 9 55
rect 4 43 9 53
rect 11 49 19 59
rect 11 47 14 49
rect 16 47 19 49
rect 11 43 19 47
rect 21 47 29 66
rect 21 45 24 47
rect 26 45 29 47
rect 21 43 29 45
rect 31 43 36 66
rect 38 64 47 66
rect 38 62 41 64
rect 43 62 47 64
rect 38 43 47 62
rect 61 67 67 69
rect 61 65 63 67
rect 65 65 67 67
rect 61 54 67 65
rect 61 38 69 54
rect 71 51 76 54
rect 71 49 78 51
rect 71 47 74 49
rect 76 47 78 49
rect 71 42 78 47
rect 71 40 74 42
rect 76 40 78 42
rect 71 38 78 40
<< alu1 >>
rect -2 67 82 72
rect -2 65 53 67
rect 55 65 63 67
rect 65 65 73 67
rect 75 65 82 67
rect -2 64 82 65
rect 2 49 18 50
rect 2 47 14 49
rect 16 47 18 49
rect 2 46 18 47
rect 2 18 6 46
rect 42 35 46 51
rect 50 48 62 51
rect 50 46 54 48
rect 56 46 62 48
rect 50 45 62 46
rect 58 37 62 45
rect 42 32 54 35
rect 42 30 44 32
rect 46 30 54 32
rect 42 29 54 30
rect 66 33 70 43
rect 66 31 67 33
rect 69 31 70 33
rect 66 27 70 31
rect 2 17 26 18
rect 2 15 22 17
rect 24 15 26 17
rect 2 14 26 15
rect 58 21 70 27
rect -2 7 82 8
rect -2 5 4 7
rect 6 5 82 7
rect -2 0 82 5
<< ptie >>
rect 50 10 56 12
rect 50 8 52 10
rect 54 8 56 10
rect 50 6 56 8
<< ntie >>
rect 51 67 57 69
rect 51 65 53 67
rect 55 65 57 67
rect 51 53 57 65
rect 71 67 77 69
rect 71 65 73 67
rect 75 65 77 67
rect 71 63 77 65
<< nmos >>
rect 10 12 12 19
rect 17 12 19 19
rect 27 12 29 19
rect 37 12 39 19
rect 57 18 59 25
rect 69 13 71 20
<< pmos >>
rect 9 43 11 59
rect 19 43 21 66
rect 29 43 31 66
rect 36 43 38 66
rect 69 38 71 54
<< polyct0 >>
rect 11 36 13 38
rect 21 31 23 33
<< polyct1 >>
rect 54 46 56 48
rect 44 30 46 32
rect 67 31 69 33
<< ndifct0 >>
rect 52 20 54 22
rect 32 15 34 17
rect 42 14 44 16
rect 63 15 65 17
rect 74 16 76 18
<< ndifct1 >>
rect 22 15 24 17
rect 4 5 6 7
<< ntiect1 >>
rect 53 65 55 67
rect 73 65 75 67
<< ptiect0 >>
rect 52 8 54 10
<< pdifct0 >>
rect 4 55 6 57
rect 24 45 26 47
rect 41 62 43 64
rect 74 47 76 49
rect 74 40 76 42
<< pdifct1 >>
rect 14 47 16 49
rect 63 65 65 67
<< alu0 >>
rect 39 62 41 64
rect 43 62 45 64
rect 39 61 45 62
rect 2 57 77 58
rect 2 55 4 57
rect 6 55 77 57
rect 2 54 77 55
rect 23 47 27 49
rect 23 45 24 47
rect 26 45 27 47
rect 23 42 27 45
rect 10 38 27 42
rect 10 36 11 38
rect 13 36 14 38
rect 10 26 14 36
rect 31 34 35 54
rect 19 33 35 34
rect 19 31 21 33
rect 23 31 35 33
rect 19 30 35 31
rect 73 49 77 54
rect 73 47 74 49
rect 76 47 77 49
rect 10 25 35 26
rect 10 22 55 25
rect 31 21 52 22
rect 31 17 35 21
rect 51 20 52 21
rect 54 20 55 22
rect 73 42 77 47
rect 73 40 74 42
rect 76 40 77 42
rect 51 18 55 20
rect 73 18 77 40
rect 61 17 67 18
rect 31 15 32 17
rect 34 15 35 17
rect 31 13 35 15
rect 40 16 46 17
rect 40 14 42 16
rect 44 14 46 16
rect 40 8 46 14
rect 61 15 63 17
rect 65 15 67 17
rect 51 10 55 12
rect 51 8 52 10
rect 54 8 55 10
rect 61 8 67 15
rect 73 16 74 18
rect 76 16 77 18
rect 73 14 77 16
<< labels >>
rlabel alu0 12 32 12 32 6 an
rlabel alu0 33 19 33 19 6 an
rlabel alu0 27 32 27 32 6 bn
rlabel alu0 25 43 25 43 6 an
rlabel alu0 43 23 43 23 6 an
rlabel alu0 39 56 39 56 6 bn
rlabel alu0 75 36 75 36 6 bn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 52 32 52 32 6 a2
rlabel alu1 44 40 44 40 6 a2
rlabel alu1 52 48 52 48 6 a1
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 60 24 60 24 6 b
rlabel polyct1 68 32 68 32 6 b
rlabel alu1 60 44 60 44 6 a1
<< end >>
