magic
tech scmos
timestamp 1199980651
<< ab >>
rect 0 0 96 88
<< nwell >>
rect -8 40 104 97
<< pwell >>
rect -8 -9 104 40
<< poly >>
rect 5 80 14 86
rect 18 80 27 86
rect 37 84 46 86
rect 37 82 42 84
rect 44 82 46 84
rect 37 80 46 82
rect 50 80 59 86
rect 69 80 78 86
rect 82 84 91 86
rect 82 82 87 84
rect 89 82 91 84
rect 82 80 91 82
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 73 77 75 80
rect 85 77 87 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 73 48 75 51
rect 85 48 87 51
rect 2 46 11 48
rect 2 44 7 46
rect 9 44 11 46
rect 2 42 11 44
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 39 46
rect 41 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 66 46 75 48
rect 66 44 71 46
rect 73 44 75 46
rect 66 42 75 44
rect 79 42 94 48
rect 2 36 17 38
rect 2 34 7 36
rect 9 34 17 36
rect 2 32 17 34
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 39 36
rect 41 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 66 36 81 38
rect 66 34 71 36
rect 73 34 81 36
rect 66 32 81 34
rect 85 32 94 38
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 73 29 75 32
rect 85 29 87 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 73 8 75 11
rect 85 8 87 11
rect 5 2 14 8
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
rect 69 2 78 8
rect 82 6 91 8
rect 82 4 87 6
rect 89 4 91 6
rect 82 2 91 4
<< ndif >>
rect 2 24 9 29
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 11 9 15
rect 11 15 21 29
rect 11 13 15 15
rect 17 13 21 15
rect 11 11 21 13
rect 23 17 30 29
rect 23 15 26 17
rect 28 15 30 17
rect 23 11 30 15
rect 34 25 41 29
rect 34 23 36 25
rect 38 23 41 25
rect 34 11 41 23
rect 43 25 53 29
rect 43 23 47 25
rect 49 23 53 25
rect 43 11 53 23
rect 55 25 62 29
rect 55 23 58 25
rect 60 23 62 25
rect 55 18 62 23
rect 55 16 58 18
rect 60 16 62 18
rect 55 11 62 16
rect 66 24 73 29
rect 66 22 68 24
rect 70 22 73 24
rect 66 17 73 22
rect 66 15 68 17
rect 70 15 73 17
rect 66 11 73 15
rect 75 16 85 29
rect 75 14 79 16
rect 81 14 85 16
rect 75 11 85 14
rect 87 11 94 29
<< pdif >>
rect 2 65 9 77
rect 2 63 4 65
rect 6 63 9 65
rect 2 58 9 63
rect 2 56 4 58
rect 6 56 9 58
rect 2 51 9 56
rect 11 73 21 77
rect 11 71 15 73
rect 17 71 21 73
rect 11 66 21 71
rect 11 64 15 66
rect 17 64 21 66
rect 11 51 21 64
rect 23 72 30 77
rect 23 70 26 72
rect 28 70 30 72
rect 23 65 30 70
rect 23 63 26 65
rect 28 63 30 65
rect 23 51 30 63
rect 34 73 41 77
rect 34 71 36 73
rect 38 71 41 73
rect 34 51 41 71
rect 43 57 53 77
rect 43 55 47 57
rect 49 55 53 57
rect 43 51 53 55
rect 55 65 62 77
rect 55 63 58 65
rect 60 63 62 65
rect 55 51 62 63
rect 66 72 73 77
rect 66 70 68 72
rect 70 70 73 72
rect 66 65 73 70
rect 66 63 68 65
rect 70 63 73 65
rect 66 58 73 63
rect 66 56 68 58
rect 70 56 73 58
rect 66 51 73 56
rect 75 73 85 77
rect 75 71 79 73
rect 81 71 85 73
rect 75 66 85 71
rect 75 64 79 66
rect 81 64 85 66
rect 75 51 85 64
rect 87 51 94 77
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect 62 85 66 90
rect 94 85 98 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 34 85
rect -2 81 34 83
rect 62 83 63 85
rect 65 84 95 85
rect 65 83 87 84
rect 62 82 87 83
rect 89 83 95 84
rect 97 83 98 85
rect 89 82 98 83
rect 62 81 98 82
rect 14 73 18 81
rect 14 71 15 73
rect 17 71 18 73
rect 14 66 18 71
rect 14 64 15 66
rect 17 64 18 66
rect 14 62 18 64
rect 46 57 50 59
rect 46 55 47 57
rect 49 55 50 57
rect 6 46 10 51
rect 6 44 7 46
rect 9 44 10 46
rect 6 36 10 44
rect 6 34 7 36
rect 9 34 10 36
rect 6 29 10 34
rect 22 46 26 51
rect 22 44 23 46
rect 25 44 26 46
rect 22 36 26 44
rect 22 34 23 36
rect 25 34 26 36
rect 22 29 26 34
rect 46 25 50 55
rect 54 50 58 59
rect 78 73 82 81
rect 78 71 79 73
rect 81 71 82 73
rect 78 66 82 71
rect 78 64 79 66
rect 81 64 82 66
rect 78 62 82 64
rect 54 46 74 50
rect 54 44 55 46
rect 57 44 58 46
rect 54 36 58 44
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 70 44 71 46
rect 73 44 74 46
rect 70 36 74 44
rect 70 34 71 36
rect 73 34 74 36
rect 70 32 74 34
rect 46 23 47 25
rect 49 23 50 25
rect 46 21 50 23
rect 14 15 18 17
rect 14 13 15 15
rect 17 13 18 15
rect 78 16 82 18
rect 78 14 79 16
rect 81 14 82 16
rect 14 7 18 13
rect 78 7 82 14
rect -2 5 34 7
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 34 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 6 98 7
rect 62 5 87 6
rect 62 3 63 5
rect 65 4 87 5
rect 89 5 98 6
rect 89 4 95 5
rect 65 3 95 4
rect 97 3 98 5
rect 62 -2 66 3
rect 94 -2 98 3
<< alu2 >>
rect -2 85 98 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 95 85
rect 97 83 98 85
rect -2 80 98 83
rect -2 5 98 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 95 5
rect 97 3 98 5
rect -2 -2 98 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
rect 93 5 99 7
rect 93 3 95 5
rect 97 3 99 5
rect 93 0 99 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
rect 93 85 99 88
rect 93 83 95 85
rect 97 83 99 85
rect 93 81 99 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
rect 73 11 75 29
rect 85 11 87 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
rect 73 51 75 77
rect 85 51 87 77
<< polyct0 >>
rect 42 82 44 84
rect 39 44 41 46
rect 39 34 41 36
<< polyct1 >>
rect 87 82 89 84
rect 7 44 9 46
rect 23 44 25 46
rect 55 44 57 46
rect 71 44 73 46
rect 7 34 9 36
rect 23 34 25 36
rect 55 34 57 36
rect 71 34 73 36
rect 87 4 89 6
<< ndifct0 >>
rect 4 22 6 24
rect 4 15 6 17
rect 26 15 28 17
rect 36 23 38 25
rect 58 23 60 25
rect 58 16 60 18
rect 68 22 70 24
rect 68 15 70 17
<< ndifct1 >>
rect 15 13 17 15
rect 47 23 49 25
rect 79 14 81 16
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< pdifct0 >>
rect 4 63 6 65
rect 4 56 6 58
rect 26 70 28 72
rect 26 63 28 65
rect 36 71 38 73
rect 58 63 60 65
rect 68 70 70 72
rect 68 63 70 65
rect 68 56 70 58
<< pdifct1 >>
rect 15 71 17 73
rect 15 64 17 66
rect 47 55 49 57
rect 79 71 81 73
rect 79 64 81 66
<< alu0 >>
rect 40 84 58 85
rect 40 82 42 84
rect 44 82 58 84
rect 40 81 58 82
rect 54 74 58 81
rect 3 65 7 67
rect 3 63 4 65
rect 6 63 7 65
rect 3 58 7 63
rect 25 73 40 74
rect 25 72 36 73
rect 25 70 26 72
rect 28 71 36 72
rect 38 71 40 73
rect 28 70 40 71
rect 54 72 71 74
rect 54 70 68 72
rect 70 70 71 72
rect 25 65 29 70
rect 25 63 26 65
rect 28 63 29 65
rect 25 61 29 63
rect 38 65 62 66
rect 38 63 58 65
rect 60 63 62 65
rect 38 62 62 63
rect 67 65 71 70
rect 67 63 68 65
rect 70 63 71 65
rect 38 58 42 62
rect 3 56 4 58
rect 6 56 42 58
rect 3 54 42 56
rect 38 46 42 48
rect 38 44 39 46
rect 41 44 42 46
rect 38 36 42 44
rect 38 34 39 36
rect 41 34 42 36
rect 38 32 42 34
rect 3 25 40 26
rect 3 24 36 25
rect 3 22 4 24
rect 6 23 36 24
rect 38 23 40 25
rect 6 22 40 23
rect 67 58 71 63
rect 67 56 68 58
rect 70 56 82 58
rect 67 54 82 56
rect 3 17 7 22
rect 57 25 61 27
rect 78 26 82 54
rect 57 23 58 25
rect 60 23 61 25
rect 57 18 61 23
rect 24 17 58 18
rect 3 15 4 17
rect 6 15 7 17
rect 3 13 7 15
rect 24 15 26 17
rect 28 16 58 17
rect 60 16 61 18
rect 28 15 61 16
rect 24 14 61 15
rect 67 24 82 26
rect 67 22 68 24
rect 70 22 82 24
rect 67 17 71 22
rect 67 15 68 17
rect 70 15 71 17
rect 67 13 71 15
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect 95 83 97 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
rect 95 3 97 5
<< labels >>
rlabel alu1 8 40 8 40 6 a1
rlabel alu1 24 40 24 40 6 a2
rlabel alu1 48 40 48 40 6 z
rlabel alu1 56 48 56 48 6 s
rlabel alu1 64 48 64 48 6 s
rlabel alu1 72 40 72 40 6 s
rlabel alu2 48 4 48 4 6 vss
rlabel alu2 48 84 48 84 6 vdd
<< end >>
