magic
tech scmos
timestamp 1199469777
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -5 48 55 105
<< pwell >>
rect -5 -5 55 48
<< poly >>
rect 13 94 15 98
rect 25 94 27 98
rect 37 85 39 90
rect 13 52 15 55
rect 25 52 27 55
rect 13 50 21 52
rect 13 49 17 50
rect 15 48 17 49
rect 19 48 21 50
rect 15 46 21 48
rect 25 50 32 52
rect 25 48 28 50
rect 30 48 32 50
rect 25 46 32 48
rect 17 39 19 46
rect 25 39 27 46
rect 37 42 39 55
rect 35 40 41 42
rect 35 38 37 40
rect 39 38 41 40
rect 35 36 41 38
rect 37 33 39 36
rect 37 13 39 18
rect 17 2 19 6
rect 25 2 27 6
<< ndif >>
rect 9 37 17 39
rect 9 35 11 37
rect 13 35 17 37
rect 9 29 17 35
rect 9 27 11 29
rect 13 27 17 29
rect 9 25 17 27
rect 12 6 17 25
rect 19 6 25 39
rect 27 33 32 39
rect 27 21 37 33
rect 27 19 31 21
rect 33 19 37 21
rect 27 18 37 19
rect 39 30 47 33
rect 39 28 43 30
rect 45 28 47 30
rect 39 22 47 28
rect 39 20 43 22
rect 45 20 47 22
rect 39 18 47 20
rect 27 11 35 18
rect 27 9 31 11
rect 33 9 35 11
rect 27 6 35 9
<< pdif >>
rect 4 92 13 94
rect 4 90 7 92
rect 9 90 13 92
rect 4 82 13 90
rect 4 80 7 82
rect 9 80 13 82
rect 4 55 13 80
rect 15 81 25 94
rect 15 79 19 81
rect 21 79 25 81
rect 15 71 25 79
rect 15 69 19 71
rect 21 69 25 71
rect 15 55 25 69
rect 27 92 35 94
rect 27 90 31 92
rect 33 90 35 92
rect 27 85 35 90
rect 27 82 37 85
rect 27 80 31 82
rect 33 80 37 82
rect 27 55 37 80
rect 39 69 44 85
rect 39 67 47 69
rect 39 65 43 67
rect 45 65 47 67
rect 39 59 47 65
rect 39 57 43 59
rect 45 57 47 59
rect 39 55 47 57
<< alu1 >>
rect -2 95 52 100
rect -2 93 43 95
rect 45 93 52 95
rect -2 92 52 93
rect -2 90 7 92
rect 9 90 31 92
rect 33 90 52 92
rect -2 88 52 90
rect 6 82 10 88
rect 6 80 7 82
rect 9 80 10 82
rect 6 78 10 80
rect 18 81 22 83
rect 18 79 19 81
rect 21 79 22 81
rect 18 73 22 79
rect 30 82 34 88
rect 30 80 31 82
rect 33 80 34 82
rect 30 78 34 80
rect 8 71 22 73
rect 8 69 19 71
rect 21 69 22 71
rect 8 67 22 69
rect 8 39 12 67
rect 28 63 32 73
rect 18 57 32 63
rect 42 67 46 69
rect 42 65 43 67
rect 45 65 46 67
rect 42 59 46 65
rect 42 57 43 59
rect 45 57 46 59
rect 18 52 22 57
rect 16 50 22 52
rect 42 51 46 57
rect 16 48 17 50
rect 19 48 22 50
rect 16 46 22 48
rect 26 50 48 51
rect 26 48 28 50
rect 30 48 48 50
rect 26 47 48 48
rect 27 40 40 42
rect 8 37 14 39
rect 8 35 11 37
rect 13 35 14 37
rect 8 29 14 35
rect 27 38 37 40
rect 39 38 40 40
rect 27 36 40 38
rect 27 33 33 36
rect 8 27 11 29
rect 13 27 14 29
rect 8 25 14 27
rect 18 27 33 33
rect 44 32 48 47
rect 42 30 48 32
rect 42 28 43 30
rect 45 28 48 30
rect 18 17 22 27
rect 30 21 34 23
rect 30 19 31 21
rect 33 19 34 21
rect 30 12 34 19
rect 42 22 48 28
rect 42 20 43 22
rect 45 20 48 22
rect 42 18 48 20
rect -2 11 52 12
rect -2 9 31 11
rect 33 9 52 11
rect -2 7 52 9
rect -2 5 43 7
rect 45 5 52 7
rect -2 0 52 5
<< ptie >>
rect 41 7 47 9
rect 41 5 43 7
rect 45 5 47 7
rect 41 3 47 5
<< ntie >>
rect 41 95 47 97
rect 41 93 43 95
rect 45 93 47 95
rect 41 91 47 93
<< nmos >>
rect 17 6 19 39
rect 25 6 27 39
rect 37 18 39 33
<< pmos >>
rect 13 55 15 94
rect 25 55 27 94
rect 37 55 39 85
<< polyct1 >>
rect 17 48 19 50
rect 28 48 30 50
rect 37 38 39 40
<< ndifct1 >>
rect 11 35 13 37
rect 11 27 13 29
rect 31 19 33 21
rect 43 28 45 30
rect 43 20 45 22
rect 31 9 33 11
<< ntiect1 >>
rect 43 93 45 95
<< ptiect1 >>
rect 43 5 45 7
<< pdifct1 >>
rect 7 90 9 92
rect 7 80 9 82
rect 19 79 21 81
rect 19 69 21 71
rect 31 90 33 92
rect 31 80 33 82
rect 43 65 45 67
rect 43 57 45 59
<< labels >>
rlabel alu1 20 25 20 25 6 a
rlabel alu1 10 50 10 50 6 z
rlabel alu1 20 55 20 55 6 b
rlabel alu1 20 75 20 75 6 z
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 35 30 35 6 a
rlabel alu1 30 65 30 65 6 b
rlabel alu1 25 94 25 94 6 vdd
<< end >>
