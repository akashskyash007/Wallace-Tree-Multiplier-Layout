magic
tech scmos
timestamp 1199541709
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -2 48 62 104
<< pwell >>
rect -2 -4 62 48
<< poly >>
rect 47 95 49 98
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 11 43 13 65
rect 23 63 25 65
rect 17 61 25 63
rect 17 59 19 61
rect 21 59 23 61
rect 17 57 23 59
rect 35 53 37 65
rect 35 51 43 53
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 27 45 33 47
rect 27 43 29 45
rect 31 43 33 45
rect 47 43 49 55
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 11 25 13 37
rect 17 41 23 43
rect 27 41 49 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 17 35 25 37
rect 23 25 25 35
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 35 27 43 29
rect 35 25 37 27
rect 47 25 49 41
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 47 2 49 5
<< ndif >>
rect 15 31 21 33
rect 15 29 17 31
rect 19 29 21 31
rect 15 25 21 29
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 15 35 19
rect 37 15 47 25
rect 39 11 47 15
rect 39 9 41 11
rect 43 9 47 11
rect 39 5 47 9
rect 49 21 57 25
rect 49 19 53 21
rect 55 19 57 21
rect 49 5 57 19
<< pdif >>
rect 3 91 9 93
rect 39 91 47 95
rect 3 89 5 91
rect 7 89 9 91
rect 3 85 9 89
rect 39 89 41 91
rect 43 89 47 91
rect 39 85 47 89
rect 3 65 11 85
rect 13 65 23 85
rect 25 81 35 85
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 65 35 69
rect 37 65 47 85
rect 39 55 47 65
rect 49 81 57 95
rect 49 79 53 81
rect 55 79 57 81
rect 49 71 57 79
rect 49 69 53 71
rect 55 69 57 71
rect 49 61 57 69
rect 49 59 53 61
rect 55 59 57 61
rect 49 55 57 59
<< alu1 >>
rect -2 95 62 100
rect -2 93 17 95
rect 19 93 29 95
rect 31 93 62 95
rect -2 91 62 93
rect -2 89 5 91
rect 7 89 41 91
rect 43 89 62 91
rect -2 88 62 89
rect 8 41 12 82
rect 8 39 9 41
rect 11 39 12 41
rect 8 38 12 39
rect 18 61 22 82
rect 28 81 32 82
rect 28 79 29 81
rect 31 79 32 81
rect 28 78 32 79
rect 29 72 31 78
rect 28 71 32 72
rect 28 69 29 71
rect 31 69 32 71
rect 28 68 32 69
rect 18 59 19 61
rect 21 59 22 61
rect 18 41 22 59
rect 29 46 31 68
rect 38 51 42 82
rect 38 49 39 51
rect 41 49 42 51
rect 28 45 32 46
rect 28 43 29 45
rect 31 43 32 45
rect 28 42 32 43
rect 18 39 19 41
rect 21 39 22 41
rect 18 38 22 39
rect 16 31 20 32
rect 29 31 31 42
rect 16 29 17 31
rect 19 29 31 31
rect 38 31 42 49
rect 38 29 39 31
rect 41 29 42 31
rect 16 28 20 29
rect 4 21 8 22
rect 28 21 32 22
rect 4 19 5 21
rect 7 19 29 21
rect 31 19 32 21
rect 4 18 8 19
rect 28 18 32 19
rect 38 18 42 29
rect 48 81 56 82
rect 48 79 53 81
rect 55 79 56 81
rect 48 78 56 79
rect 48 72 52 78
rect 48 71 56 72
rect 48 69 53 71
rect 55 69 56 71
rect 48 68 56 69
rect 48 62 52 68
rect 48 61 56 62
rect 48 59 53 61
rect 55 59 56 61
rect 48 58 56 59
rect 48 22 52 58
rect 48 21 56 22
rect 48 19 53 21
rect 55 19 56 21
rect 48 18 56 19
rect -2 11 62 12
rect -2 9 41 11
rect 43 9 62 11
rect -2 7 62 9
rect -2 5 5 7
rect 7 5 17 7
rect 19 5 29 7
rect 31 5 62 7
rect -2 0 62 5
<< ptie >>
rect 3 7 33 9
rect 3 5 5 7
rect 7 5 17 7
rect 19 5 29 7
rect 31 5 33 7
rect 3 3 33 5
<< ntie >>
rect 15 95 33 97
rect 15 93 17 95
rect 19 93 29 95
rect 31 93 33 95
rect 15 91 33 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 47 5 49 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 55 49 95
<< polyct1 >>
rect 19 59 21 61
rect 39 49 41 51
rect 29 43 31 45
rect 9 39 11 41
rect 19 39 21 41
rect 39 29 41 31
<< ndifct1 >>
rect 17 29 19 31
rect 5 19 7 21
rect 29 19 31 21
rect 41 9 43 11
rect 53 19 55 21
<< ntiect1 >>
rect 17 93 19 95
rect 29 93 31 95
<< ptiect1 >>
rect 5 5 7 7
rect 17 5 19 7
rect 29 5 31 7
<< pdifct1 >>
rect 5 89 7 91
rect 41 89 43 91
rect 29 79 31 81
rect 29 69 31 71
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
<< labels >>
rlabel alu1 10 60 10 60 6 i0
rlabel polyct1 20 60 20 60 6 i1
rlabel ptiect1 30 6 30 6 6 vss
rlabel polyct1 40 50 40 50 6 i2
rlabel ntiect1 30 94 30 94 6 vdd
rlabel alu1 50 50 50 50 6 q
<< end >>
