magic
tech scmos
timestamp 1199201899
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 31 66 33 71
rect 41 66 43 71
rect 9 61 11 65
rect 19 61 21 65
rect 31 47 33 50
rect 30 45 37 47
rect 9 39 11 45
rect 19 42 21 45
rect 30 43 33 45
rect 35 43 37 45
rect 19 40 26 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 19 38 22 40
rect 24 38 26 40
rect 19 36 26 38
rect 30 41 37 43
rect 9 33 15 35
rect 13 24 15 33
rect 23 28 25 36
rect 30 28 32 41
rect 41 37 43 50
rect 41 35 47 37
rect 41 33 43 35
rect 45 33 47 35
rect 37 31 47 33
rect 37 28 39 31
rect 13 13 15 18
rect 23 13 25 18
rect 30 13 32 18
rect 37 13 39 18
<< ndif >>
rect 18 24 23 28
rect 3 18 13 24
rect 15 22 23 24
rect 15 20 18 22
rect 20 20 23 22
rect 15 18 23 20
rect 25 18 30 28
rect 32 18 37 28
rect 39 22 50 28
rect 39 20 45 22
rect 47 20 50 22
rect 39 18 50 20
rect 3 11 10 18
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
<< pdif >>
rect 23 71 29 73
rect 23 69 25 71
rect 27 69 29 71
rect 23 66 29 69
rect 23 61 31 66
rect 4 58 9 61
rect 2 56 9 58
rect 2 54 4 56
rect 6 54 9 56
rect 2 49 9 54
rect 2 47 4 49
rect 6 47 9 49
rect 2 45 9 47
rect 11 59 19 61
rect 11 57 14 59
rect 16 57 19 59
rect 11 45 19 57
rect 21 50 31 61
rect 33 61 41 66
rect 33 59 36 61
rect 38 59 41 61
rect 33 54 41 59
rect 33 52 36 54
rect 38 52 41 54
rect 33 50 41 52
rect 43 64 50 66
rect 43 62 46 64
rect 48 62 50 64
rect 43 50 50 62
rect 21 45 26 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 71 58 79
rect -2 69 25 71
rect 27 69 58 71
rect -2 68 58 69
rect 2 56 7 63
rect 2 54 4 56
rect 6 54 7 56
rect 2 50 7 54
rect 2 49 6 50
rect 2 47 4 49
rect 2 22 6 47
rect 21 50 31 54
rect 21 47 25 50
rect 18 41 25 47
rect 42 46 47 55
rect 31 45 47 46
rect 31 43 33 45
rect 35 43 47 45
rect 31 42 47 43
rect 21 40 25 41
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 21 38 22 40
rect 24 38 25 40
rect 21 34 31 38
rect 41 35 47 38
rect 41 33 43 35
rect 45 33 47 35
rect 41 30 47 33
rect 10 26 31 30
rect 35 26 47 30
rect 35 22 39 26
rect 2 17 15 22
rect 25 18 39 22
rect -2 11 58 12
rect -2 9 6 11
rect 8 9 58 11
rect -2 1 58 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 13 18 15 24
rect 23 18 25 28
rect 30 18 32 28
rect 37 18 39 28
<< pmos >>
rect 9 45 11 61
rect 19 45 21 61
rect 31 50 33 66
rect 41 50 43 66
<< polyct1 >>
rect 33 43 35 45
rect 11 35 13 37
rect 22 38 24 40
rect 43 33 45 35
<< ndifct0 >>
rect 18 20 20 22
rect 45 20 47 22
<< ndifct1 >>
rect 6 9 8 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 14 57 16 59
rect 36 59 38 61
rect 36 52 38 54
rect 46 62 48 64
<< pdifct1 >>
rect 25 69 27 71
rect 4 54 6 56
rect 4 47 6 49
<< alu0 >>
rect 45 64 49 68
rect 13 61 39 63
rect 13 59 36 61
rect 38 59 39 61
rect 45 62 46 64
rect 48 62 49 64
rect 45 60 49 62
rect 13 57 14 59
rect 16 57 17 59
rect 13 55 17 57
rect 35 54 39 59
rect 6 45 7 50
rect 35 52 36 54
rect 38 52 39 54
rect 35 50 39 52
rect 6 22 22 23
rect 15 20 18 22
rect 20 20 22 22
rect 15 19 22 20
rect 43 22 49 23
rect 43 20 45 22
rect 47 20 49 22
rect 43 12 49 20
<< labels >>
rlabel alu0 37 56 37 56 6 n3
rlabel alu0 26 61 26 61 6 n3
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 44 20 44 6 a3
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 36 20 36 20 6 a1
rlabel alu1 28 20 28 20 6 a1
rlabel alu1 28 28 28 28 6 b
rlabel alu1 28 36 28 36 6 a3
rlabel alu1 36 44 36 44 6 a2
rlabel alu1 28 52 28 52 6 a3
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 32 44 32 6 a1
rlabel alu1 44 48 44 48 6 a2
<< end >>
