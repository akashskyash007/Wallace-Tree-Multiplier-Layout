magic
tech scmos
timestamp 1199202023
<< ab >>
rect 0 0 32 80
<< nwell >>
rect -5 36 37 88
<< pwell >>
rect -5 -8 37 36
<< poly >>
rect 9 70 11 74
rect 21 60 23 65
rect 9 39 11 42
rect 21 39 23 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 21 37 27 39
rect 21 35 23 37
rect 25 35 27 37
rect 21 33 27 35
rect 9 30 11 33
rect 21 30 23 33
rect 21 16 23 21
rect 9 11 11 16
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 16 9 19
rect 11 21 21 30
rect 23 28 30 30
rect 23 26 26 28
rect 28 26 30 28
rect 23 24 30 26
rect 23 21 28 24
rect 11 20 19 21
rect 11 18 15 20
rect 17 18 19 20
rect 11 16 19 18
<< pdif >>
rect 4 63 9 70
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 68 19 70
rect 11 66 15 68
rect 17 66 19 68
rect 11 60 19 66
rect 11 42 21 60
rect 23 55 28 60
rect 23 53 30 55
rect 23 51 26 53
rect 28 51 30 53
rect 23 49 30 51
rect 23 42 28 49
<< alu1 >>
rect -2 81 34 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 34 81
rect -2 68 34 79
rect 2 62 7 63
rect 2 61 15 62
rect 2 59 4 61
rect 6 59 15 61
rect 2 58 15 59
rect 2 54 6 58
rect 2 52 4 54
rect 2 30 6 52
rect 26 39 30 47
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 18 37 30 39
rect 18 35 23 37
rect 25 35 30 37
rect 18 33 30 35
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect -2 1 34 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 34 1
rect -2 -2 34 -1
<< ptie >>
rect 0 1 32 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 32 1
rect 0 -3 32 -1
<< ntie >>
rect 0 81 32 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 32 81
rect 0 77 32 79
<< nmos >>
rect 9 16 11 30
rect 21 21 23 30
<< pmos >>
rect 9 42 11 70
rect 21 42 23 60
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 23 35 25 37
<< ndifct0 >>
rect 26 26 28 28
rect 15 18 17 20
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
<< pdifct0 >>
rect 15 66 17 68
rect 26 51 28 53
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
<< alu0 >>
rect 13 66 15 68
rect 17 66 19 68
rect 13 65 19 66
rect 6 50 7 58
rect 10 53 30 54
rect 10 51 26 53
rect 28 51 30 53
rect 10 50 30 51
rect 10 37 14 50
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 10 28 30 29
rect 10 26 26 28
rect 28 26 30 28
rect 10 25 30 26
rect 13 20 19 21
rect 13 18 15 20
rect 17 18 19 20
rect 13 12 19 18
<< labels >>
rlabel alu0 12 39 12 39 6 an
rlabel alu0 20 27 20 27 6 an
rlabel alu0 20 52 20 52 6 an
rlabel alu1 4 40 4 40 6 z
rlabel alu1 16 6 16 6 6 vss
rlabel alu1 12 60 12 60 6 z
rlabel alu1 16 74 16 74 6 vdd
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 40 28 40 6 a
<< end >>
