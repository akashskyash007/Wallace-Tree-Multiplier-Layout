magic
tech scmos
timestamp 1199541918
<< ab >>
rect 0 0 210 100
<< nwell >>
rect -2 48 212 104
<< pwell >>
rect -2 -4 212 48
<< poly >>
rect 81 95 83 98
rect 93 95 95 98
rect 105 95 107 98
rect 117 95 119 98
rect 11 83 13 86
rect 23 83 25 86
rect 35 83 37 86
rect 47 83 49 86
rect 57 83 59 86
rect 11 43 13 65
rect 23 43 25 65
rect 35 53 37 65
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 25 43
rect 17 39 19 41
rect 21 39 25 41
rect 17 37 25 39
rect 33 51 43 53
rect 33 49 39 51
rect 41 49 43 51
rect 33 47 43 49
rect 11 27 13 37
rect 21 29 23 37
rect 33 25 35 47
rect 47 43 49 57
rect 57 53 59 57
rect 131 83 133 86
rect 143 83 145 86
rect 153 83 155 86
rect 165 83 167 86
rect 57 51 63 53
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 45 37 53 39
rect 45 25 47 37
rect 57 25 59 47
rect 81 43 83 55
rect 93 43 95 55
rect 75 41 95 43
rect 75 39 77 41
rect 79 39 95 41
rect 75 37 95 39
rect 81 25 83 37
rect 93 25 95 37
rect 105 43 107 55
rect 117 43 119 55
rect 131 43 133 69
rect 143 67 145 69
rect 153 67 155 69
rect 141 65 145 67
rect 151 65 155 67
rect 177 79 179 82
rect 187 79 189 82
rect 197 79 199 82
rect 141 43 143 65
rect 151 43 153 65
rect 165 63 167 65
rect 163 61 167 63
rect 163 43 165 61
rect 177 53 179 65
rect 187 53 189 65
rect 177 51 183 53
rect 177 49 179 51
rect 181 49 183 51
rect 105 41 123 43
rect 105 39 119 41
rect 121 39 123 41
rect 105 37 123 39
rect 127 41 133 43
rect 127 39 129 41
rect 131 39 133 41
rect 127 37 133 39
rect 137 41 143 43
rect 137 39 139 41
rect 141 39 143 41
rect 137 37 143 39
rect 147 41 153 43
rect 147 39 149 41
rect 151 39 153 41
rect 147 37 153 39
rect 157 41 165 43
rect 157 39 159 41
rect 161 39 165 41
rect 157 37 165 39
rect 105 25 107 37
rect 117 25 119 37
rect 131 25 133 37
rect 141 25 143 37
rect 151 25 153 37
rect 163 27 165 37
rect 175 47 183 49
rect 187 51 193 53
rect 187 49 189 51
rect 191 49 193 51
rect 187 47 193 49
rect 11 14 13 17
rect 21 14 23 17
rect 33 14 35 17
rect 45 14 47 17
rect 57 14 59 17
rect 175 25 177 47
rect 187 29 189 47
rect 185 27 189 29
rect 197 43 199 65
rect 197 41 203 43
rect 197 39 199 41
rect 201 39 203 41
rect 197 37 203 39
rect 185 25 187 27
rect 197 25 199 37
rect 131 14 133 17
rect 141 14 143 17
rect 151 14 153 17
rect 163 14 165 17
rect 175 14 177 17
rect 185 14 187 17
rect 197 14 199 17
rect 81 2 83 5
rect 93 2 95 5
rect 105 2 107 5
rect 117 2 119 5
<< ndif >>
rect 17 27 21 29
rect 3 17 11 27
rect 13 17 21 27
rect 23 25 31 29
rect 159 25 163 27
rect 23 21 33 25
rect 23 19 27 21
rect 29 19 33 21
rect 23 17 33 19
rect 35 21 45 25
rect 35 19 39 21
rect 41 19 45 21
rect 35 17 45 19
rect 47 17 57 25
rect 59 21 67 25
rect 59 19 63 21
rect 65 19 67 21
rect 59 17 67 19
rect 73 21 81 25
rect 73 19 75 21
rect 77 19 81 21
rect 3 11 9 17
rect 49 11 55 17
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
rect 73 11 81 19
rect 73 9 75 11
rect 77 9 81 11
rect 73 5 81 9
rect 83 21 93 25
rect 83 19 87 21
rect 89 19 93 21
rect 83 5 93 19
rect 95 11 105 25
rect 95 9 99 11
rect 101 9 105 11
rect 95 5 105 9
rect 107 21 117 25
rect 107 19 111 21
rect 113 19 117 21
rect 107 5 117 19
rect 119 17 131 25
rect 133 17 141 25
rect 143 17 151 25
rect 153 21 163 25
rect 153 19 157 21
rect 159 19 163 21
rect 153 17 163 19
rect 165 25 169 27
rect 165 21 175 25
rect 165 19 169 21
rect 171 19 175 21
rect 165 17 175 19
rect 177 17 185 25
rect 187 21 197 25
rect 187 19 191 21
rect 193 19 197 21
rect 187 17 197 19
rect 199 21 207 25
rect 199 19 203 21
rect 205 19 207 21
rect 199 17 207 19
rect 119 11 129 17
rect 179 11 183 17
rect 119 9 123 11
rect 125 9 129 11
rect 119 5 129 9
rect 178 9 184 11
rect 178 7 180 9
rect 182 7 184 9
rect 178 5 184 7
<< pdif >>
rect 15 91 21 93
rect 73 91 81 95
rect 15 89 17 91
rect 19 89 21 91
rect 15 83 21 89
rect 73 89 75 91
rect 77 89 81 91
rect 3 81 11 83
rect 3 79 5 81
rect 7 79 11 81
rect 3 65 11 79
rect 13 65 23 83
rect 25 81 35 83
rect 25 79 29 81
rect 31 79 35 81
rect 25 65 35 79
rect 37 71 47 83
rect 37 69 41 71
rect 43 69 47 71
rect 37 65 47 69
rect 40 57 47 65
rect 49 57 57 83
rect 59 81 67 83
rect 59 79 63 81
rect 65 79 67 81
rect 59 57 67 79
rect 73 55 81 89
rect 83 71 93 95
rect 83 69 87 71
rect 89 69 93 71
rect 83 61 93 69
rect 83 59 87 61
rect 89 59 93 61
rect 83 55 93 59
rect 95 91 105 95
rect 95 89 99 91
rect 101 89 105 91
rect 95 55 105 89
rect 107 71 117 95
rect 107 69 111 71
rect 113 69 117 71
rect 107 61 117 69
rect 107 59 111 61
rect 113 59 117 61
rect 107 55 117 59
rect 119 91 129 95
rect 119 89 123 91
rect 125 89 129 91
rect 146 93 152 95
rect 146 91 148 93
rect 150 91 152 93
rect 146 89 152 91
rect 119 83 129 89
rect 147 83 151 89
rect 119 69 131 83
rect 133 81 143 83
rect 133 79 137 81
rect 139 79 143 81
rect 133 69 143 79
rect 145 69 153 83
rect 155 81 165 83
rect 155 79 159 81
rect 161 79 165 81
rect 155 69 165 79
rect 119 55 127 69
rect 157 65 165 69
rect 167 79 174 83
rect 201 81 207 83
rect 201 79 203 81
rect 205 79 207 81
rect 167 71 177 79
rect 167 69 171 71
rect 173 69 177 71
rect 167 65 177 69
rect 179 65 187 79
rect 189 65 197 79
rect 199 65 207 79
<< alu1 >>
rect -2 95 212 100
rect -2 93 31 95
rect 33 93 39 95
rect 41 93 47 95
rect 49 93 55 95
rect 57 93 63 95
rect 65 93 161 95
rect 163 93 169 95
rect 171 93 177 95
rect 179 93 185 95
rect 187 93 193 95
rect 195 93 212 95
rect -2 91 148 93
rect 150 91 212 93
rect -2 89 17 91
rect 19 89 75 91
rect 77 89 99 91
rect 101 89 123 91
rect 125 89 212 91
rect -2 88 212 89
rect 4 81 8 82
rect 28 81 32 82
rect 62 81 66 82
rect 136 81 140 82
rect 158 81 162 82
rect 202 81 206 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 63 81
rect 65 79 66 81
rect 4 78 8 79
rect 28 78 32 79
rect 62 78 66 79
rect 75 79 123 81
rect 8 41 12 72
rect 8 39 9 41
rect 11 39 12 41
rect 8 18 12 39
rect 18 41 22 72
rect 40 71 44 72
rect 75 71 77 79
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 29 69 41 71
rect 43 69 77 71
rect 29 22 31 69
rect 40 68 44 69
rect 38 51 42 62
rect 38 49 39 51
rect 41 49 42 51
rect 38 28 42 49
rect 48 41 52 62
rect 48 39 49 41
rect 51 39 52 41
rect 48 28 52 39
rect 58 51 62 62
rect 58 49 59 51
rect 61 49 62 51
rect 58 28 62 49
rect 75 42 77 69
rect 86 71 92 72
rect 86 69 87 71
rect 89 69 92 71
rect 86 68 92 69
rect 88 62 92 68
rect 86 61 92 62
rect 86 59 87 61
rect 89 59 92 61
rect 86 58 92 59
rect 75 41 80 42
rect 75 39 77 41
rect 79 39 80 41
rect 76 38 80 39
rect 88 22 92 58
rect 26 21 31 22
rect 26 19 27 21
rect 29 19 31 21
rect 38 21 42 22
rect 62 21 66 22
rect 38 19 39 21
rect 41 19 63 21
rect 65 19 66 21
rect 26 18 30 19
rect 38 18 42 19
rect 62 18 66 19
rect 74 21 78 22
rect 74 19 75 21
rect 77 19 78 21
rect 74 12 78 19
rect 86 21 92 22
rect 86 19 87 21
rect 89 19 92 21
rect 86 18 92 19
rect 108 71 114 72
rect 108 69 111 71
rect 113 69 114 71
rect 121 71 123 79
rect 136 79 137 81
rect 139 79 159 81
rect 161 79 203 81
rect 205 79 206 81
rect 136 78 140 79
rect 158 78 162 79
rect 202 78 206 79
rect 169 71 174 72
rect 121 69 161 71
rect 108 68 114 69
rect 108 62 112 68
rect 108 61 114 62
rect 108 59 111 61
rect 113 59 114 61
rect 108 58 114 59
rect 108 22 112 58
rect 118 41 122 42
rect 118 39 119 41
rect 121 39 122 41
rect 118 38 122 39
rect 128 41 132 62
rect 128 39 129 41
rect 131 39 132 41
rect 128 38 132 39
rect 138 41 142 62
rect 138 39 139 41
rect 141 39 142 41
rect 119 31 121 38
rect 119 29 131 31
rect 108 21 114 22
rect 108 19 111 21
rect 113 19 114 21
rect 129 21 131 29
rect 138 28 142 39
rect 148 41 152 62
rect 159 42 161 69
rect 169 69 171 71
rect 173 69 174 71
rect 169 68 174 69
rect 148 39 149 41
rect 151 39 152 41
rect 148 28 152 39
rect 158 41 162 42
rect 158 39 159 41
rect 161 39 162 41
rect 158 38 162 39
rect 169 31 171 68
rect 159 29 171 31
rect 178 51 182 62
rect 178 49 179 51
rect 181 49 182 51
rect 159 22 161 29
rect 178 28 182 49
rect 188 51 192 72
rect 188 49 189 51
rect 191 49 192 51
rect 188 28 192 49
rect 198 41 202 72
rect 198 39 199 41
rect 201 39 202 41
rect 198 28 202 39
rect 156 21 161 22
rect 129 19 157 21
rect 159 19 161 21
rect 108 18 114 19
rect 156 18 161 19
rect 168 21 172 22
rect 190 21 194 22
rect 168 19 169 21
rect 171 19 191 21
rect 193 19 194 21
rect 168 18 172 19
rect 190 18 194 19
rect 202 21 206 22
rect 202 19 203 21
rect 205 19 206 21
rect 202 12 206 19
rect -2 11 212 12
rect -2 9 5 11
rect 7 9 51 11
rect 53 9 75 11
rect 77 9 99 11
rect 101 9 123 11
rect 125 9 212 11
rect -2 7 19 9
rect 21 7 29 9
rect 31 7 39 9
rect 41 7 137 9
rect 139 7 147 9
rect 149 7 157 9
rect 159 7 168 9
rect 170 7 180 9
rect 182 7 193 9
rect 195 7 201 9
rect 203 7 212 9
rect -2 0 212 7
<< ptie >>
rect 17 9 43 11
rect 17 7 19 9
rect 21 7 29 9
rect 31 7 39 9
rect 41 7 43 9
rect 17 5 43 7
rect 135 9 172 11
rect 135 7 137 9
rect 139 7 147 9
rect 149 7 157 9
rect 159 7 168 9
rect 170 7 172 9
rect 135 5 172 7
rect 191 9 205 11
rect 191 7 193 9
rect 195 7 201 9
rect 203 7 205 9
rect 191 5 205 7
<< ntie >>
rect 29 95 67 97
rect 159 95 197 97
rect 29 93 31 95
rect 33 93 39 95
rect 41 93 47 95
rect 49 93 55 95
rect 57 93 63 95
rect 65 93 67 95
rect 29 91 67 93
rect 159 93 161 95
rect 163 93 169 95
rect 171 93 177 95
rect 179 93 185 95
rect 187 93 193 95
rect 195 93 197 95
rect 159 91 197 93
<< nmos >>
rect 11 17 13 27
rect 21 17 23 29
rect 33 17 35 25
rect 45 17 47 25
rect 57 17 59 25
rect 81 5 83 25
rect 93 5 95 25
rect 105 5 107 25
rect 117 5 119 25
rect 131 17 133 25
rect 141 17 143 25
rect 151 17 153 25
rect 163 17 165 27
rect 175 17 177 25
rect 185 17 187 25
rect 197 17 199 25
<< pmos >>
rect 11 65 13 83
rect 23 65 25 83
rect 35 65 37 83
rect 47 57 49 83
rect 57 57 59 83
rect 81 55 83 95
rect 93 55 95 95
rect 105 55 107 95
rect 117 55 119 95
rect 131 69 133 83
rect 143 69 145 83
rect 153 69 155 83
rect 165 65 167 83
rect 177 65 179 79
rect 187 65 189 79
rect 197 65 199 79
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 39 49 41 51
rect 59 49 61 51
rect 49 39 51 41
rect 77 39 79 41
rect 179 49 181 51
rect 119 39 121 41
rect 129 39 131 41
rect 139 39 141 41
rect 149 39 151 41
rect 159 39 161 41
rect 189 49 191 51
rect 199 39 201 41
<< ndifct1 >>
rect 27 19 29 21
rect 39 19 41 21
rect 63 19 65 21
rect 75 19 77 21
rect 5 9 7 11
rect 51 9 53 11
rect 75 9 77 11
rect 87 19 89 21
rect 99 9 101 11
rect 111 19 113 21
rect 157 19 159 21
rect 169 19 171 21
rect 191 19 193 21
rect 203 19 205 21
rect 123 9 125 11
rect 180 7 182 9
<< ntiect1 >>
rect 31 93 33 95
rect 39 93 41 95
rect 47 93 49 95
rect 55 93 57 95
rect 63 93 65 95
rect 161 93 163 95
rect 169 93 171 95
rect 177 93 179 95
rect 185 93 187 95
rect 193 93 195 95
<< ptiect1 >>
rect 19 7 21 9
rect 29 7 31 9
rect 39 7 41 9
rect 137 7 139 9
rect 147 7 149 9
rect 157 7 159 9
rect 168 7 170 9
rect 193 7 195 9
rect 201 7 203 9
<< pdifct1 >>
rect 17 89 19 91
rect 75 89 77 91
rect 5 79 7 81
rect 29 79 31 81
rect 41 69 43 71
rect 63 79 65 81
rect 87 69 89 71
rect 87 59 89 61
rect 99 89 101 91
rect 111 69 113 71
rect 111 59 113 61
rect 123 89 125 91
rect 148 91 150 93
rect 137 79 139 81
rect 159 79 161 81
rect 203 79 205 81
rect 171 69 173 71
<< labels >>
rlabel alu1 10 45 10 45 6 a1
rlabel alu1 20 50 20 50 6 b1
rlabel alu1 60 45 60 45 6 b2
rlabel alu1 50 45 50 45 6 a2
rlabel alu1 40 45 40 45 6 cin1
rlabel alu1 105 6 105 6 6 vss
rlabel alu1 110 45 110 45 6 sout
rlabel alu1 90 45 90 45 6 cout
rlabel alu1 105 94 105 94 6 vdd
rlabel alu1 150 45 150 45 6 cin2
rlabel alu1 140 45 140 45 6 b3
rlabel alu1 130 50 130 50 6 a3
rlabel alu1 180 45 180 45 6 cin3
rlabel alu1 200 50 200 50 6 b4
rlabel polyct1 190 50 190 50 6 a4
<< end >>
