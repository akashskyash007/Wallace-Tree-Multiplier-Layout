magic
tech scmos
timestamp 1199202778
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 11 70 13 74
rect 21 70 23 74
rect 37 70 39 74
rect 49 70 51 74
rect 11 53 13 56
rect 21 53 23 56
rect 11 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 12 30 14 33
rect 19 30 21 47
rect 37 39 39 42
rect 33 37 39 39
rect 33 35 35 37
rect 37 35 39 37
rect 49 39 51 42
rect 49 37 55 39
rect 49 35 51 37
rect 53 35 55 37
rect 26 33 39 35
rect 26 30 28 33
rect 36 30 38 33
rect 43 30 45 35
rect 49 33 55 35
rect 50 30 52 33
rect 12 11 14 16
rect 19 8 21 16
rect 26 12 28 16
rect 36 12 38 16
rect 43 8 45 16
rect 50 11 52 16
rect 19 6 45 8
<< ndif >>
rect 2 20 12 30
rect 2 18 4 20
rect 6 18 12 20
rect 2 16 12 18
rect 14 16 19 30
rect 21 16 26 30
rect 28 21 36 30
rect 28 19 31 21
rect 33 19 36 21
rect 28 16 36 19
rect 38 16 43 30
rect 45 16 50 30
rect 52 20 60 30
rect 52 18 55 20
rect 57 18 60 20
rect 52 16 60 18
<< pdif >>
rect 3 68 11 70
rect 3 66 6 68
rect 8 66 11 68
rect 3 56 11 66
rect 13 61 21 70
rect 13 59 16 61
rect 18 59 21 61
rect 13 56 21 59
rect 23 68 37 70
rect 23 66 29 68
rect 31 66 37 68
rect 23 56 37 66
rect 25 42 37 56
rect 39 61 49 70
rect 39 59 43 61
rect 45 59 49 61
rect 39 53 49 59
rect 39 51 43 53
rect 45 51 49 53
rect 39 42 49 51
rect 51 68 59 70
rect 51 66 54 68
rect 56 66 59 68
rect 51 61 59 66
rect 51 59 54 61
rect 56 59 59 61
rect 51 42 59 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 61 47 62
rect 2 59 16 61
rect 18 59 43 61
rect 45 59 47 61
rect 2 58 47 59
rect 2 29 6 58
rect 17 51 23 54
rect 17 49 19 51
rect 21 49 23 51
rect 41 53 47 58
rect 41 51 43 53
rect 45 51 47 53
rect 41 50 47 51
rect 17 46 23 49
rect 17 42 31 46
rect 38 42 47 46
rect 38 38 42 42
rect 12 37 26 38
rect 13 35 26 37
rect 12 34 26 35
rect 33 37 42 38
rect 33 35 35 37
rect 37 35 42 37
rect 33 34 42 35
rect 49 37 55 38
rect 49 35 51 37
rect 53 35 55 37
rect 22 30 26 34
rect 49 30 55 35
rect 2 25 15 29
rect 22 26 55 30
rect 11 22 15 25
rect 11 21 35 22
rect 11 19 31 21
rect 33 19 35 21
rect 11 18 35 19
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 12 16 14 30
rect 19 16 21 30
rect 26 16 28 30
rect 36 16 38 30
rect 43 16 45 30
rect 50 16 52 30
<< pmos >>
rect 11 56 13 70
rect 21 56 23 70
rect 37 42 39 70
rect 49 42 51 70
<< polyct0 >>
rect 11 35 12 37
<< polyct1 >>
rect 19 49 21 51
rect 12 35 13 37
rect 35 35 37 37
rect 51 35 53 37
<< ndifct0 >>
rect 4 18 6 20
rect 55 18 57 20
<< ndifct1 >>
rect 31 19 33 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 6 66 8 68
rect 29 66 31 68
rect 54 66 56 68
rect 54 59 56 61
<< pdifct1 >>
rect 16 59 18 61
rect 43 59 45 61
rect 43 51 45 53
<< alu0 >>
rect 4 66 6 68
rect 8 66 10 68
rect 4 65 10 66
rect 27 66 29 68
rect 31 66 33 68
rect 27 65 33 66
rect 52 66 54 68
rect 56 66 58 68
rect 52 61 58 66
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
rect 10 38 16 39
rect 10 37 12 38
rect 10 35 11 37
rect 10 34 12 35
rect 10 33 22 34
rect 3 20 7 22
rect 3 18 4 20
rect 6 18 7 20
rect 54 20 58 22
rect 54 18 55 20
rect 57 18 58 20
rect 3 12 7 18
rect 54 12 58 18
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 60 12 60 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 48 20 48 6 b
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 44 44 44 6 c
rlabel alu1 44 56 44 56 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 32 52 32 6 a
<< end >>
