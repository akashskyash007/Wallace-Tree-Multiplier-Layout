magic
tech scmos
timestamp 1199542787
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 19 94 21 98
rect 27 94 29 98
rect 35 94 37 98
rect 43 94 45 98
rect 19 53 21 56
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 11 47 23 49
rect 11 25 13 47
rect 27 43 29 56
rect 35 53 37 56
rect 43 53 45 56
rect 35 51 39 53
rect 43 51 49 53
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 23 37 33 39
rect 23 25 25 37
rect 37 33 39 51
rect 47 43 49 51
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 35 27 43 29
rect 35 24 37 27
rect 47 25 49 37
rect 11 11 13 15
rect 23 11 25 15
rect 35 10 37 14
rect 47 11 49 15
<< ndif >>
rect 3 15 11 25
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 15 23 19
rect 25 24 30 25
rect 42 24 47 25
rect 25 15 35 24
rect 3 11 9 15
rect 27 14 35 15
rect 37 21 47 24
rect 37 19 41 21
rect 43 19 47 21
rect 37 15 47 19
rect 49 15 57 25
rect 37 14 45 15
rect 27 11 33 14
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 27 9 29 11
rect 31 9 33 11
rect 51 11 57 15
rect 27 7 33 9
rect 51 9 53 11
rect 55 9 57 11
rect 51 6 57 9
<< pdif >>
rect 14 85 19 94
rect 7 81 19 85
rect 7 79 9 81
rect 11 79 19 81
rect 7 71 19 79
rect 7 69 9 71
rect 11 69 19 71
rect 7 61 19 69
rect 7 59 9 61
rect 11 59 19 61
rect 7 56 19 59
rect 21 56 27 94
rect 29 56 35 94
rect 37 56 43 94
rect 45 91 53 94
rect 45 89 49 91
rect 51 89 53 91
rect 45 56 53 89
rect 7 55 13 56
<< alu1 >>
rect -2 91 62 100
rect -2 89 49 91
rect 51 89 62 91
rect -2 88 62 89
rect 8 81 12 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 71 12 79
rect 8 69 9 71
rect 11 69 12 71
rect 8 61 12 69
rect 8 59 9 61
rect 11 59 12 61
rect 8 22 12 59
rect 18 51 22 83
rect 18 49 19 51
rect 21 49 22 51
rect 18 27 22 49
rect 28 41 32 83
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 31 42 83
rect 38 29 39 31
rect 41 29 42 31
rect 38 27 42 29
rect 48 41 52 83
rect 48 39 49 41
rect 51 39 52 41
rect 48 27 52 39
rect 8 21 45 22
rect 8 19 17 21
rect 19 19 41 21
rect 43 19 45 21
rect 8 18 45 19
rect 8 17 12 18
rect -2 11 62 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 53 11
rect 55 9 62 11
rect -2 0 62 9
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 14 37 24
rect 47 15 49 25
<< pmos >>
rect 19 56 21 94
rect 27 56 29 94
rect 35 56 37 94
rect 43 56 45 94
<< polyct1 >>
rect 19 49 21 51
rect 29 39 31 41
rect 49 39 51 41
rect 39 29 41 31
<< ndifct1 >>
rect 17 19 19 21
rect 41 19 43 21
rect 5 9 7 11
rect 29 9 31 11
rect 53 9 55 11
<< pdifct1 >>
rect 9 79 11 81
rect 9 69 11 71
rect 9 59 11 61
rect 49 89 51 91
<< labels >>
rlabel alu1 10 50 10 50 6 nq
rlabel alu1 20 20 20 20 6 nq
rlabel alu1 20 55 20 55 6 i1
rlabel alu1 30 20 30 20 6 nq
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 40 20 40 20 6 nq
rlabel alu1 30 55 30 55 6 i0
rlabel alu1 40 55 40 55 6 i2
rlabel alu1 30 94 30 94 6 vdd
rlabel alu1 50 55 50 55 6 i3
<< end >>
