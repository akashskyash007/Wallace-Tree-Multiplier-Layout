magic
tech scmos
timestamp 1199202250
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 10 65 12 69
rect 20 57 22 61
rect 10 36 12 41
rect 20 36 22 41
rect 10 34 30 36
rect 10 26 12 34
rect 20 32 26 34
rect 28 32 30 34
rect 20 30 30 32
rect 20 26 22 30
rect 10 11 12 16
rect 20 11 22 16
<< ndif >>
rect 2 17 10 26
rect 2 15 4 17
rect 6 16 10 17
rect 12 24 20 26
rect 12 22 15 24
rect 17 22 20 24
rect 12 16 20 22
rect 22 20 30 26
rect 22 18 26 20
rect 28 18 30 20
rect 22 16 30 18
rect 6 15 8 16
rect 2 13 8 15
<< pdif >>
rect 2 63 10 65
rect 2 61 5 63
rect 7 61 10 63
rect 2 56 10 61
rect 2 54 5 56
rect 7 54 10 56
rect 2 41 10 54
rect 12 57 17 65
rect 12 49 20 57
rect 12 47 15 49
rect 17 47 20 49
rect 12 41 20 47
rect 22 55 30 57
rect 22 53 25 55
rect 27 53 30 55
rect 22 48 30 53
rect 22 46 25 48
rect 27 46 30 48
rect 22 41 30 46
<< alu1 >>
rect -2 67 34 72
rect -2 65 24 67
rect 26 65 34 67
rect -2 64 34 65
rect 2 49 19 50
rect 2 47 15 49
rect 17 47 19 49
rect 2 46 19 47
rect 2 27 6 46
rect 17 38 30 42
rect 26 34 30 38
rect 28 32 30 34
rect 26 29 30 32
rect 2 24 22 27
rect 2 22 15 24
rect 17 22 22 24
rect 2 21 22 22
rect -2 7 34 8
rect -2 5 5 7
rect 7 5 25 7
rect 27 5 34 7
rect -2 0 34 5
<< ptie >>
rect 3 7 29 9
rect 3 5 5 7
rect 7 5 25 7
rect 27 5 29 7
rect 3 3 29 5
<< ntie >>
rect 22 67 28 69
rect 22 65 24 67
rect 26 65 28 67
rect 22 63 28 65
<< nmos >>
rect 10 16 12 26
rect 20 16 22 26
<< pmos >>
rect 10 41 12 65
rect 20 41 22 57
<< polyct1 >>
rect 26 32 28 34
<< ndifct0 >>
rect 4 15 6 17
rect 26 18 28 20
<< ndifct1 >>
rect 15 22 17 24
<< ntiect1 >>
rect 24 65 26 67
<< ptiect1 >>
rect 5 5 7 7
rect 25 5 27 7
<< pdifct0 >>
rect 5 61 7 63
rect 5 54 7 56
rect 25 53 27 55
rect 25 46 27 48
<< pdifct1 >>
rect 15 47 17 49
<< alu0 >>
rect 3 63 9 64
rect 3 61 5 63
rect 7 61 9 63
rect 3 56 9 61
rect 3 54 5 56
rect 7 54 9 56
rect 3 53 9 54
rect 23 55 29 64
rect 23 53 25 55
rect 27 53 29 55
rect 23 48 29 53
rect 23 46 25 48
rect 27 46 29 48
rect 23 45 29 46
rect 24 31 26 38
rect 25 20 29 22
rect 25 18 26 20
rect 28 18 29 20
rect 2 17 8 18
rect 2 15 4 17
rect 6 15 8 17
rect 2 8 8 15
rect 25 8 29 18
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 24 20 24 6 z
rlabel alu1 20 40 20 40 6 a
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 32 28 32 6 a
<< end >>
