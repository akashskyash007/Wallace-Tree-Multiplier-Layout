magic
tech scmos
timestamp 1199201727
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 55 70 57 74
rect 65 70 67 74
rect 35 64 37 69
rect 45 64 47 69
rect 35 47 37 50
rect 45 47 47 50
rect 35 45 48 47
rect 38 43 44 45
rect 46 43 48 45
rect 9 39 11 42
rect 19 39 21 42
rect 38 41 48 43
rect 9 37 21 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 26 37 33 39
rect 26 35 28 37
rect 30 35 33 37
rect 26 33 33 35
rect 9 30 11 33
rect 19 30 21 33
rect 31 30 33 33
rect 38 30 40 41
rect 55 39 57 43
rect 65 40 67 43
rect 52 37 58 39
rect 65 38 78 40
rect 52 35 54 37
rect 56 35 58 37
rect 45 33 58 35
rect 69 37 78 38
rect 69 35 74 37
rect 76 35 78 37
rect 45 30 47 33
rect 55 30 57 33
rect 62 30 64 34
rect 69 33 78 35
rect 69 30 71 33
rect 9 11 11 16
rect 19 11 21 16
rect 31 11 33 16
rect 38 8 40 16
rect 45 12 47 16
rect 55 12 57 16
rect 62 8 64 16
rect 69 11 71 16
rect 38 6 64 8
<< ndif >>
rect 2 20 9 30
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 26 19 30
rect 11 24 14 26
rect 16 24 19 26
rect 11 16 19 24
rect 21 16 31 30
rect 33 16 38 30
rect 40 16 45 30
rect 47 20 55 30
rect 47 18 50 20
rect 52 18 55 20
rect 47 16 55 18
rect 57 16 62 30
rect 64 16 69 30
rect 71 20 78 30
rect 71 18 74 20
rect 76 18 78 20
rect 71 16 78 18
rect 23 11 29 16
rect 23 9 25 11
rect 27 9 29 11
rect 23 7 29 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 42 9 59
rect 11 53 19 70
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 68 33 70
rect 21 66 27 68
rect 29 66 33 68
rect 21 64 33 66
rect 49 64 55 70
rect 21 61 35 64
rect 21 59 27 61
rect 29 59 35 61
rect 21 50 35 59
rect 37 61 45 64
rect 37 59 40 61
rect 42 59 45 61
rect 37 54 45 59
rect 37 52 40 54
rect 42 52 45 54
rect 37 50 45 52
rect 47 62 55 64
rect 47 60 50 62
rect 52 60 55 62
rect 47 50 55 60
rect 21 42 33 50
rect 50 43 55 50
rect 57 61 65 70
rect 57 59 60 61
rect 62 59 65 61
rect 57 54 65 59
rect 57 52 60 54
rect 62 52 65 54
rect 57 43 65 52
rect 67 68 75 70
rect 67 66 70 68
rect 72 66 75 68
rect 67 61 75 66
rect 67 59 70 61
rect 72 59 75 61
rect 67 43 75 59
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 13 53 17 55
rect 13 51 14 53
rect 16 51 17 53
rect 13 47 17 51
rect 2 46 17 47
rect 2 44 14 46
rect 16 44 17 46
rect 2 42 17 44
rect 2 30 6 42
rect 2 26 17 30
rect 2 25 14 26
rect 13 24 14 25
rect 16 24 17 26
rect 13 22 17 24
rect 34 38 38 47
rect 66 46 70 55
rect 42 45 70 46
rect 42 43 44 45
rect 46 43 70 45
rect 42 42 70 43
rect 74 38 78 39
rect 34 37 58 38
rect 34 35 54 37
rect 56 35 58 37
rect 34 34 58 35
rect 72 37 78 38
rect 72 35 74 37
rect 76 35 78 37
rect 72 30 78 35
rect 29 26 78 30
rect 58 17 62 26
rect -2 11 82 12
rect -2 9 25 11
rect 27 9 82 11
rect -2 1 82 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 31 16 33 30
rect 38 16 40 30
rect 45 16 47 30
rect 55 16 57 30
rect 62 16 64 30
rect 69 16 71 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 35 50 37 64
rect 45 50 47 64
rect 55 43 57 70
rect 65 43 67 70
<< polyct0 >>
rect 17 35 19 37
rect 28 35 30 37
<< polyct1 >>
rect 44 43 46 45
rect 54 35 56 37
rect 74 35 76 37
<< ndifct0 >>
rect 4 18 6 20
rect 50 18 52 20
rect 74 18 76 20
<< ndifct1 >>
rect 14 24 16 26
rect 25 9 27 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 27 66 29 68
rect 27 59 29 61
rect 40 59 42 61
rect 40 52 42 54
rect 50 60 52 62
rect 60 59 62 61
rect 60 52 62 54
rect 70 66 72 68
rect 70 59 72 61
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 25 66 27 68
rect 29 66 31 68
rect 25 61 31 66
rect 25 59 27 61
rect 29 59 31 61
rect 25 58 31 59
rect 39 61 43 63
rect 39 59 40 61
rect 42 59 43 61
rect 39 54 43 59
rect 49 62 53 68
rect 68 66 70 68
rect 72 66 74 68
rect 49 60 50 62
rect 52 60 53 62
rect 49 58 53 60
rect 59 61 63 63
rect 59 59 60 61
rect 62 59 63 61
rect 59 54 63 59
rect 68 61 74 66
rect 68 59 70 61
rect 72 59 74 61
rect 68 58 74 59
rect 20 52 40 54
rect 42 52 60 54
rect 62 52 63 54
rect 20 50 63 52
rect 20 38 24 50
rect 15 37 24 38
rect 15 35 17 37
rect 19 35 24 37
rect 15 34 24 35
rect 20 21 24 34
rect 27 37 31 39
rect 27 35 28 37
rect 30 35 31 37
rect 27 30 31 35
rect 27 26 29 30
rect 2 20 8 21
rect 2 18 4 20
rect 6 18 8 20
rect 2 12 8 18
rect 20 20 54 21
rect 20 18 50 20
rect 52 18 54 20
rect 20 17 54 18
rect 73 20 77 22
rect 73 18 74 20
rect 76 18 77 20
rect 73 12 77 18
<< labels >>
rlabel alu0 19 36 19 36 6 zn
rlabel alu0 37 19 37 19 6 zn
rlabel alu0 41 56 41 56 6 zn
rlabel alu0 61 56 61 56 6 zn
rlabel alu1 12 28 12 28 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 c
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 36 44 36 6 c
rlabel alu1 52 36 52 36 6 c
rlabel alu1 52 28 52 28 6 a
rlabel alu1 52 44 52 44 6 b
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 24 60 24 6 a
rlabel alu1 76 36 76 36 6 a
rlabel alu1 68 28 68 28 6 a
rlabel alu1 60 44 60 44 6 b
rlabel alu1 68 52 68 52 6 b
<< end >>
