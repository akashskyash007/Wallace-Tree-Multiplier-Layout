magic
tech scmos
timestamp 1199201944
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 67 11 72
rect 19 67 21 72
rect 29 67 31 72
rect 39 67 41 72
rect 49 67 51 72
rect 59 67 61 72
rect 9 39 11 50
rect 19 47 21 50
rect 29 47 31 50
rect 19 45 31 47
rect 25 43 27 45
rect 29 43 31 45
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 25 37 31 43
rect 39 39 41 50
rect 49 39 51 42
rect 25 35 27 37
rect 29 35 31 37
rect 9 33 15 35
rect 19 33 31 35
rect 35 37 41 39
rect 35 35 37 37
rect 39 35 41 37
rect 35 33 41 35
rect 45 37 51 39
rect 45 35 47 37
rect 49 35 51 37
rect 59 35 61 42
rect 45 33 51 35
rect 55 33 70 35
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 30 38 33
rect 48 30 50 33
rect 55 30 57 33
rect 64 31 66 33
rect 68 31 70 33
rect 12 15 14 19
rect 19 15 21 19
rect 29 8 31 13
rect 36 8 38 13
rect 64 29 70 31
rect 48 6 50 10
rect 55 6 57 10
<< ndif >>
rect 3 19 12 30
rect 14 19 19 30
rect 21 23 29 30
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 3 11 10 19
rect 24 13 29 19
rect 31 13 36 30
rect 38 14 48 30
rect 38 13 42 14
rect 3 9 6 11
rect 8 9 10 11
rect 3 7 10 9
rect 40 12 42 13
rect 44 12 48 14
rect 40 10 48 12
rect 50 10 55 30
rect 57 23 62 30
rect 57 21 64 23
rect 57 19 60 21
rect 62 19 64 21
rect 57 17 64 19
rect 57 10 62 17
<< pdif >>
rect 2 65 9 67
rect 2 63 4 65
rect 6 63 9 65
rect 2 50 9 63
rect 11 61 19 67
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 50 19 52
rect 21 65 29 67
rect 21 63 24 65
rect 26 63 29 65
rect 21 50 29 63
rect 31 61 39 67
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 50 39 52
rect 41 65 49 67
rect 41 63 44 65
rect 46 63 49 65
rect 41 50 49 63
rect 43 42 49 50
rect 51 61 59 67
rect 51 59 54 61
rect 56 59 59 61
rect 51 54 59 59
rect 51 52 54 54
rect 56 52 59 54
rect 51 42 59 52
rect 61 65 69 67
rect 61 63 64 65
rect 66 63 69 65
rect 61 57 69 63
rect 61 55 64 57
rect 66 55 69 57
rect 61 42 69 55
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 13 61 17 63
rect 33 61 38 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 55 17 59
rect 2 54 17 55
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 2 52 14 54
rect 16 52 34 54
rect 36 52 38 54
rect 2 50 38 52
rect 2 22 6 50
rect 17 45 31 46
rect 17 43 27 45
rect 29 43 31 45
rect 17 42 31 43
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 50 41 62 47
rect 22 23 28 24
rect 22 22 24 23
rect 2 21 24 22
rect 26 21 28 23
rect 2 18 28 21
rect 50 25 54 41
rect 66 33 70 39
rect 68 31 70 33
rect 58 25 70 31
rect -2 11 74 12
rect -2 9 6 11
rect 8 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 12 19 14 30
rect 19 19 21 30
rect 29 13 31 30
rect 36 13 38 30
rect 48 10 50 30
rect 55 10 57 30
<< pmos >>
rect 9 50 11 67
rect 19 50 21 67
rect 29 50 31 67
rect 39 50 41 67
rect 49 42 51 67
rect 59 42 61 67
<< polyct0 >>
rect 11 35 13 37
rect 37 35 39 37
rect 47 35 49 37
<< polyct1 >>
rect 27 43 29 45
rect 27 35 29 37
rect 66 31 68 33
<< ndifct0 >>
rect 42 12 44 14
rect 60 19 62 21
<< ndifct1 >>
rect 24 21 26 23
rect 6 9 8 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 4 63 6 65
rect 24 63 26 65
rect 44 63 46 65
rect 54 59 56 61
rect 54 52 56 54
rect 64 63 66 65
rect 64 55 66 57
<< pdifct1 >>
rect 14 59 16 61
rect 14 52 16 54
rect 34 59 36 61
rect 34 52 36 54
<< alu0 >>
rect 3 65 7 68
rect 3 63 4 65
rect 6 63 7 65
rect 23 65 27 68
rect 23 63 24 65
rect 26 63 27 65
rect 43 65 47 68
rect 43 63 44 65
rect 46 63 47 65
rect 63 65 67 68
rect 63 63 64 65
rect 66 63 67 65
rect 3 61 7 63
rect 23 61 27 63
rect 43 61 47 63
rect 53 61 57 63
rect 53 59 54 61
rect 56 59 57 61
rect 53 54 57 59
rect 42 52 54 54
rect 56 52 57 54
rect 63 57 67 63
rect 63 55 64 57
rect 66 55 67 57
rect 63 53 67 55
rect 42 50 57 52
rect 42 46 46 50
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 31 14 35
rect 36 42 46 46
rect 36 37 40 42
rect 36 35 37 37
rect 39 35 40 37
rect 36 31 40 35
rect 45 37 50 38
rect 45 35 47 37
rect 49 35 50 37
rect 45 34 50 35
rect 10 27 40 31
rect 36 22 40 27
rect 65 31 66 35
rect 36 21 64 22
rect 36 19 60 21
rect 62 19 64 21
rect 36 18 64 19
rect 40 14 46 15
rect 40 12 42 14
rect 44 12 46 14
<< labels >>
rlabel alu0 12 33 12 33 6 an
rlabel alu0 38 32 38 32 6 an
rlabel alu0 50 20 50 20 6 an
rlabel alu0 55 56 55 56 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 44 20 44 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 52 36 52 36 6 a1
rlabel alu1 36 60 36 60 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 28 60 28 6 a2
rlabel alu1 68 32 68 32 6 a2
rlabel alu1 60 44 60 44 6 a1
<< end >>
