magic
tech scmos
timestamp 1199202699
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 10 57 16 59
rect 10 55 12 57
rect 14 55 16 57
rect 10 53 16 55
rect 10 50 12 53
rect 20 50 22 55
rect 10 35 12 38
rect 20 35 22 38
rect 9 32 12 35
rect 16 33 23 35
rect 9 26 11 32
rect 16 31 19 33
rect 21 31 23 33
rect 16 29 23 31
rect 16 26 18 29
rect 9 13 11 18
rect 16 13 18 18
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 20 9 22
rect 4 18 9 20
rect 11 18 16 26
rect 18 18 27 26
rect 20 17 27 18
rect 20 15 22 17
rect 24 15 27 17
rect 20 13 27 15
<< pdif >>
rect 2 65 8 67
rect 2 63 4 65
rect 6 63 8 65
rect 2 50 8 63
rect 2 38 10 50
rect 12 42 20 50
rect 12 40 15 42
rect 17 40 20 42
rect 12 38 20 40
rect 22 48 30 50
rect 22 46 26 48
rect 28 46 30 48
rect 22 38 30 46
<< alu1 >>
rect -2 67 34 72
rect -2 65 17 67
rect 19 65 25 67
rect 27 65 34 67
rect -2 64 4 65
rect 6 64 34 65
rect 9 57 23 58
rect 9 55 12 57
rect 14 55 23 57
rect 9 54 23 55
rect 9 46 15 54
rect 2 40 15 42
rect 17 40 19 42
rect 2 38 19 40
rect 2 26 6 38
rect 17 33 23 34
rect 17 31 19 33
rect 21 31 23 33
rect 17 27 23 31
rect 2 24 7 26
rect 2 22 4 24
rect 6 22 7 24
rect 2 20 7 22
rect 17 21 30 27
rect -2 7 34 8
rect -2 5 5 7
rect 7 5 25 7
rect 27 5 34 7
rect -2 0 34 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 23 7 29 9
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< ntie >>
rect 15 67 29 69
rect 15 65 17 67
rect 19 65 25 67
rect 27 65 29 67
rect 15 63 29 65
<< nmos >>
rect 9 18 11 26
rect 16 18 18 26
<< pmos >>
rect 10 38 12 50
rect 20 38 22 50
<< polyct1 >>
rect 12 55 14 57
rect 19 31 21 33
<< ndifct0 >>
rect 22 15 24 17
<< ndifct1 >>
rect 4 22 6 24
<< ntiect1 >>
rect 17 65 19 67
rect 25 65 27 67
<< ptiect1 >>
rect 5 5 7 7
rect 25 5 27 7
<< pdifct0 >>
rect 4 63 6 64
rect 26 46 28 48
<< pdifct1 >>
rect 4 64 6 65
rect 15 40 17 42
<< alu0 >>
rect 2 63 4 64
rect 6 63 8 64
rect 2 62 8 63
rect 26 49 30 64
rect 24 48 30 49
rect 24 46 26 48
rect 28 46 30 48
rect 24 45 30 46
rect 13 42 19 43
rect 20 17 26 18
rect 20 15 22 17
rect 24 15 26 17
rect 20 8 26 15
<< labels >>
rlabel alu1 4 28 4 28 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 12 52 12 52 6 b
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 28 20 28 6 a
rlabel alu1 20 56 20 56 6 b
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 24 28 24 6 a
<< end >>
