magic
tech scmos
timestamp 1199202540
<< ab >>
rect 0 0 96 80
<< nwell >>
rect -5 36 101 88
<< pwell >>
rect -5 -8 101 36
<< poly >>
rect 29 70 31 74
rect 39 70 41 74
rect 9 65 11 70
rect 19 65 21 70
rect 9 47 11 50
rect 19 47 21 50
rect 9 45 21 47
rect 9 43 11 45
rect 13 43 15 45
rect 9 41 15 43
rect 51 70 53 74
rect 61 70 63 74
rect 71 70 73 74
rect 81 60 83 65
rect 71 47 73 50
rect 81 47 83 50
rect 71 45 83 47
rect 71 43 75 45
rect 77 43 83 45
rect 9 28 11 41
rect 29 37 31 42
rect 15 35 31 37
rect 39 39 41 42
rect 51 39 53 42
rect 61 39 63 42
rect 71 41 83 43
rect 39 37 53 39
rect 57 37 63 39
rect 39 35 45 37
rect 47 35 49 37
rect 15 33 17 35
rect 19 33 21 35
rect 15 31 21 33
rect 29 28 31 35
rect 36 33 49 35
rect 57 35 59 37
rect 61 35 63 37
rect 57 33 63 35
rect 71 35 77 37
rect 71 33 73 35
rect 75 33 77 35
rect 36 28 38 33
rect 47 28 49 33
rect 54 31 66 33
rect 54 28 56 31
rect 64 28 66 31
rect 71 31 77 33
rect 71 28 73 31
rect 81 28 83 41
rect 9 8 11 13
rect 29 6 31 10
rect 36 6 38 10
rect 47 8 49 13
rect 54 8 56 13
rect 64 8 66 13
rect 71 8 73 13
rect 81 8 83 13
<< ndif >>
rect 2 26 9 28
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 4 13 9 22
rect 11 25 18 28
rect 11 23 14 25
rect 16 23 18 25
rect 11 17 18 23
rect 22 26 29 28
rect 22 24 24 26
rect 26 24 29 26
rect 22 22 29 24
rect 11 15 14 17
rect 16 15 18 17
rect 11 13 18 15
rect 24 10 29 22
rect 31 10 36 28
rect 38 14 47 28
rect 38 12 41 14
rect 43 13 47 14
rect 49 13 54 28
rect 56 21 64 28
rect 56 19 59 21
rect 61 19 64 21
rect 56 13 64 19
rect 66 13 71 28
rect 73 17 81 28
rect 73 15 76 17
rect 78 15 81 17
rect 73 13 81 15
rect 83 26 90 28
rect 83 24 86 26
rect 88 24 90 26
rect 83 22 90 24
rect 83 13 88 22
rect 43 12 45 13
rect 38 10 45 12
<< pdif >>
rect 43 71 49 73
rect 43 70 45 71
rect 23 65 29 70
rect 2 63 9 65
rect 2 61 4 63
rect 6 61 9 63
rect 2 50 9 61
rect 11 61 19 65
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 50 19 52
rect 21 63 29 65
rect 21 61 24 63
rect 26 61 29 63
rect 21 50 29 61
rect 23 42 29 50
rect 31 62 39 70
rect 31 60 34 62
rect 36 60 39 62
rect 31 46 39 60
rect 31 44 34 46
rect 36 44 39 46
rect 31 42 39 44
rect 41 69 45 70
rect 47 70 49 71
rect 47 69 51 70
rect 41 42 51 69
rect 53 62 61 70
rect 53 60 56 62
rect 58 60 61 62
rect 53 55 61 60
rect 53 53 56 55
rect 58 53 61 55
rect 53 42 61 53
rect 63 68 71 70
rect 63 66 66 68
rect 68 66 71 68
rect 63 61 71 66
rect 63 59 66 61
rect 68 59 71 61
rect 63 50 71 59
rect 73 60 78 70
rect 73 54 81 60
rect 73 52 76 54
rect 78 52 81 54
rect 73 50 81 52
rect 83 58 90 60
rect 83 56 86 58
rect 88 56 90 58
rect 83 50 90 56
rect 63 42 69 50
<< alu1 >>
rect -2 81 98 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 98 81
rect -2 71 98 79
rect -2 69 45 71
rect 47 69 98 71
rect -2 68 98 69
rect 2 47 6 55
rect 2 45 14 47
rect 2 43 11 45
rect 13 43 14 45
rect 2 41 14 43
rect 26 46 39 47
rect 26 44 34 46
rect 36 44 39 46
rect 26 42 39 44
rect 26 22 30 42
rect 74 45 86 47
rect 74 43 75 45
rect 77 43 86 45
rect 74 41 86 43
rect 82 33 86 41
rect 26 21 63 22
rect 26 19 59 21
rect 61 19 63 21
rect 26 18 63 19
rect -2 1 98 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 98 1
rect -2 -2 98 -1
<< ptie >>
rect 0 1 96 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 96 1
rect 0 -3 96 -1
<< ntie >>
rect 0 81 96 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 96 81
rect 0 77 96 79
<< nmos >>
rect 9 13 11 28
rect 29 10 31 28
rect 36 10 38 28
rect 47 13 49 28
rect 54 13 56 28
rect 64 13 66 28
rect 71 13 73 28
rect 81 13 83 28
<< pmos >>
rect 9 50 11 65
rect 19 50 21 65
rect 29 42 31 70
rect 39 42 41 70
rect 51 42 53 70
rect 61 42 63 70
rect 71 50 73 70
rect 81 50 83 60
<< polyct0 >>
rect 45 35 47 37
rect 17 33 19 35
rect 59 35 61 37
rect 73 33 75 35
<< polyct1 >>
rect 11 43 13 45
rect 75 43 77 45
<< ndifct0 >>
rect 4 24 6 26
rect 14 23 16 25
rect 24 24 26 26
rect 14 15 16 17
rect 41 12 43 14
rect 76 15 78 17
rect 86 24 88 26
<< ndifct1 >>
rect 59 19 61 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
<< pdifct0 >>
rect 4 61 6 63
rect 14 59 16 61
rect 14 52 16 54
rect 24 61 26 63
rect 34 60 36 62
rect 56 60 58 62
rect 56 53 58 55
rect 66 66 68 68
rect 66 59 68 61
rect 76 52 78 54
rect 86 56 88 58
<< pdifct1 >>
rect 34 44 36 46
rect 45 69 47 71
<< alu0 >>
rect 3 63 7 68
rect 23 63 27 68
rect 64 66 66 68
rect 68 66 70 68
rect 3 61 4 63
rect 6 61 7 63
rect 3 59 7 61
rect 12 61 17 63
rect 12 59 14 61
rect 16 59 17 61
rect 23 61 24 63
rect 26 61 27 63
rect 23 59 27 61
rect 32 62 60 63
rect 32 60 34 62
rect 36 60 56 62
rect 58 60 60 62
rect 32 59 60 60
rect 12 55 17 59
rect 55 55 60 59
rect 64 61 70 66
rect 64 59 66 61
rect 68 59 70 61
rect 64 58 70 59
rect 85 58 89 68
rect 85 56 86 58
rect 88 56 89 58
rect 12 54 49 55
rect 12 52 14 54
rect 16 52 49 54
rect 12 51 49 52
rect 55 53 56 55
rect 58 53 60 55
rect 55 51 60 53
rect 67 54 80 55
rect 85 54 89 56
rect 67 52 76 54
rect 78 52 80 54
rect 67 51 80 52
rect 18 36 22 51
rect 45 47 49 51
rect 3 35 22 36
rect 3 33 17 35
rect 19 33 22 35
rect 3 32 22 33
rect 45 43 62 47
rect 3 26 7 32
rect 3 24 4 26
rect 6 24 7 26
rect 3 22 7 24
rect 13 25 17 27
rect 13 23 14 25
rect 16 23 17 25
rect 22 26 26 27
rect 22 24 24 26
rect 22 23 26 24
rect 13 17 17 23
rect 43 37 52 38
rect 43 35 45 37
rect 47 35 52 37
rect 43 34 52 35
rect 48 29 52 34
rect 58 37 62 43
rect 58 35 59 37
rect 61 35 62 37
rect 58 33 62 35
rect 67 36 71 51
rect 67 35 77 36
rect 67 33 73 35
rect 75 33 77 35
rect 67 32 77 33
rect 67 29 71 32
rect 48 27 71 29
rect 48 26 90 27
rect 48 25 86 26
rect 67 24 86 25
rect 88 24 90 26
rect 67 23 90 24
rect 13 15 14 17
rect 16 15 17 17
rect 75 17 79 19
rect 75 15 76 17
rect 78 15 79 17
rect 13 12 17 15
rect 39 14 45 15
rect 39 12 41 14
rect 43 12 45 14
rect 75 12 79 15
<< labels >>
rlabel alu0 5 29 5 29 6 bn
rlabel alu0 12 34 12 34 6 bn
rlabel alu0 14 57 14 57 6 bn
rlabel alu0 47 36 47 36 6 an
rlabel alu0 60 40 60 40 6 bn
rlabel alu0 30 53 30 53 6 bn
rlabel alu0 72 34 72 34 6 an
rlabel alu0 78 25 78 25 6 an
rlabel alu0 73 53 73 53 6 an
rlabel polyct1 12 44 12 44 6 b
rlabel alu1 4 48 4 48 6 b
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 36 28 36 6 z
rlabel alu1 36 44 36 44 6 z
rlabel alu1 48 6 48 6 6 vss
rlabel ndifct1 60 20 60 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 48 74 48 74 6 vdd
rlabel alu1 84 40 84 40 6 a
rlabel polyct1 76 44 76 44 6 a
<< end >>
