magic
tech scmos
timestamp 1199202970
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 9 34 11 43
rect 16 40 18 43
rect 26 40 28 43
rect 33 40 35 43
rect 43 40 45 43
rect 16 38 29 40
rect 33 38 45 40
rect 50 39 52 43
rect 60 39 62 43
rect 23 37 29 38
rect 23 35 25 37
rect 27 35 29 37
rect 9 32 19 34
rect 13 30 15 32
rect 17 30 19 32
rect 13 28 19 30
rect 23 33 29 35
rect 36 36 42 38
rect 36 34 38 36
rect 40 34 42 36
rect 50 37 62 39
rect 67 38 69 43
rect 50 35 52 37
rect 54 35 62 37
rect 50 34 62 35
rect 13 25 15 28
rect 23 25 25 33
rect 36 32 42 34
rect 47 32 62 34
rect 66 36 72 38
rect 66 34 68 36
rect 70 34 72 36
rect 66 32 72 34
rect 37 29 39 32
rect 47 29 49 32
rect 59 29 61 32
rect 69 29 71 32
rect 13 6 15 10
rect 23 6 25 10
rect 37 6 39 10
rect 47 6 49 10
rect 59 6 61 10
rect 69 6 71 10
<< ndif >>
rect 27 25 37 29
rect 4 14 13 25
rect 4 12 8 14
rect 10 12 13 14
rect 4 10 13 12
rect 15 21 23 25
rect 15 19 18 21
rect 20 19 23 21
rect 15 10 23 19
rect 25 14 37 25
rect 25 12 30 14
rect 32 12 37 14
rect 25 10 37 12
rect 39 21 47 29
rect 39 19 42 21
rect 44 19 47 21
rect 39 10 47 19
rect 49 14 59 29
rect 49 12 53 14
rect 55 12 59 14
rect 49 10 59 12
rect 61 21 69 29
rect 61 19 64 21
rect 66 19 69 21
rect 61 10 69 19
rect 71 21 78 29
rect 71 19 74 21
rect 76 19 78 21
rect 71 14 78 19
rect 71 12 74 14
rect 76 12 78 14
rect 71 10 78 12
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 43 9 59
rect 11 43 16 70
rect 18 55 26 70
rect 18 53 21 55
rect 23 53 26 55
rect 18 47 26 53
rect 18 45 21 47
rect 23 45 26 47
rect 18 43 26 45
rect 28 43 33 70
rect 35 68 43 70
rect 35 66 38 68
rect 40 66 43 68
rect 35 61 43 66
rect 35 59 38 61
rect 40 59 43 61
rect 35 43 43 59
rect 45 43 50 70
rect 52 55 60 70
rect 52 53 55 55
rect 57 53 60 55
rect 52 47 60 53
rect 52 45 55 47
rect 57 45 60 47
rect 52 43 60 45
rect 62 43 67 70
rect 69 68 77 70
rect 69 66 72 68
rect 74 66 77 68
rect 69 61 77 66
rect 69 59 72 61
rect 74 59 77 61
rect 69 43 77 59
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 18 55 24 57
rect 18 53 21 55
rect 23 54 24 55
rect 23 53 55 54
rect 57 53 63 54
rect 18 50 63 53
rect 18 47 24 50
rect 2 45 21 47
rect 23 45 24 47
rect 2 42 24 45
rect 29 42 49 46
rect 2 22 6 42
rect 29 38 33 42
rect 45 38 49 42
rect 23 37 33 38
rect 23 35 25 37
rect 27 35 33 37
rect 23 34 33 35
rect 45 37 56 38
rect 45 35 52 37
rect 54 35 56 37
rect 45 34 56 35
rect 65 36 71 38
rect 65 34 68 36
rect 70 34 71 36
rect 14 32 18 34
rect 14 30 15 32
rect 17 30 18 32
rect 65 30 71 34
rect 14 26 71 30
rect 2 21 68 22
rect 2 19 18 21
rect 20 19 42 21
rect 44 19 64 21
rect 66 19 68 21
rect 2 18 68 19
rect -2 1 82 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 13 10 15 25
rect 23 10 25 25
rect 37 10 39 29
rect 47 10 49 29
rect 59 10 61 29
rect 69 10 71 29
<< pmos >>
rect 9 43 11 70
rect 16 43 18 70
rect 26 43 28 70
rect 33 43 35 70
rect 43 43 45 70
rect 50 43 52 70
rect 60 43 62 70
rect 67 43 69 70
<< polyct0 >>
rect 38 34 40 36
<< polyct1 >>
rect 25 35 27 37
rect 15 30 17 32
rect 52 35 54 37
rect 68 34 70 36
<< ndifct0 >>
rect 8 12 10 14
rect 30 12 32 14
rect 53 12 55 14
rect 74 19 76 21
rect 74 12 76 14
<< ndifct1 >>
rect 18 19 20 21
rect 42 19 44 21
rect 64 19 66 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 38 66 40 68
rect 38 59 40 61
rect 55 54 57 55
rect 55 45 57 47
rect 72 66 74 68
rect 72 59 74 61
<< pdifct1 >>
rect 21 53 23 55
rect 21 45 23 47
rect 55 53 57 54
<< alu0 >>
rect 2 66 4 68
rect 6 66 8 68
rect 2 61 8 66
rect 2 59 4 61
rect 6 59 8 61
rect 2 58 8 59
rect 36 66 38 68
rect 40 66 42 68
rect 36 61 42 66
rect 36 59 38 61
rect 40 59 42 61
rect 36 58 42 59
rect 70 66 72 68
rect 74 66 76 68
rect 70 61 76 66
rect 70 59 72 61
rect 74 59 76 61
rect 70 58 76 59
rect 54 55 58 57
rect 54 54 55 55
rect 57 54 58 55
rect 54 47 58 50
rect 54 45 55 47
rect 57 45 58 47
rect 54 43 58 45
rect 37 36 41 38
rect 37 34 38 36
rect 40 34 41 36
rect 37 30 41 34
rect 72 21 78 22
rect 72 19 74 21
rect 76 19 78 21
rect 6 14 12 15
rect 6 12 8 14
rect 10 12 12 14
rect 28 14 34 15
rect 28 12 30 14
rect 32 12 34 14
rect 51 14 57 15
rect 51 12 53 14
rect 55 12 57 14
rect 72 14 78 19
rect 72 12 74 14
rect 76 12 78 14
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 12 44 12 44 6 z
rlabel alu1 28 36 28 36 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 20 44 20 6 z
rlabel alu1 44 28 44 28 6 a
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 44 44 44 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 52 20 52 20 6 z
rlabel alu1 52 28 52 28 6 a
rlabel alu1 60 20 60 20 6 z
rlabel alu1 60 28 60 28 6 a
rlabel alu1 52 36 52 36 6 b
rlabel alu1 60 52 60 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 68 32 68 32 6 a
<< end >>
