magic
tech scmos
timestamp 1199542480
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 11 95 13 98
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 11 43 13 55
rect 23 43 25 55
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 25 43
rect 17 39 19 41
rect 21 39 25 41
rect 17 37 25 39
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 55
rect 47 43 49 55
rect 35 41 43 43
rect 35 39 39 41
rect 41 39 43 41
rect 35 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 35 25 37 37
rect 47 25 49 37
rect 11 2 13 5
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
<< ndif >>
rect 15 31 21 33
rect 15 29 17 31
rect 19 29 21 31
rect 15 25 21 29
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 5 11 19
rect 13 5 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 5 35 19
rect 37 11 47 25
rect 37 9 41 11
rect 43 9 47 11
rect 37 5 47 9
rect 49 21 57 25
rect 49 19 53 21
rect 55 19 57 21
rect 49 5 57 19
<< pdif >>
rect 3 91 11 95
rect 3 89 5 91
rect 7 89 11 91
rect 3 55 11 89
rect 13 55 23 95
rect 25 81 35 95
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 61 35 69
rect 25 59 29 61
rect 31 59 35 61
rect 25 55 35 59
rect 37 55 47 95
rect 49 91 57 95
rect 49 89 53 91
rect 55 89 57 91
rect 49 73 57 89
rect 49 55 55 73
<< alu1 >>
rect -2 91 72 100
rect -2 89 5 91
rect 7 89 53 91
rect 55 89 72 91
rect -2 88 72 89
rect 8 41 12 82
rect 8 39 9 41
rect 11 39 12 41
rect 8 38 12 39
rect 18 41 22 82
rect 18 39 19 41
rect 21 39 22 41
rect 18 38 22 39
rect 28 81 32 82
rect 28 79 29 81
rect 31 79 32 81
rect 28 71 32 79
rect 28 69 29 71
rect 31 69 32 71
rect 28 61 32 69
rect 28 59 29 61
rect 31 59 32 61
rect 28 32 32 59
rect 16 31 32 32
rect 16 29 17 31
rect 19 29 32 31
rect 16 28 32 29
rect 38 41 42 82
rect 38 39 39 41
rect 41 39 42 41
rect 38 28 42 39
rect 48 41 52 82
rect 62 59 66 88
rect 62 57 63 59
rect 65 57 66 59
rect 62 56 66 57
rect 48 39 49 41
rect 51 39 52 41
rect 48 28 52 39
rect 4 21 8 22
rect 28 21 32 22
rect 52 21 56 22
rect 4 19 5 21
rect 7 19 29 21
rect 31 19 53 21
rect 55 19 56 21
rect 4 18 8 19
rect 28 18 32 19
rect 52 18 56 19
rect -2 11 72 12
rect -2 9 41 11
rect 43 9 72 11
rect -2 0 72 9
<< ntie >>
rect 61 59 67 67
rect 61 57 63 59
rect 65 57 67 59
rect 61 55 67 57
<< nmos >>
rect 11 5 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
<< pmos >>
rect 11 55 13 95
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 39 39 41 41
rect 49 39 51 41
<< ndifct1 >>
rect 17 29 19 31
rect 5 19 7 21
rect 29 19 31 21
rect 41 9 43 11
rect 53 19 55 21
<< ntiect1 >>
rect 63 57 65 59
<< pdifct1 >>
rect 5 89 7 91
rect 29 79 31 81
rect 29 69 31 71
rect 29 59 31 61
rect 53 89 55 91
<< labels >>
rlabel alu1 10 60 10 60 6 i0
rlabel alu1 30 55 30 55 6 nq
rlabel alu1 20 60 20 60 6 i1
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 50 55 50 55 6 i2
rlabel alu1 40 55 40 55 6 i3
rlabel alu1 35 94 35 94 6 vdd
<< end >>
