magic
tech scmos
timestamp 1199468882
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -2 48 52 104
<< pwell >>
rect -2 -4 52 48
<< poly >>
rect 13 78 15 83
rect 25 74 27 79
rect 37 74 39 79
rect 13 47 15 58
rect 25 54 27 58
rect 25 52 33 54
rect 25 51 29 52
rect 27 50 29 51
rect 31 50 33 52
rect 27 48 33 50
rect 37 53 39 58
rect 37 51 43 53
rect 37 49 39 51
rect 41 49 43 51
rect 13 45 23 47
rect 13 43 19 45
rect 21 43 23 45
rect 13 41 23 43
rect 15 38 17 41
rect 29 31 31 48
rect 37 47 43 49
rect 37 31 39 47
rect 15 23 17 28
rect 29 12 31 17
rect 37 12 39 17
<< ndif >>
rect 7 36 15 38
rect 7 34 9 36
rect 11 34 15 36
rect 7 32 15 34
rect 10 28 15 32
rect 17 31 27 38
rect 17 28 29 31
rect 19 21 29 28
rect 19 19 22 21
rect 24 19 29 21
rect 19 17 29 19
rect 31 17 37 31
rect 39 29 47 31
rect 39 27 43 29
rect 45 27 47 29
rect 39 21 47 27
rect 39 19 43 21
rect 45 19 47 21
rect 39 17 47 19
<< pdif >>
rect 17 81 23 83
rect 17 79 19 81
rect 21 79 23 81
rect 41 81 47 83
rect 41 79 43 81
rect 45 79 47 81
rect 17 78 23 79
rect 8 72 13 78
rect 5 70 13 72
rect 5 68 7 70
rect 9 68 13 70
rect 5 62 13 68
rect 5 60 7 62
rect 9 60 13 62
rect 5 58 13 60
rect 15 74 23 78
rect 41 74 47 79
rect 15 58 25 74
rect 27 62 37 74
rect 27 60 31 62
rect 33 60 37 62
rect 27 58 37 60
rect 39 58 47 74
<< alu1 >>
rect -2 95 52 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 52 95
rect -2 88 52 93
rect 18 81 22 88
rect 18 79 19 81
rect 21 79 22 81
rect 18 77 22 79
rect 42 81 46 88
rect 42 79 43 81
rect 45 79 46 81
rect 42 77 46 79
rect 6 70 23 72
rect 6 68 7 70
rect 9 68 23 70
rect 27 68 42 73
rect 6 62 12 68
rect 6 60 7 62
rect 9 60 12 62
rect 6 58 12 60
rect 8 36 12 58
rect 8 34 9 36
rect 11 34 12 36
rect 8 32 12 34
rect 18 62 34 64
rect 18 60 31 62
rect 33 60 34 62
rect 18 58 34 60
rect 18 45 22 58
rect 18 43 19 45
rect 21 43 22 45
rect 18 30 22 43
rect 28 52 32 54
rect 28 50 29 52
rect 31 50 32 52
rect 28 42 32 50
rect 38 51 42 68
rect 38 49 39 51
rect 41 49 42 51
rect 38 47 42 49
rect 28 37 43 42
rect 18 29 47 30
rect 18 27 43 29
rect 45 27 47 29
rect 18 26 47 27
rect 20 21 26 22
rect 20 19 22 21
rect 24 19 26 21
rect 20 12 26 19
rect 41 21 47 26
rect 41 19 43 21
rect 45 19 47 21
rect 41 18 47 19
rect -2 7 52 12
rect -2 5 9 7
rect 11 5 17 7
rect 19 5 52 7
rect -2 0 52 5
<< ptie >>
rect 7 7 21 9
rect 7 5 9 7
rect 11 5 17 7
rect 19 5 21 7
rect 7 3 21 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 15 28 17 38
rect 29 17 31 31
rect 37 17 39 31
<< pmos >>
rect 13 58 15 78
rect 25 58 27 74
rect 37 58 39 74
<< polyct1 >>
rect 29 50 31 52
rect 39 49 41 51
rect 19 43 21 45
<< ndifct1 >>
rect 9 34 11 36
rect 22 19 24 21
rect 43 27 45 29
rect 43 19 45 21
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 9 5 11 7
rect 17 5 19 7
<< pdifct1 >>
rect 19 79 21 81
rect 43 79 45 81
rect 7 68 9 70
rect 7 60 9 62
rect 31 60 33 62
<< labels >>
rlabel alu1 20 45 20 45 6 zn
rlabel alu1 10 55 10 55 6 z
rlabel alu1 20 70 20 70 6 z
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 45 30 45 6 a
rlabel alu1 26 61 26 61 6 zn
rlabel alu1 30 70 30 70 6 b
rlabel alu1 25 94 25 94 6 vdd
rlabel alu1 44 24 44 24 6 zn
rlabel alu1 32 28 32 28 6 zn
rlabel alu1 40 40 40 40 6 a
rlabel alu1 40 60 40 60 6 b
<< end >>
