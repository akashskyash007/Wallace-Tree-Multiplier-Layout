magic
tech scmos
timestamp 1199470545
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -2 48 82 104
<< pwell >>
rect -2 -4 82 48
<< poly >>
rect 47 87 49 92
rect 55 87 57 92
rect 67 87 69 92
rect 11 75 13 80
rect 31 82 37 84
rect 31 80 33 82
rect 35 80 37 82
rect 23 75 25 80
rect 31 78 37 80
rect 35 75 37 78
rect 11 38 13 55
rect 23 46 25 55
rect 35 50 37 55
rect 47 53 49 67
rect 55 63 57 67
rect 67 63 69 67
rect 53 61 59 63
rect 53 59 55 61
rect 57 59 59 61
rect 53 57 59 59
rect 63 61 69 63
rect 63 59 65 61
rect 67 59 69 61
rect 63 57 69 59
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 47 46 49 47
rect 23 44 33 46
rect 27 42 29 44
rect 31 42 33 44
rect 27 40 33 42
rect 41 44 49 46
rect 11 36 23 38
rect 17 34 19 36
rect 21 34 23 36
rect 17 32 23 34
rect 21 29 23 32
rect 29 29 31 40
rect 41 29 43 44
rect 57 31 59 57
rect 53 29 59 31
rect 53 26 55 29
rect 65 26 67 57
rect 21 12 23 17
rect 29 12 31 17
rect 41 12 43 17
rect 53 12 55 17
rect 65 12 67 17
<< ndif >>
rect 12 17 21 29
rect 23 17 29 29
rect 31 21 41 29
rect 31 19 35 21
rect 37 19 41 21
rect 31 17 41 19
rect 43 26 48 29
rect 43 21 53 26
rect 43 19 47 21
rect 49 19 53 21
rect 43 17 53 19
rect 55 21 65 26
rect 55 19 59 21
rect 61 19 65 21
rect 55 17 65 19
rect 67 21 76 26
rect 67 19 71 21
rect 73 19 76 21
rect 67 17 76 19
rect 12 11 19 17
rect 12 9 15 11
rect 17 9 19 11
rect 12 7 19 9
<< pdif >>
rect 59 91 65 93
rect 59 89 61 91
rect 63 89 65 91
rect 59 87 65 89
rect 15 81 21 83
rect 15 79 17 81
rect 19 79 21 81
rect 15 75 21 79
rect 42 75 47 87
rect 6 69 11 75
rect 3 67 11 69
rect 3 65 5 67
rect 7 65 11 67
rect 3 59 11 65
rect 3 57 5 59
rect 7 57 11 59
rect 3 55 11 57
rect 13 55 23 75
rect 25 71 35 75
rect 25 69 29 71
rect 31 69 35 71
rect 25 55 35 69
rect 37 67 47 75
rect 49 67 55 87
rect 57 67 67 87
rect 69 81 74 87
rect 69 79 77 81
rect 69 77 73 79
rect 75 77 77 79
rect 69 71 77 77
rect 69 69 73 71
rect 75 69 77 71
rect 69 67 77 69
rect 37 61 45 67
rect 37 59 41 61
rect 43 59 45 61
rect 37 57 45 59
rect 37 55 42 57
<< alu1 >>
rect -2 95 82 100
rect -2 93 9 95
rect 11 93 19 95
rect 21 93 82 95
rect -2 91 82 93
rect -2 89 61 91
rect 63 89 82 91
rect -2 88 82 89
rect 16 81 20 88
rect 16 79 17 81
rect 19 79 20 81
rect 16 77 20 79
rect 31 82 62 83
rect 31 80 33 82
rect 35 80 62 82
rect 31 78 62 80
rect 4 71 52 72
rect 4 69 29 71
rect 31 69 52 71
rect 4 68 52 69
rect 4 67 8 68
rect 4 65 5 67
rect 7 65 8 67
rect 4 59 8 65
rect 4 57 5 59
rect 7 57 8 59
rect 18 57 32 63
rect 4 22 8 57
rect 18 36 22 53
rect 28 44 32 57
rect 28 42 29 44
rect 31 42 32 44
rect 28 37 32 42
rect 38 61 44 63
rect 38 59 41 61
rect 43 59 44 61
rect 38 43 44 59
rect 48 62 52 68
rect 58 71 62 78
rect 72 79 76 81
rect 72 77 73 79
rect 75 77 76 79
rect 72 71 76 77
rect 58 67 68 71
rect 48 61 59 62
rect 48 59 55 61
rect 57 59 59 61
rect 48 58 59 59
rect 64 61 68 67
rect 64 59 65 61
rect 67 59 68 61
rect 64 57 68 59
rect 72 69 73 71
rect 75 69 76 71
rect 72 53 76 69
rect 48 51 76 53
rect 48 49 49 51
rect 51 49 76 51
rect 48 47 62 49
rect 38 37 52 43
rect 18 34 19 36
rect 21 34 22 36
rect 18 33 22 34
rect 18 27 42 33
rect 4 21 39 22
rect 4 19 35 21
rect 37 19 39 21
rect 4 18 39 19
rect 46 21 52 37
rect 46 19 47 21
rect 49 19 52 21
rect 46 17 52 19
rect 58 21 62 47
rect 58 19 59 21
rect 61 19 62 21
rect 58 17 62 19
rect 70 21 74 23
rect 70 19 71 21
rect 73 19 74 21
rect 70 12 74 19
rect -2 11 82 12
rect -2 9 15 11
rect 17 9 82 11
rect -2 7 82 9
rect -2 5 29 7
rect 31 5 39 7
rect 41 5 82 7
rect -2 0 82 5
<< ptie >>
rect 27 7 43 9
rect 27 5 29 7
rect 31 5 39 7
rect 41 5 43 7
rect 27 3 43 5
<< ntie >>
rect 7 95 23 97
rect 7 93 9 95
rect 11 93 19 95
rect 21 93 23 95
rect 7 91 23 93
<< nmos >>
rect 21 17 23 29
rect 29 17 31 29
rect 41 17 43 29
rect 53 17 55 26
rect 65 17 67 26
<< pmos >>
rect 11 55 13 75
rect 23 55 25 75
rect 35 55 37 75
rect 47 67 49 87
rect 55 67 57 87
rect 67 67 69 87
<< polyct1 >>
rect 33 80 35 82
rect 55 59 57 61
rect 65 59 67 61
rect 49 49 51 51
rect 29 42 31 44
rect 19 34 21 36
<< ndifct1 >>
rect 35 19 37 21
rect 47 19 49 21
rect 59 19 61 21
rect 71 19 73 21
rect 15 9 17 11
<< ntiect1 >>
rect 9 93 11 95
rect 19 93 21 95
<< ptiect1 >>
rect 29 5 31 7
rect 39 5 41 7
<< pdifct1 >>
rect 61 89 63 91
rect 17 79 19 81
rect 5 65 7 67
rect 5 57 7 59
rect 29 69 31 71
rect 73 77 75 79
rect 73 69 75 71
rect 41 59 43 61
<< labels >>
rlabel alu1 6 45 6 45 6 an
rlabel alu1 20 40 20 40 6 a1
rlabel alu1 20 60 20 60 6 a2
rlabel ptiect1 40 6 40 6 6 vss
rlabel alu1 21 20 21 20 6 an
rlabel alu1 30 30 30 30 6 a1
rlabel alu1 40 30 40 30 6 a1
rlabel alu1 30 50 30 50 6 a2
rlabel alu1 40 50 40 50 6 z
rlabel alu1 40 80 40 80 6 b
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 50 30 50 30 6 z
rlabel alu1 60 35 60 35 6 bn
rlabel alu1 53 60 53 60 6 an
rlabel alu1 28 70 28 70 6 an
rlabel alu1 60 75 60 75 6 b
rlabel alu1 50 80 50 80 6 b
rlabel alu1 62 51 62 51 6 bn
rlabel alu1 74 65 74 65 6 bn
<< end >>
