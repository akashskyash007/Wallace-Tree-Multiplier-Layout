magic
tech scmos
timestamp 1199542838
<< ab >>
rect 0 0 100 100
<< nwell >>
rect -2 48 102 104
<< pwell >>
rect -2 -4 102 48
<< poly >>
rect 73 95 75 98
rect 85 95 87 98
rect 13 85 15 88
rect 25 85 27 88
rect 37 85 39 88
rect 61 75 63 78
rect 13 43 15 65
rect 7 41 15 43
rect 7 39 9 41
rect 11 39 15 41
rect 7 37 15 39
rect 13 25 15 37
rect 25 43 27 65
rect 37 43 39 65
rect 61 53 63 55
rect 61 51 69 53
rect 61 49 65 51
rect 67 49 69 51
rect 61 47 69 49
rect 25 41 33 43
rect 25 39 29 41
rect 31 39 33 41
rect 25 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 25 25 27 37
rect 37 25 39 37
rect 61 25 63 47
rect 73 43 75 55
rect 85 43 87 55
rect 67 41 87 43
rect 67 39 69 41
rect 71 39 87 41
rect 67 37 87 39
rect 73 25 75 37
rect 85 25 87 37
rect 13 12 15 15
rect 25 12 27 15
rect 37 12 39 15
rect 61 12 63 15
rect 73 2 75 5
rect 85 2 87 5
<< ndif >>
rect 5 15 13 25
rect 15 21 25 25
rect 15 19 19 21
rect 21 19 25 21
rect 15 15 25 19
rect 27 15 37 25
rect 39 15 47 25
rect 53 21 61 25
rect 53 19 55 21
rect 57 19 61 21
rect 53 15 61 19
rect 63 21 73 25
rect 63 19 67 21
rect 69 19 73 21
rect 63 15 73 19
rect 5 11 11 15
rect 5 9 7 11
rect 9 9 11 11
rect 41 11 47 15
rect 41 9 43 11
rect 45 9 47 11
rect 5 7 11 9
rect 41 7 47 9
rect 65 11 73 15
rect 65 9 67 11
rect 69 9 73 11
rect 65 5 73 9
rect 75 21 85 25
rect 75 19 79 21
rect 81 19 85 21
rect 75 5 85 19
rect 87 21 95 25
rect 87 19 91 21
rect 93 19 95 21
rect 87 11 95 19
rect 87 9 91 11
rect 93 9 95 11
rect 87 5 95 9
<< pdif >>
rect 5 91 11 93
rect 65 91 73 95
rect 5 89 7 91
rect 9 89 11 91
rect 5 85 11 89
rect 65 89 67 91
rect 69 89 73 91
rect 5 65 13 85
rect 15 81 25 85
rect 15 79 19 81
rect 21 79 25 81
rect 15 65 25 79
rect 27 71 37 85
rect 27 69 31 71
rect 33 69 37 71
rect 27 65 37 69
rect 39 81 47 85
rect 39 79 43 81
rect 45 79 47 81
rect 39 65 47 79
rect 65 81 73 89
rect 65 79 67 81
rect 69 79 73 81
rect 65 75 73 79
rect 53 61 61 75
rect 53 59 55 61
rect 57 59 61 61
rect 53 55 61 59
rect 63 55 73 75
rect 75 81 85 95
rect 75 79 79 81
rect 81 79 85 81
rect 75 71 85 79
rect 75 69 79 71
rect 81 69 85 71
rect 75 61 85 69
rect 75 59 79 61
rect 81 59 85 61
rect 75 55 85 59
rect 87 91 95 95
rect 87 89 91 91
rect 93 89 95 91
rect 87 81 95 89
rect 87 79 91 81
rect 93 79 95 81
rect 87 71 95 79
rect 87 69 91 71
rect 93 69 95 71
rect 87 61 95 69
rect 87 59 91 61
rect 93 59 95 61
rect 87 55 95 59
<< alu1 >>
rect -2 95 102 100
rect -2 93 19 95
rect 21 93 31 95
rect 33 93 43 95
rect 45 93 55 95
rect 57 93 102 95
rect -2 91 102 93
rect -2 89 7 91
rect 9 89 67 91
rect 69 89 91 91
rect 93 89 102 91
rect -2 88 102 89
rect 8 41 12 82
rect 18 81 22 82
rect 42 81 46 82
rect 18 79 19 81
rect 21 79 43 81
rect 45 79 46 81
rect 18 78 22 79
rect 42 78 46 79
rect 66 81 70 88
rect 66 79 67 81
rect 69 79 70 81
rect 66 78 70 79
rect 78 81 82 82
rect 78 79 79 81
rect 81 79 82 81
rect 30 71 34 72
rect 78 71 82 79
rect 8 39 9 41
rect 11 39 12 41
rect 8 18 12 39
rect 19 69 31 71
rect 33 69 67 71
rect 19 22 21 69
rect 30 68 34 69
rect 28 41 32 62
rect 28 39 29 41
rect 31 39 32 41
rect 18 21 22 22
rect 18 19 19 21
rect 21 19 22 21
rect 18 18 22 19
rect 28 18 32 39
rect 38 41 42 62
rect 54 61 58 62
rect 54 59 55 61
rect 57 59 58 61
rect 54 58 58 59
rect 38 39 39 41
rect 41 39 42 41
rect 38 18 42 39
rect 55 41 57 58
rect 65 52 67 69
rect 78 69 79 71
rect 81 69 82 71
rect 78 61 82 69
rect 78 59 79 61
rect 81 59 82 61
rect 64 51 68 52
rect 64 49 65 51
rect 67 49 68 51
rect 64 48 68 49
rect 68 41 72 42
rect 55 39 69 41
rect 71 39 72 41
rect 55 22 57 39
rect 68 38 72 39
rect 54 21 58 22
rect 54 19 55 21
rect 57 19 58 21
rect 54 18 58 19
rect 66 21 70 22
rect 66 19 67 21
rect 69 19 70 21
rect 66 12 70 19
rect 78 21 82 59
rect 90 81 94 88
rect 90 79 91 81
rect 93 79 94 81
rect 90 71 94 79
rect 90 69 91 71
rect 93 69 94 71
rect 90 61 94 69
rect 90 59 91 61
rect 93 59 94 61
rect 90 58 94 59
rect 78 19 79 21
rect 81 19 82 21
rect 78 18 82 19
rect 90 21 94 22
rect 90 19 91 21
rect 93 19 94 21
rect 90 12 94 19
rect -2 11 102 12
rect -2 9 7 11
rect 9 9 43 11
rect 45 9 67 11
rect 69 9 91 11
rect 93 9 102 11
rect -2 7 102 9
rect -2 5 19 7
rect 21 5 31 7
rect 33 5 102 7
rect -2 0 102 5
<< ptie >>
rect 17 7 35 9
rect 17 5 19 7
rect 21 5 31 7
rect 33 5 35 7
rect 17 3 35 5
<< ntie >>
rect 17 95 59 97
rect 17 93 19 95
rect 21 93 31 95
rect 33 93 43 95
rect 45 93 55 95
rect 57 93 59 95
rect 17 91 59 93
<< nmos >>
rect 13 15 15 25
rect 25 15 27 25
rect 37 15 39 25
rect 61 15 63 25
rect 73 5 75 25
rect 85 5 87 25
<< pmos >>
rect 13 65 15 85
rect 25 65 27 85
rect 37 65 39 85
rect 61 55 63 75
rect 73 55 75 95
rect 85 55 87 95
<< polyct1 >>
rect 9 39 11 41
rect 65 49 67 51
rect 29 39 31 41
rect 39 39 41 41
rect 69 39 71 41
<< ndifct1 >>
rect 19 19 21 21
rect 55 19 57 21
rect 67 19 69 21
rect 7 9 9 11
rect 43 9 45 11
rect 67 9 69 11
rect 79 19 81 21
rect 91 19 93 21
rect 91 9 93 11
<< ntiect1 >>
rect 19 93 21 95
rect 31 93 33 95
rect 43 93 45 95
rect 55 93 57 95
<< ptiect1 >>
rect 19 5 21 7
rect 31 5 33 7
<< pdifct1 >>
rect 7 89 9 91
rect 67 89 69 91
rect 19 79 21 81
rect 31 69 33 71
rect 43 79 45 81
rect 67 79 69 81
rect 55 59 57 61
rect 79 79 81 81
rect 79 69 81 71
rect 79 59 81 61
rect 91 89 93 91
rect 91 79 93 81
rect 91 69 93 71
rect 91 59 93 61
<< labels >>
rlabel alu1 10 50 10 50 6 i2
rlabel polyct1 40 40 40 40 6 i0
rlabel polyct1 30 40 30 40 6 i1
rlabel alu1 50 6 50 6 6 vss
rlabel alu1 50 94 50 94 6 vdd
rlabel alu1 80 50 80 50 6 nq
<< end >>
