magic
tech scmos
timestamp 1199202897
<< ab >>
rect 0 0 32 72
<< nwell >>
rect -5 32 37 77
<< pwell >>
rect -5 -5 37 32
<< poly >>
rect 12 66 14 70
rect 19 66 21 70
rect 12 43 14 46
rect 9 41 15 43
rect 9 39 11 41
rect 13 39 15 41
rect 9 37 15 39
rect 10 25 12 37
rect 19 34 21 46
rect 19 32 25 34
rect 19 30 21 32
rect 23 30 25 32
rect 19 28 25 30
rect 20 25 22 28
rect 10 14 12 19
rect 20 14 22 19
<< ndif >>
rect 2 23 10 25
rect 2 21 4 23
rect 6 21 10 23
rect 2 19 10 21
rect 12 23 20 25
rect 12 21 15 23
rect 17 21 20 23
rect 12 19 20 21
rect 22 23 30 25
rect 22 21 26 23
rect 28 21 30 23
rect 22 19 30 21
<< pdif >>
rect 7 60 12 66
rect 5 58 12 60
rect 5 56 7 58
rect 9 56 12 58
rect 5 54 12 56
rect 7 46 12 54
rect 14 46 19 66
rect 21 64 30 66
rect 21 62 26 64
rect 28 62 30 64
rect 21 57 30 62
rect 21 55 26 57
rect 28 55 30 57
rect 21 46 30 55
<< alu1 >>
rect -2 64 34 72
rect 2 58 11 59
rect 2 56 7 58
rect 9 56 11 58
rect 2 55 11 56
rect 2 33 6 55
rect 18 46 22 51
rect 10 42 22 46
rect 10 41 14 42
rect 10 39 11 41
rect 13 39 14 41
rect 10 37 14 39
rect 26 35 30 43
rect 2 29 14 33
rect 18 32 30 35
rect 18 30 21 32
rect 23 30 30 32
rect 18 29 30 30
rect 10 24 14 29
rect 10 23 19 24
rect 10 21 15 23
rect 17 21 19 23
rect 10 20 19 21
rect -2 7 34 8
rect -2 5 5 7
rect 7 5 25 7
rect 27 5 34 7
rect -2 0 34 5
<< ptie >>
rect 3 7 29 9
rect 3 5 5 7
rect 7 5 25 7
rect 27 5 29 7
rect 3 3 29 5
<< nmos >>
rect 10 19 12 25
rect 20 19 22 25
<< pmos >>
rect 12 46 14 66
rect 19 46 21 66
<< polyct1 >>
rect 11 39 13 41
rect 21 30 23 32
<< ndifct0 >>
rect 4 21 6 23
rect 26 21 28 23
<< ndifct1 >>
rect 15 21 17 23
<< ptiect1 >>
rect 5 5 7 7
rect 25 5 27 7
<< pdifct0 >>
rect 26 62 28 64
rect 26 55 28 57
<< pdifct1 >>
rect 7 56 9 58
<< alu0 >>
rect 25 62 26 64
rect 28 62 29 64
rect 25 57 29 62
rect 25 55 26 57
rect 28 55 29 57
rect 25 53 29 55
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 8 7 21
rect 25 23 29 25
rect 25 21 26 23
rect 28 21 29 23
rect 25 8 29 21
<< labels >>
rlabel alu1 4 44 4 44 6 z
rlabel alu1 12 24 12 24 6 z
rlabel polyct1 12 40 12 40 6 b
rlabel alu1 16 4 16 4 6 vss
rlabel alu1 20 32 20 32 6 a
rlabel alu1 20 48 20 48 6 b
rlabel alu1 16 68 16 68 6 vdd
rlabel alu1 28 36 28 36 6 a
<< end >>
