magic
tech scmos
timestamp 1199202835
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 59 11 64
rect 19 59 21 64
rect 29 59 31 64
rect 39 59 41 64
rect 9 34 11 49
rect 19 44 21 49
rect 16 42 24 44
rect 16 40 18 42
rect 20 40 24 42
rect 16 38 24 40
rect 9 32 15 34
rect 9 30 11 32
rect 13 30 15 32
rect 9 28 17 30
rect 15 25 17 28
rect 22 25 24 38
rect 29 43 31 49
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 29 37 35 39
rect 29 25 31 37
rect 39 34 41 49
rect 39 32 47 34
rect 39 30 43 32
rect 45 30 47 32
rect 36 28 47 30
rect 36 25 38 28
rect 15 8 17 13
rect 22 8 24 13
rect 29 8 31 13
rect 36 8 38 13
<< ndif >>
rect 10 19 15 25
rect 8 17 15 19
rect 8 15 10 17
rect 12 15 15 17
rect 8 13 15 15
rect 17 13 22 25
rect 24 13 29 25
rect 31 13 36 25
rect 38 17 49 25
rect 38 15 44 17
rect 46 15 49 17
rect 38 13 49 15
<< pdif >>
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 49 9 55
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 49 19 52
rect 21 57 29 59
rect 21 55 24 57
rect 26 55 29 57
rect 21 49 29 55
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 49 39 52
rect 41 57 49 59
rect 41 55 45 57
rect 47 55 49 57
rect 41 49 49 55
<< alu1 >>
rect -2 67 58 72
rect -2 65 49 67
rect 51 65 58 67
rect -2 64 58 65
rect 33 54 38 59
rect 33 52 34 54
rect 36 52 38 54
rect 33 50 38 52
rect 2 46 38 50
rect 2 13 6 46
rect 10 32 14 35
rect 10 30 11 32
rect 13 30 14 32
rect 10 25 14 30
rect 25 41 38 42
rect 42 41 46 51
rect 25 39 31 41
rect 33 39 38 41
rect 25 38 38 39
rect 18 29 30 34
rect 34 29 38 38
rect 42 32 46 35
rect 42 30 43 32
rect 45 30 46 32
rect 10 21 22 25
rect 18 13 22 21
rect 26 13 30 29
rect 42 25 46 30
rect 34 21 46 25
rect 34 13 38 21
rect -2 7 58 8
rect -2 5 5 7
rect 7 5 48 7
rect 50 5 58 7
rect -2 0 58 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 45 7 53 9
rect 45 5 48 7
rect 50 5 53 7
rect 45 3 53 5
<< ntie >>
rect 47 67 53 69
rect 47 65 49 67
rect 51 65 53 67
rect 47 63 53 65
<< nmos >>
rect 15 13 17 25
rect 22 13 24 25
rect 29 13 31 25
rect 36 13 38 25
<< pmos >>
rect 9 49 11 59
rect 19 49 21 59
rect 29 49 31 59
rect 39 49 41 59
<< polyct0 >>
rect 18 40 20 42
<< polyct1 >>
rect 11 30 13 32
rect 31 39 33 41
rect 43 30 45 32
<< ndifct0 >>
rect 10 15 12 17
rect 44 15 46 17
<< ntiect1 >>
rect 49 65 51 67
<< ptiect1 >>
rect 5 5 7 7
rect 48 5 50 7
<< pdifct0 >>
rect 4 55 6 57
rect 14 52 16 54
rect 24 55 26 57
rect 45 55 47 57
<< pdifct1 >>
rect 34 52 36 54
<< alu0 >>
rect 2 57 8 64
rect 2 55 4 57
rect 6 55 8 57
rect 22 57 28 64
rect 2 54 8 55
rect 13 54 17 56
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 43 57 49 64
rect 43 55 45 57
rect 47 55 49 57
rect 43 54 49 55
rect 13 52 14 54
rect 16 52 17 54
rect 13 50 17 52
rect 16 42 22 43
rect 34 42 42 43
rect 16 40 18 42
rect 20 40 22 42
rect 16 39 22 40
rect 18 34 22 39
rect 38 41 42 42
rect 38 38 46 41
rect 6 17 14 18
rect 6 15 10 17
rect 12 15 14 17
rect 6 14 14 15
rect 42 17 48 18
rect 42 15 44 17
rect 46 15 48 17
rect 42 8 48 15
<< labels >>
rlabel alu1 4 28 4 28 6 z
rlabel alu1 20 16 20 16 6 d
rlabel alu1 12 28 12 28 6 d
rlabel alu1 20 32 20 32 6 c
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 16 36 16 6 a
rlabel alu1 28 20 28 20 6 c
rlabel alu1 36 32 36 32 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 28 44 28 6 a
rlabel alu1 44 48 44 48 6 b
<< end >>
