magic
tech scmos
timestamp 1199202145
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 26 65 48 67
rect 56 65 58 70
rect 9 54 11 59
rect 19 54 21 59
rect 26 54 28 65
rect 46 62 48 65
rect 36 54 38 59
rect 9 33 11 38
rect 19 33 21 38
rect 26 35 28 38
rect 36 35 38 38
rect 9 31 21 33
rect 9 28 11 31
rect 5 26 11 28
rect 19 26 21 31
rect 25 33 31 35
rect 25 31 27 33
rect 29 31 31 33
rect 25 29 31 31
rect 36 33 42 35
rect 36 31 38 33
rect 40 31 42 33
rect 36 29 42 31
rect 26 26 28 29
rect 36 26 38 29
rect 46 26 48 46
rect 56 43 58 46
rect 56 41 63 43
rect 56 39 59 41
rect 61 39 63 41
rect 56 37 63 39
rect 56 26 58 37
rect 5 24 7 26
rect 9 24 11 26
rect 5 22 11 24
rect 9 19 11 22
rect 19 14 21 19
rect 26 14 28 19
rect 36 14 38 19
rect 46 14 48 19
rect 9 7 11 12
rect 56 11 58 16
<< ndif >>
rect 13 19 19 26
rect 21 19 26 26
rect 28 24 36 26
rect 28 22 31 24
rect 33 22 36 24
rect 28 19 36 22
rect 38 23 46 26
rect 38 21 41 23
rect 43 21 46 23
rect 38 19 46 21
rect 48 23 56 26
rect 48 21 51 23
rect 53 21 56 23
rect 48 19 56 21
rect 2 16 9 19
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 12 17 19
rect 50 16 56 19
rect 58 24 65 26
rect 58 22 61 24
rect 63 22 65 24
rect 58 20 65 22
rect 58 16 63 20
rect 13 7 19 12
rect 13 5 15 7
rect 17 5 19 7
rect 13 3 19 5
<< pdif >>
rect 13 67 19 69
rect 13 65 15 67
rect 17 65 19 67
rect 13 61 19 65
rect 13 54 17 61
rect 50 62 56 65
rect 41 54 46 62
rect 2 52 9 54
rect 2 50 4 52
rect 6 50 9 52
rect 2 45 9 50
rect 2 43 4 45
rect 6 43 9 45
rect 2 41 9 43
rect 4 38 9 41
rect 11 38 19 54
rect 21 38 26 54
rect 28 50 36 54
rect 28 48 31 50
rect 33 48 36 50
rect 28 38 36 48
rect 38 52 46 54
rect 38 50 41 52
rect 43 50 46 52
rect 38 46 46 50
rect 48 60 56 62
rect 48 58 51 60
rect 53 58 56 60
rect 48 46 56 58
rect 58 59 63 65
rect 58 57 65 59
rect 58 55 61 57
rect 63 55 65 57
rect 58 50 65 55
rect 58 48 61 50
rect 63 48 65 50
rect 58 46 65 48
rect 38 38 43 46
<< alu1 >>
rect -2 67 74 72
rect -2 65 5 67
rect 7 65 15 67
rect 17 65 74 67
rect -2 64 74 65
rect 10 50 35 51
rect 10 48 31 50
rect 33 48 35 50
rect 10 47 35 48
rect 10 45 22 47
rect 2 27 6 35
rect 2 26 14 27
rect 2 24 7 26
rect 9 24 14 26
rect 2 21 14 24
rect 18 25 22 45
rect 26 37 38 43
rect 26 33 30 37
rect 58 41 70 43
rect 58 39 59 41
rect 61 39 70 41
rect 58 37 70 39
rect 26 31 27 33
rect 29 31 30 33
rect 26 29 30 31
rect 66 29 70 37
rect 18 24 35 25
rect 18 22 31 24
rect 33 22 35 24
rect 18 21 35 22
rect -2 7 74 8
rect -2 5 15 7
rect 17 5 27 7
rect 29 5 64 7
rect 66 5 74 7
rect -2 0 74 5
<< ptie >>
rect 25 7 68 9
rect 25 5 27 7
rect 29 5 64 7
rect 66 5 68 7
rect 25 3 68 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 19 19 21 26
rect 26 19 28 26
rect 36 19 38 26
rect 46 19 48 26
rect 9 12 11 19
rect 56 16 58 26
<< pmos >>
rect 9 38 11 54
rect 19 38 21 54
rect 26 38 28 54
rect 36 38 38 54
rect 46 46 48 62
rect 56 46 58 65
<< polyct0 >>
rect 38 31 40 33
<< polyct1 >>
rect 27 31 29 33
rect 59 39 61 41
rect 7 24 9 26
<< ndifct0 >>
rect 41 21 43 23
rect 51 21 53 23
rect 4 14 6 16
rect 61 22 63 24
<< ndifct1 >>
rect 31 22 33 24
rect 15 5 17 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 27 5 29 7
rect 64 5 66 7
<< pdifct0 >>
rect 4 50 6 52
rect 4 43 6 45
rect 41 50 43 52
rect 51 58 53 60
rect 61 55 63 57
rect 61 48 63 50
<< pdifct1 >>
rect 15 65 17 67
rect 31 48 33 50
<< alu0 >>
rect 50 60 54 64
rect 3 55 44 59
rect 50 58 51 60
rect 53 58 54 60
rect 50 56 54 58
rect 60 57 64 59
rect 3 52 7 55
rect 3 50 4 52
rect 6 50 7 52
rect 40 52 44 55
rect 3 45 7 50
rect 40 50 41 52
rect 43 50 44 52
rect 60 55 61 57
rect 63 55 64 57
rect 60 50 64 55
rect 40 48 44 50
rect 50 48 61 50
rect 63 48 64 50
rect 3 43 4 45
rect 6 43 7 45
rect 3 41 7 43
rect 50 46 64 48
rect 50 34 54 46
rect 36 33 62 34
rect 36 31 38 33
rect 40 31 62 33
rect 36 30 62 31
rect 58 25 62 30
rect 40 23 44 25
rect 40 21 41 23
rect 43 21 44 23
rect 40 17 44 21
rect 2 16 44 17
rect 2 14 4 16
rect 6 14 44 16
rect 2 13 44 14
rect 50 23 54 25
rect 50 21 51 23
rect 53 21 54 23
rect 58 24 65 25
rect 58 22 61 24
rect 63 22 65 24
rect 58 21 65 22
rect 50 8 54 21
<< labels >>
rlabel alu0 5 50 5 50 6 n1
rlabel alu0 23 15 23 15 6 n3
rlabel alu0 42 19 42 19 6 n3
rlabel alu0 42 53 42 53 6 n1
rlabel alu0 49 32 49 32 6 cn
rlabel alu0 60 27 60 27 6 cn
rlabel alu0 62 52 62 52 6 cn
rlabel alu1 4 28 4 28 6 a
rlabel alu1 12 24 12 24 6 a
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 36 20 36 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 36 40 36 40 6 b
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 68 36 68 36 6 c
rlabel polyct1 60 40 60 40 6 c
<< end >>
