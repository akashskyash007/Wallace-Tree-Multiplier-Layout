magic
tech scmos
timestamp 1199203115
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 10 70 12 74
rect 22 70 24 74
rect 29 70 31 74
rect 39 70 41 74
rect 46 70 48 74
rect 10 39 12 42
rect 22 39 24 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 29 37 41 39
rect 29 35 35 37
rect 37 35 41 37
rect 29 33 41 35
rect 46 39 48 42
rect 46 37 55 39
rect 46 35 51 37
rect 53 35 55 37
rect 46 33 55 35
rect 9 30 11 33
rect 30 30 32 33
rect 46 30 48 33
rect 20 24 22 29
rect 9 9 11 12
rect 20 9 22 12
rect 9 7 22 9
rect 30 6 32 10
rect 46 6 48 10
<< ndif >>
rect 4 23 9 30
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 12 9 17
rect 11 28 18 30
rect 11 26 14 28
rect 16 26 18 28
rect 11 24 18 26
rect 25 24 30 30
rect 11 12 20 24
rect 22 21 30 24
rect 22 19 25 21
rect 27 19 30 21
rect 22 12 30 19
rect 25 10 30 12
rect 32 14 46 30
rect 32 12 38 14
rect 40 12 46 14
rect 32 10 46 12
rect 48 23 53 30
rect 48 21 55 23
rect 48 19 51 21
rect 53 19 55 21
rect 48 17 55 19
rect 48 10 53 17
<< pdif >>
rect 5 63 10 70
rect 2 61 10 63
rect 2 59 4 61
rect 6 59 10 61
rect 2 54 10 59
rect 2 52 4 54
rect 6 52 10 54
rect 2 50 10 52
rect 5 42 10 50
rect 12 68 22 70
rect 12 66 16 68
rect 18 66 22 68
rect 12 42 22 66
rect 24 42 29 70
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 42 39 52
rect 41 42 46 70
rect 48 68 57 70
rect 48 66 52 68
rect 54 66 57 68
rect 48 61 57 66
rect 48 59 52 61
rect 54 59 57 61
rect 48 42 57 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 61 38 62
rect 2 59 4 61
rect 6 59 34 61
rect 36 59 38 61
rect 2 58 38 59
rect 2 54 6 58
rect 2 52 4 54
rect 2 29 6 52
rect 33 54 38 58
rect 17 47 23 54
rect 33 52 34 54
rect 36 52 38 54
rect 33 50 38 52
rect 10 42 23 47
rect 42 46 46 55
rect 10 37 14 42
rect 33 41 46 46
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 19 37 27 38
rect 19 35 21 37
rect 23 35 27 37
rect 19 34 27 35
rect 33 37 39 41
rect 33 35 35 37
rect 37 35 39 37
rect 33 34 39 35
rect 50 37 55 47
rect 50 35 51 37
rect 53 35 55 37
rect 23 30 27 34
rect 50 30 55 35
rect 2 28 18 29
rect 2 26 14 28
rect 16 26 18 28
rect 23 26 55 30
rect 2 25 18 26
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 12 11 30
rect 20 12 22 24
rect 30 10 32 30
rect 46 10 48 30
<< pmos >>
rect 10 42 12 70
rect 22 42 24 70
rect 29 42 31 70
rect 39 42 41 70
rect 46 42 48 70
<< polyct1 >>
rect 11 35 13 37
rect 21 35 23 37
rect 35 35 37 37
rect 51 35 53 37
<< ndifct0 >>
rect 4 19 6 21
rect 25 19 27 21
rect 38 12 40 14
rect 51 19 53 21
<< ndifct1 >>
rect 14 26 16 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 16 66 18 68
rect 52 66 54 68
rect 52 59 54 61
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
rect 34 59 36 61
rect 34 52 36 54
<< alu0 >>
rect 14 66 16 68
rect 18 66 20 68
rect 14 65 20 66
rect 50 66 52 68
rect 54 66 56 68
rect 50 61 56 66
rect 50 59 52 61
rect 54 59 56 61
rect 50 58 56 59
rect 6 50 7 58
rect 2 21 55 22
rect 2 19 4 21
rect 6 19 25 21
rect 27 19 51 21
rect 53 19 55 21
rect 2 18 55 19
rect 36 14 42 15
rect 36 12 38 14
rect 40 12 42 14
<< labels >>
rlabel alu0 28 20 28 20 6 n1
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 28 28 28 6 a1
rlabel alu1 20 48 20 48 6 b
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 28 36 28 6 a1
rlabel alu1 44 28 44 28 6 a1
rlabel alu1 36 40 36 40 6 a2
rlabel alu1 44 48 44 48 6 a2
rlabel alu1 32 74 32 74 6 vdd
rlabel polyct1 52 36 52 36 6 a1
<< end >>
