magic
tech scmos
timestamp 1199543935
<< ab >>
rect 0 0 280 100
<< nwell >>
rect -2 48 282 104
<< pwell >>
rect -2 -4 282 48
<< poly >>
rect 27 95 29 98
rect 39 95 41 98
rect 51 95 53 98
rect 59 95 61 98
rect 71 95 73 98
rect 83 95 85 98
rect 91 95 93 98
rect 195 95 197 98
rect 207 95 209 98
rect 219 95 221 98
rect 231 95 233 98
rect 243 95 245 98
rect 255 95 257 98
rect 267 95 269 98
rect 121 85 123 88
rect 147 85 149 88
rect 159 85 161 88
rect 171 85 173 88
rect 183 85 185 88
rect 15 69 17 72
rect 15 53 17 55
rect 7 51 17 53
rect 7 49 9 51
rect 11 49 17 51
rect 7 47 17 49
rect 15 37 17 47
rect 27 53 29 75
rect 39 73 41 75
rect 33 71 41 73
rect 33 69 35 71
rect 37 69 41 71
rect 33 67 41 69
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 15 26 17 29
rect 27 23 29 47
rect 39 41 41 67
rect 51 63 53 75
rect 47 61 53 63
rect 47 59 49 61
rect 51 59 53 61
rect 47 57 53 59
rect 47 51 53 53
rect 59 51 61 75
rect 71 73 73 75
rect 83 73 85 75
rect 47 49 49 51
rect 51 49 61 51
rect 47 47 53 49
rect 39 39 53 41
rect 33 31 41 33
rect 33 29 35 31
rect 37 29 41 31
rect 33 27 41 29
rect 39 23 41 27
rect 51 23 53 39
rect 59 23 61 49
rect 69 71 73 73
rect 79 71 85 73
rect 69 33 71 71
rect 79 53 81 71
rect 91 63 93 75
rect 103 69 105 72
rect 85 61 93 63
rect 85 59 87 61
rect 89 59 93 61
rect 85 57 93 59
rect 195 73 197 75
rect 195 71 203 73
rect 195 69 199 71
rect 201 69 203 71
rect 195 67 203 69
rect 75 51 81 53
rect 103 51 105 55
rect 121 53 123 65
rect 147 63 149 65
rect 159 63 161 65
rect 171 63 173 65
rect 141 61 149 63
rect 157 61 163 63
rect 75 49 77 51
rect 79 49 105 51
rect 75 47 81 49
rect 79 39 81 47
rect 65 31 71 33
rect 65 29 67 31
rect 69 29 71 31
rect 65 27 71 29
rect 75 37 81 39
rect 85 41 93 43
rect 85 39 87 41
rect 89 39 93 41
rect 85 37 93 39
rect 103 37 105 49
rect 117 51 123 53
rect 117 49 119 51
rect 121 49 123 51
rect 117 47 123 49
rect 129 51 135 53
rect 141 51 143 61
rect 157 59 159 61
rect 161 59 163 61
rect 157 57 163 59
rect 169 61 175 63
rect 169 59 171 61
rect 173 59 175 61
rect 169 57 175 59
rect 167 51 173 53
rect 183 51 185 65
rect 207 63 209 75
rect 201 61 209 63
rect 201 59 203 61
rect 205 59 209 61
rect 201 57 209 59
rect 219 51 221 75
rect 231 73 233 75
rect 225 71 233 73
rect 225 69 227 71
rect 229 69 233 71
rect 225 67 233 69
rect 243 53 245 75
rect 243 51 251 53
rect 129 49 131 51
rect 133 49 169 51
rect 171 49 233 51
rect 129 47 135 49
rect 75 23 77 37
rect 81 31 87 33
rect 81 29 83 31
rect 85 29 87 31
rect 81 27 87 29
rect 71 21 77 23
rect 71 19 73 21
rect 83 19 85 27
rect 91 19 93 37
rect 103 26 105 29
rect 121 25 123 47
rect 141 29 143 49
rect 167 47 173 49
rect 147 41 153 43
rect 177 41 185 43
rect 219 41 227 43
rect 147 39 149 41
rect 151 39 179 41
rect 181 39 223 41
rect 225 39 227 41
rect 147 37 153 39
rect 177 37 185 39
rect 157 31 163 33
rect 157 29 159 31
rect 161 29 163 31
rect 141 27 149 29
rect 157 27 163 29
rect 169 31 175 33
rect 169 29 171 31
rect 173 29 175 31
rect 169 27 175 29
rect 147 25 149 27
rect 159 25 161 27
rect 171 25 173 27
rect 183 25 185 37
rect 219 37 227 39
rect 201 31 209 33
rect 201 29 203 31
rect 205 29 209 31
rect 201 27 209 29
rect 27 8 29 11
rect 39 8 41 11
rect 51 8 53 11
rect 59 8 61 11
rect 195 21 203 23
rect 195 19 199 21
rect 201 19 203 21
rect 195 17 203 19
rect 195 15 197 17
rect 207 15 209 27
rect 219 25 221 37
rect 231 25 233 49
rect 243 49 247 51
rect 249 49 251 51
rect 243 47 251 49
rect 255 43 257 55
rect 267 43 269 55
rect 245 41 269 43
rect 245 39 247 41
rect 249 39 269 41
rect 245 37 269 39
rect 243 31 251 33
rect 243 29 247 31
rect 249 29 251 31
rect 243 27 251 29
rect 243 25 245 27
rect 255 25 257 37
rect 267 25 269 37
rect 121 12 123 15
rect 147 12 149 15
rect 159 12 161 15
rect 171 12 173 15
rect 183 12 185 15
rect 71 4 73 7
rect 83 4 85 7
rect 91 4 93 7
rect 219 12 221 15
rect 231 12 233 15
rect 243 12 245 15
rect 195 2 197 5
rect 207 2 209 5
rect 255 2 257 5
rect 267 2 269 5
<< ndif >>
rect 7 29 15 37
rect 17 33 25 37
rect 17 31 21 33
rect 23 31 25 33
rect 17 29 25 31
rect 7 21 13 29
rect 43 31 49 33
rect 43 29 45 31
rect 47 29 49 31
rect 43 23 49 29
rect 7 19 9 21
rect 11 19 13 21
rect 7 17 13 19
rect 19 21 27 23
rect 19 19 21 21
rect 23 19 27 21
rect 19 11 27 19
rect 29 11 39 23
rect 41 11 51 23
rect 53 11 59 23
rect 61 21 69 23
rect 61 19 65 21
rect 67 19 69 21
rect 95 35 103 37
rect 95 33 97 35
rect 99 33 103 35
rect 95 29 103 33
rect 105 29 117 37
rect 107 25 117 29
rect 95 21 101 23
rect 95 19 97 21
rect 99 19 101 21
rect 61 11 71 19
rect 63 7 71 11
rect 73 11 83 19
rect 73 9 77 11
rect 79 9 83 11
rect 73 7 83 9
rect 85 7 91 19
rect 93 9 101 19
rect 107 15 121 25
rect 123 21 133 25
rect 123 19 129 21
rect 131 19 133 21
rect 123 15 133 19
rect 139 21 147 25
rect 139 19 141 21
rect 143 19 147 21
rect 139 15 147 19
rect 149 15 159 25
rect 161 15 171 25
rect 173 21 183 25
rect 173 19 177 21
rect 179 19 183 21
rect 173 15 183 19
rect 185 15 193 25
rect 211 21 219 25
rect 211 19 213 21
rect 215 19 219 21
rect 211 15 219 19
rect 221 21 231 25
rect 221 19 225 21
rect 227 19 231 21
rect 221 15 231 19
rect 233 15 243 25
rect 245 21 255 25
rect 245 19 249 21
rect 251 19 255 21
rect 245 15 255 19
rect 107 11 117 15
rect 107 9 109 11
rect 111 9 117 11
rect 151 11 157 15
rect 151 9 153 11
rect 155 9 157 11
rect 93 7 97 9
rect 107 7 117 9
rect 151 7 157 9
rect 187 5 195 15
rect 197 11 207 15
rect 197 9 201 11
rect 203 9 207 11
rect 197 5 207 9
rect 209 5 217 15
rect 247 11 255 15
rect 247 9 249 11
rect 251 9 255 11
rect 247 5 255 9
rect 257 21 267 25
rect 257 19 261 21
rect 263 19 267 21
rect 257 5 267 19
rect 269 21 277 25
rect 269 19 273 21
rect 275 19 277 21
rect 269 11 277 19
rect 269 9 273 11
rect 275 9 277 11
rect 269 5 277 9
<< pdif >>
rect 7 81 13 83
rect 7 79 9 81
rect 11 79 13 81
rect 7 69 13 79
rect 19 81 27 95
rect 19 79 21 81
rect 23 79 27 81
rect 19 75 27 79
rect 29 75 39 95
rect 41 75 51 95
rect 53 75 59 95
rect 61 81 71 95
rect 61 79 65 81
rect 67 79 71 81
rect 61 75 71 79
rect 73 91 83 95
rect 73 89 77 91
rect 79 89 83 91
rect 73 75 83 89
rect 85 75 91 95
rect 93 81 101 95
rect 93 79 97 81
rect 99 79 101 81
rect 93 75 101 79
rect 107 91 117 93
rect 151 93 157 95
rect 151 91 153 93
rect 155 91 157 93
rect 107 89 109 91
rect 111 89 117 91
rect 107 85 117 89
rect 151 85 157 91
rect 187 85 195 95
rect 7 55 15 69
rect 17 61 25 69
rect 17 59 21 61
rect 23 59 25 61
rect 17 55 25 59
rect 43 71 49 75
rect 43 69 45 71
rect 47 69 49 71
rect 43 67 49 69
rect 107 69 121 85
rect 95 61 103 69
rect 95 59 97 61
rect 99 59 103 61
rect 95 55 103 59
rect 105 65 121 69
rect 123 71 133 85
rect 123 69 129 71
rect 131 69 133 71
rect 123 65 133 69
rect 139 71 147 85
rect 139 69 141 71
rect 143 69 147 71
rect 139 65 147 69
rect 149 65 159 85
rect 161 65 171 85
rect 173 71 183 85
rect 173 69 177 71
rect 179 69 183 71
rect 173 65 183 69
rect 185 75 195 85
rect 197 91 207 95
rect 197 89 201 91
rect 203 89 207 91
rect 197 75 207 89
rect 209 81 219 95
rect 209 79 213 81
rect 215 79 219 81
rect 209 75 219 79
rect 221 81 231 95
rect 221 79 225 81
rect 227 79 231 81
rect 221 75 231 79
rect 233 75 243 95
rect 245 91 255 95
rect 245 89 249 91
rect 251 89 255 91
rect 245 81 255 89
rect 245 79 249 81
rect 251 79 255 81
rect 245 75 255 79
rect 185 65 193 75
rect 105 55 117 65
rect 247 71 255 75
rect 247 69 249 71
rect 251 69 255 71
rect 247 61 255 69
rect 247 59 249 61
rect 251 59 255 61
rect 247 55 255 59
rect 257 81 267 95
rect 257 79 261 81
rect 263 79 267 81
rect 257 71 267 79
rect 257 69 261 71
rect 263 69 267 71
rect 257 61 267 69
rect 257 59 261 61
rect 263 59 267 61
rect 257 55 267 59
rect 269 91 277 95
rect 269 89 273 91
rect 275 89 277 91
rect 269 81 277 89
rect 269 79 273 81
rect 275 79 277 81
rect 269 71 277 79
rect 269 69 273 71
rect 275 69 277 71
rect 269 61 277 69
rect 269 59 273 61
rect 275 59 277 61
rect 269 55 277 59
<< alu1 >>
rect -2 95 282 100
rect -2 93 127 95
rect 129 93 141 95
rect 143 93 165 95
rect 167 93 177 95
rect 179 93 282 95
rect -2 91 153 93
rect 155 91 282 93
rect -2 89 77 91
rect 79 89 109 91
rect 111 89 201 91
rect 203 89 249 91
rect 251 89 273 91
rect 275 89 282 91
rect -2 88 282 89
rect 8 81 12 88
rect 8 79 9 81
rect 11 79 12 81
rect 8 78 12 79
rect 20 81 68 82
rect 20 79 21 81
rect 23 79 65 81
rect 67 79 68 81
rect 20 78 68 79
rect 96 81 161 82
rect 212 81 216 82
rect 96 79 97 81
rect 99 79 162 81
rect 96 78 162 79
rect 96 72 100 78
rect 8 71 38 72
rect 8 69 35 71
rect 37 69 38 71
rect 8 68 38 69
rect 44 71 111 72
rect 44 69 45 71
rect 47 69 112 71
rect 44 68 112 69
rect 8 51 12 68
rect 20 61 52 62
rect 8 49 9 51
rect 11 49 12 51
rect 8 28 12 49
rect 18 59 21 61
rect 23 59 49 61
rect 51 59 52 61
rect 18 58 52 59
rect 18 34 22 58
rect 28 51 32 52
rect 28 49 29 51
rect 31 49 32 51
rect 28 41 32 49
rect 39 51 52 52
rect 39 49 49 51
rect 51 49 52 51
rect 39 48 52 49
rect 58 42 62 68
rect 55 41 62 42
rect 54 39 62 41
rect 68 52 72 62
rect 78 61 90 62
rect 78 59 87 61
rect 89 59 90 61
rect 78 58 90 59
rect 96 61 100 62
rect 96 59 97 61
rect 99 59 102 61
rect 96 58 102 59
rect 87 52 89 58
rect 68 51 80 52
rect 68 49 77 51
rect 79 49 80 51
rect 68 48 80 49
rect 87 48 92 52
rect 54 38 61 39
rect 68 38 72 48
rect 87 42 89 48
rect 78 41 90 42
rect 78 39 87 41
rect 89 39 90 41
rect 78 38 90 39
rect 18 33 24 34
rect 18 31 21 33
rect 23 32 24 33
rect 54 32 58 38
rect 98 36 102 58
rect 96 35 102 36
rect 96 33 97 35
rect 99 33 102 35
rect 96 32 100 33
rect 23 31 38 32
rect 20 30 35 31
rect 21 29 35 30
rect 37 29 38 31
rect 21 28 38 29
rect 44 31 58 32
rect 44 29 45 31
rect 47 29 58 31
rect 66 31 100 32
rect 66 29 67 31
rect 69 29 83 31
rect 85 29 100 31
rect 44 28 57 29
rect 66 28 99 29
rect 108 22 112 68
rect 8 21 12 22
rect 8 19 9 21
rect 11 19 12 21
rect 8 12 12 19
rect 20 21 24 22
rect 64 21 68 22
rect 20 19 21 21
rect 23 19 65 21
rect 67 19 68 21
rect 20 18 24 19
rect 64 18 68 19
rect 96 21 112 22
rect 96 19 97 21
rect 99 19 112 21
rect 118 51 122 72
rect 118 49 119 51
rect 121 49 122 51
rect 96 18 111 19
rect 118 18 122 49
rect 128 71 132 72
rect 128 69 129 71
rect 131 69 132 71
rect 128 52 132 69
rect 140 71 144 72
rect 140 69 141 71
rect 143 70 151 71
rect 143 69 152 70
rect 140 68 152 69
rect 141 67 152 68
rect 128 51 134 52
rect 128 49 131 51
rect 133 49 134 51
rect 128 48 134 49
rect 128 21 132 48
rect 148 41 152 67
rect 148 39 149 41
rect 151 39 152 41
rect 148 23 152 39
rect 158 61 162 78
rect 212 79 213 81
rect 215 79 216 81
rect 212 72 216 79
rect 224 81 239 82
rect 248 81 252 88
rect 224 79 225 81
rect 227 79 240 81
rect 224 78 240 79
rect 176 71 191 72
rect 198 71 216 72
rect 226 71 230 72
rect 176 69 177 71
rect 179 69 192 71
rect 176 68 192 69
rect 198 69 199 71
rect 201 69 216 71
rect 198 68 216 69
rect 188 62 192 68
rect 158 59 159 61
rect 161 59 162 61
rect 158 31 162 59
rect 170 61 181 62
rect 188 61 206 62
rect 170 59 171 61
rect 173 59 182 61
rect 170 58 182 59
rect 158 29 159 31
rect 161 29 162 31
rect 168 51 172 52
rect 168 49 169 51
rect 171 49 172 51
rect 168 32 172 49
rect 178 41 182 58
rect 178 39 179 41
rect 181 39 182 41
rect 178 38 182 39
rect 188 59 203 61
rect 205 59 206 61
rect 188 58 206 59
rect 188 32 192 58
rect 168 31 174 32
rect 168 29 171 31
rect 173 29 174 31
rect 158 28 162 29
rect 170 28 174 29
rect 188 31 206 32
rect 188 29 203 31
rect 205 29 206 31
rect 188 28 206 29
rect 141 22 152 23
rect 188 22 192 28
rect 212 22 216 68
rect 224 69 227 71
rect 229 69 230 71
rect 224 68 230 69
rect 224 42 228 68
rect 222 41 228 42
rect 222 39 223 41
rect 225 39 228 41
rect 236 42 240 78
rect 248 79 249 81
rect 251 79 252 81
rect 248 71 252 79
rect 248 69 249 71
rect 251 69 252 71
rect 248 61 252 69
rect 248 59 249 61
rect 251 59 252 61
rect 248 58 252 59
rect 258 81 264 82
rect 258 79 261 81
rect 263 79 264 81
rect 258 78 264 79
rect 272 81 276 88
rect 272 79 273 81
rect 275 79 276 81
rect 258 72 262 78
rect 258 71 264 72
rect 258 69 261 71
rect 263 69 264 71
rect 258 68 264 69
rect 272 71 276 79
rect 272 69 273 71
rect 275 69 276 71
rect 258 62 262 68
rect 258 61 264 62
rect 258 59 261 61
rect 263 59 264 61
rect 258 58 264 59
rect 272 61 276 69
rect 272 59 273 61
rect 275 59 276 61
rect 272 58 276 59
rect 258 52 262 58
rect 246 51 263 52
rect 246 49 247 51
rect 249 49 263 51
rect 246 48 263 49
rect 236 41 250 42
rect 236 39 247 41
rect 249 39 250 41
rect 222 38 226 39
rect 236 38 250 39
rect 236 22 240 38
rect 258 32 262 48
rect 246 31 263 32
rect 246 29 247 31
rect 249 29 263 31
rect 246 28 263 29
rect 258 22 262 28
rect 128 19 129 21
rect 131 19 132 21
rect 128 18 132 19
rect 140 21 152 22
rect 140 19 141 21
rect 143 20 152 21
rect 176 21 192 22
rect 143 19 151 20
rect 176 19 177 21
rect 179 19 192 21
rect 198 21 216 22
rect 198 19 199 21
rect 201 19 213 21
rect 215 19 216 21
rect 140 18 144 19
rect 176 18 191 19
rect 198 18 216 19
rect 224 21 240 22
rect 224 19 225 21
rect 227 19 240 21
rect 248 21 252 22
rect 248 19 249 21
rect 251 19 252 21
rect 224 18 239 19
rect 248 12 252 19
rect 258 21 264 22
rect 258 19 261 21
rect 263 19 264 21
rect 258 18 264 19
rect 272 21 276 22
rect 272 19 273 21
rect 275 19 276 21
rect 272 12 276 19
rect -2 11 282 12
rect -2 9 77 11
rect 79 9 109 11
rect 111 9 153 11
rect 155 9 201 11
rect 203 9 249 11
rect 251 9 273 11
rect 275 9 282 11
rect -2 7 282 9
rect -2 5 127 7
rect 129 5 141 7
rect 143 5 165 7
rect 167 5 177 7
rect 179 5 225 7
rect 227 5 237 7
rect 239 5 282 7
rect -2 0 282 5
<< ptie >>
rect 125 7 145 9
rect 163 7 181 9
rect 125 5 127 7
rect 129 5 141 7
rect 143 5 145 7
rect 125 3 145 5
rect 163 5 165 7
rect 167 5 177 7
rect 179 5 181 7
rect 223 7 241 9
rect 223 5 225 7
rect 227 5 237 7
rect 239 5 241 7
rect 163 3 181 5
rect 223 3 241 5
<< ntie >>
rect 125 95 145 97
rect 163 95 181 97
rect 125 93 127 95
rect 129 93 141 95
rect 143 93 145 95
rect 125 91 145 93
rect 163 93 165 95
rect 167 93 177 95
rect 179 93 181 95
rect 163 91 181 93
<< nmos >>
rect 15 29 17 37
rect 27 11 29 23
rect 39 11 41 23
rect 51 11 53 23
rect 59 11 61 23
rect 103 29 105 37
rect 71 7 73 19
rect 83 7 85 19
rect 91 7 93 19
rect 121 15 123 25
rect 147 15 149 25
rect 159 15 161 25
rect 171 15 173 25
rect 183 15 185 25
rect 219 15 221 25
rect 231 15 233 25
rect 243 15 245 25
rect 195 5 197 15
rect 207 5 209 15
rect 255 5 257 25
rect 267 5 269 25
<< pmos >>
rect 27 75 29 95
rect 39 75 41 95
rect 51 75 53 95
rect 59 75 61 95
rect 71 75 73 95
rect 83 75 85 95
rect 91 75 93 95
rect 15 55 17 69
rect 103 55 105 69
rect 121 65 123 85
rect 147 65 149 85
rect 159 65 161 85
rect 171 65 173 85
rect 183 65 185 85
rect 195 75 197 95
rect 207 75 209 95
rect 219 75 221 95
rect 231 75 233 95
rect 243 75 245 95
rect 255 55 257 95
rect 267 55 269 95
<< polyct1 >>
rect 9 49 11 51
rect 35 69 37 71
rect 29 49 31 51
rect 49 59 51 61
rect 49 49 51 51
rect 35 29 37 31
rect 87 59 89 61
rect 199 69 201 71
rect 77 49 79 51
rect 67 29 69 31
rect 87 39 89 41
rect 119 49 121 51
rect 159 59 161 61
rect 171 59 173 61
rect 203 59 205 61
rect 227 69 229 71
rect 131 49 133 51
rect 169 49 171 51
rect 83 29 85 31
rect 149 39 151 41
rect 179 39 181 41
rect 223 39 225 41
rect 159 29 161 31
rect 171 29 173 31
rect 203 29 205 31
rect 199 19 201 21
rect 247 49 249 51
rect 247 39 249 41
rect 247 29 249 31
<< ndifct1 >>
rect 21 31 23 33
rect 45 29 47 31
rect 9 19 11 21
rect 21 19 23 21
rect 65 19 67 21
rect 97 33 99 35
rect 97 19 99 21
rect 77 9 79 11
rect 129 19 131 21
rect 141 19 143 21
rect 177 19 179 21
rect 213 19 215 21
rect 225 19 227 21
rect 249 19 251 21
rect 109 9 111 11
rect 153 9 155 11
rect 201 9 203 11
rect 249 9 251 11
rect 261 19 263 21
rect 273 19 275 21
rect 273 9 275 11
<< ntiect1 >>
rect 127 93 129 95
rect 141 93 143 95
rect 165 93 167 95
rect 177 93 179 95
<< ptiect1 >>
rect 127 5 129 7
rect 141 5 143 7
rect 165 5 167 7
rect 177 5 179 7
rect 225 5 227 7
rect 237 5 239 7
<< pdifct1 >>
rect 9 79 11 81
rect 21 79 23 81
rect 65 79 67 81
rect 77 89 79 91
rect 97 79 99 81
rect 153 91 155 93
rect 109 89 111 91
rect 21 59 23 61
rect 45 69 47 71
rect 97 59 99 61
rect 129 69 131 71
rect 141 69 143 71
rect 177 69 179 71
rect 201 89 203 91
rect 213 79 215 81
rect 225 79 227 81
rect 249 89 251 91
rect 249 79 251 81
rect 249 69 251 71
rect 249 59 251 61
rect 261 79 263 81
rect 261 69 263 71
rect 261 59 263 61
rect 273 89 275 91
rect 273 79 275 81
rect 273 69 275 71
rect 273 59 275 61
<< labels >>
rlabel polyct1 30 50 30 50 6 i2
rlabel polyct1 10 50 10 50 6 cmd1
rlabel alu1 80 40 80 40 6 i0
rlabel polyct1 50 50 50 50 6 i1
rlabel alu1 70 50 70 50 6 cmd0
rlabel alu1 80 60 80 60 6 i0
rlabel alu1 120 45 120 45 6 ck
rlabel alu1 90 50 90 50 6 i0
rlabel alu1 140 6 140 6 6 vss
rlabel alu1 140 94 140 94 6 vdd
rlabel alu1 260 50 260 50 6 q
<< end >>
