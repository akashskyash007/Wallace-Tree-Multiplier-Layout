magic
tech scmos
timestamp 1199202827
<< ab >>
rect 0 0 128 72
<< nwell >>
rect -5 32 133 77
<< pwell >>
rect -5 -5 133 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 40 65 42 70
rect 50 65 52 70
rect 60 65 62 70
rect 70 65 72 70
rect 97 65 99 70
rect 107 65 109 70
rect 117 65 119 70
rect 9 35 11 39
rect 19 35 21 39
rect 40 35 42 38
rect 50 35 52 38
rect 60 35 62 38
rect 70 35 72 38
rect 97 35 99 38
rect 107 35 109 38
rect 117 35 119 38
rect 2 33 11 35
rect 2 31 4 33
rect 6 31 11 33
rect 2 29 11 31
rect 9 26 11 29
rect 16 33 23 35
rect 16 31 19 33
rect 21 31 23 33
rect 33 33 45 35
rect 33 31 35 33
rect 37 31 45 33
rect 16 29 28 31
rect 16 26 18 29
rect 26 26 28 29
rect 33 29 45 31
rect 33 26 35 29
rect 43 26 45 29
rect 50 33 62 35
rect 50 31 52 33
rect 54 31 62 33
rect 50 29 62 31
rect 50 26 52 29
rect 60 26 62 29
rect 67 33 73 35
rect 67 31 69 33
rect 71 31 73 33
rect 97 33 119 35
rect 97 31 99 33
rect 101 31 107 33
rect 109 31 119 33
rect 67 29 73 31
rect 77 29 119 31
rect 67 26 69 29
rect 77 26 79 29
rect 87 26 89 29
rect 97 26 99 29
rect 107 26 109 29
rect 117 26 119 29
rect 107 11 109 16
rect 117 11 119 16
rect 9 2 11 6
rect 16 2 18 6
rect 26 2 28 6
rect 33 2 35 6
rect 43 2 45 6
rect 50 2 52 6
rect 60 2 62 6
rect 67 2 69 6
rect 77 2 79 6
rect 87 2 89 6
rect 97 2 99 6
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 6 9 13
rect 11 6 16 26
rect 18 10 26 26
rect 18 8 21 10
rect 23 8 26 10
rect 18 6 26 8
rect 28 6 33 26
rect 35 17 43 26
rect 35 15 38 17
rect 40 15 43 17
rect 35 6 43 15
rect 45 6 50 26
rect 52 10 60 26
rect 52 8 55 10
rect 57 8 60 10
rect 52 6 60 8
rect 62 6 67 26
rect 69 24 77 26
rect 69 22 72 24
rect 74 22 77 24
rect 69 17 77 22
rect 69 15 72 17
rect 74 15 77 17
rect 69 6 77 15
rect 79 24 87 26
rect 79 22 82 24
rect 84 22 87 24
rect 79 6 87 22
rect 89 17 97 26
rect 89 15 92 17
rect 94 15 97 17
rect 89 6 97 15
rect 99 24 107 26
rect 99 22 102 24
rect 104 22 107 24
rect 99 16 107 22
rect 109 20 117 26
rect 109 18 112 20
rect 114 18 117 20
rect 109 16 117 18
rect 119 24 126 26
rect 119 22 122 24
rect 124 22 126 24
rect 119 20 126 22
rect 119 16 124 20
rect 99 6 104 16
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 39 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 39 19 48
rect 21 64 28 66
rect 21 62 24 64
rect 26 62 28 64
rect 21 57 28 62
rect 21 55 24 57
rect 26 55 28 57
rect 21 39 28 55
rect 33 63 40 65
rect 33 61 35 63
rect 37 61 40 63
rect 33 56 40 61
rect 33 54 35 56
rect 37 54 40 56
rect 33 38 40 54
rect 42 56 50 65
rect 42 54 45 56
rect 47 54 50 56
rect 42 49 50 54
rect 42 47 45 49
rect 47 47 50 49
rect 42 38 50 47
rect 52 63 60 65
rect 52 61 55 63
rect 57 61 60 63
rect 52 56 60 61
rect 52 54 55 56
rect 57 54 60 56
rect 52 38 60 54
rect 62 56 70 65
rect 62 54 65 56
rect 67 54 70 56
rect 62 49 70 54
rect 62 47 65 49
rect 67 47 70 49
rect 62 38 70 47
rect 72 59 77 65
rect 92 59 97 65
rect 72 57 97 59
rect 72 55 75 57
rect 77 55 83 57
rect 85 55 92 57
rect 94 55 97 57
rect 72 38 97 55
rect 99 56 107 65
rect 99 54 102 56
rect 104 54 107 56
rect 99 49 107 54
rect 99 47 102 49
rect 104 47 107 49
rect 99 38 107 47
rect 109 63 117 65
rect 109 61 112 63
rect 114 61 117 63
rect 109 56 117 61
rect 109 54 112 56
rect 114 54 117 56
rect 109 38 117 54
rect 119 51 124 65
rect 119 49 126 51
rect 119 47 122 49
rect 124 47 126 49
rect 119 42 126 47
rect 119 40 122 42
rect 124 40 126 42
rect 119 38 126 40
<< alu1 >>
rect -2 67 130 72
rect -2 65 83 67
rect 85 65 130 67
rect -2 64 130 65
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 2 42 6 51
rect 13 50 17 55
rect 44 56 48 58
rect 44 54 45 56
rect 47 54 48 56
rect 44 50 48 54
rect 64 56 70 59
rect 64 54 65 56
rect 67 54 70 56
rect 101 56 105 58
rect 101 54 102 56
rect 104 54 105 56
rect 64 50 70 54
rect 101 50 105 54
rect 121 50 126 51
rect 13 48 14 50
rect 16 49 126 50
rect 16 48 45 49
rect 13 47 45 48
rect 47 47 65 49
rect 67 47 102 49
rect 104 47 122 49
rect 124 47 126 49
rect 13 46 126 47
rect 2 38 64 42
rect 2 33 7 38
rect 2 31 4 33
rect 6 31 7 33
rect 2 29 7 31
rect 17 33 29 34
rect 17 31 19 33
rect 21 31 29 33
rect 17 30 29 31
rect 33 33 39 38
rect 60 34 64 38
rect 33 31 35 33
rect 37 31 39 33
rect 33 30 39 31
rect 43 33 56 34
rect 43 31 52 33
rect 54 31 56 33
rect 43 30 56 31
rect 60 33 73 34
rect 60 31 69 33
rect 71 31 73 33
rect 60 30 73 31
rect 25 26 29 30
rect 43 26 47 30
rect 82 26 86 46
rect 121 42 126 46
rect 97 34 103 42
rect 121 40 122 42
rect 124 40 126 42
rect 97 33 111 34
rect 97 31 99 33
rect 101 31 107 33
rect 109 31 111 33
rect 97 30 111 31
rect 25 22 47 26
rect 80 24 106 26
rect 80 22 82 24
rect 84 22 102 24
rect 104 22 106 24
rect 121 24 126 40
rect 121 22 122 24
rect 124 22 126 24
rect 80 21 106 22
rect 121 13 126 22
rect -2 7 130 8
rect -2 5 113 7
rect 115 5 121 7
rect 123 5 130 7
rect -2 0 130 5
<< ptie >>
rect 111 7 125 9
rect 111 5 113 7
rect 115 5 121 7
rect 123 5 125 7
rect 111 3 125 5
<< ntie >>
rect 81 67 88 69
rect 81 65 83 67
rect 85 65 88 67
rect 81 63 88 65
<< nmos >>
rect 9 6 11 26
rect 16 6 18 26
rect 26 6 28 26
rect 33 6 35 26
rect 43 6 45 26
rect 50 6 52 26
rect 60 6 62 26
rect 67 6 69 26
rect 77 6 79 26
rect 87 6 89 26
rect 97 6 99 26
rect 107 16 109 26
rect 117 16 119 26
<< pmos >>
rect 9 39 11 66
rect 19 39 21 66
rect 40 38 42 65
rect 50 38 52 65
rect 60 38 62 65
rect 70 38 72 65
rect 97 38 99 65
rect 107 38 109 65
rect 117 38 119 65
<< polyct1 >>
rect 4 31 6 33
rect 19 31 21 33
rect 35 31 37 33
rect 52 31 54 33
rect 69 31 71 33
rect 99 31 101 33
rect 107 31 109 33
<< ndifct0 >>
rect 4 22 6 24
rect 4 15 6 17
rect 21 8 23 10
rect 38 15 40 17
rect 55 8 57 10
rect 72 22 74 24
rect 72 15 74 17
rect 92 15 94 17
rect 112 18 114 20
<< ndifct1 >>
rect 82 22 84 24
rect 102 22 104 24
rect 122 22 124 24
<< ntiect1 >>
rect 83 65 85 67
<< ptiect1 >>
rect 113 5 115 7
rect 121 5 123 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 24 62 26 64
rect 24 55 26 57
rect 35 61 37 63
rect 35 54 37 56
rect 55 61 57 63
rect 55 54 57 56
rect 75 55 77 57
rect 83 55 85 57
rect 92 55 94 57
rect 112 61 114 63
rect 112 54 114 56
<< pdifct1 >>
rect 14 55 16 57
rect 14 48 16 50
rect 45 54 47 56
rect 45 47 47 49
rect 65 54 67 56
rect 65 47 67 49
rect 102 54 104 56
rect 102 47 104 49
rect 122 47 124 49
rect 122 40 124 42
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 22 57 28 62
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 33 63 39 64
rect 33 61 35 63
rect 37 61 39 63
rect 33 56 39 61
rect 53 63 59 64
rect 53 61 55 63
rect 57 61 59 63
rect 33 54 35 56
rect 37 54 39 56
rect 33 53 39 54
rect 53 56 59 61
rect 53 54 55 56
rect 57 54 59 56
rect 53 53 59 54
rect 73 58 79 64
rect 90 58 96 64
rect 110 63 116 64
rect 110 61 112 63
rect 114 61 116 63
rect 73 57 96 58
rect 73 55 75 57
rect 77 55 83 57
rect 85 55 92 57
rect 94 55 96 57
rect 73 54 96 55
rect 110 56 116 61
rect 110 54 112 56
rect 114 54 116 56
rect 110 53 116 54
rect 2 24 8 25
rect 2 22 4 24
rect 6 22 8 24
rect 71 24 75 26
rect 71 22 72 24
rect 74 22 75 24
rect 2 18 8 22
rect 71 18 75 22
rect 111 20 115 22
rect 111 18 112 20
rect 114 18 115 20
rect 2 17 115 18
rect 2 15 4 17
rect 6 15 38 17
rect 40 15 72 17
rect 74 15 92 17
rect 94 15 115 17
rect 2 14 115 15
rect 19 10 25 11
rect 19 8 21 10
rect 23 8 25 10
rect 53 10 59 11
rect 53 8 55 10
rect 57 8 59 10
<< labels >>
rlabel alu0 5 19 5 19 6 n2
rlabel alu0 73 20 73 20 6 n2
rlabel alu0 58 16 58 16 6 n2
rlabel polyct1 20 32 20 32 6 a
rlabel alu1 4 40 4 40 6 b
rlabel alu1 12 40 12 40 6 b
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 44 24 44 24 6 a
rlabel alu1 36 24 36 24 6 a
rlabel alu1 28 24 28 24 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 36 36 36 6 b
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 64 4 64 4 6 vss
rlabel alu1 68 32 68 32 6 b
rlabel alu1 52 32 52 32 6 a
rlabel alu1 52 40 52 40 6 b
rlabel alu1 60 40 60 40 6 b
rlabel alu1 52 48 52 48 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 60 48 60 48 6 z
rlabel alu1 64 68 64 68 6 vdd
rlabel alu1 100 24 100 24 6 z
rlabel alu1 92 24 92 24 6 z
rlabel alu1 84 36 84 36 6 z
rlabel alu1 100 36 100 36 6 c
rlabel alu1 76 48 76 48 6 z
rlabel alu1 100 48 100 48 6 z
rlabel alu1 92 48 92 48 6 z
rlabel polyct1 108 32 108 32 6 c
rlabel alu1 124 32 124 32 6 z
rlabel alu1 108 48 108 48 6 z
rlabel alu1 116 48 116 48 6 z
<< end >>
