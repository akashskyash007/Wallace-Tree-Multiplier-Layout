magic
tech scmos
timestamp 1199202753
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 30 67 32 72
rect 37 67 39 72
rect 9 60 11 65
rect 19 60 21 65
rect 9 49 11 52
rect 9 47 15 49
rect 9 45 11 47
rect 13 45 15 47
rect 9 43 15 45
rect 9 30 11 43
rect 19 39 21 52
rect 30 49 32 52
rect 25 47 32 49
rect 25 45 27 47
rect 29 45 32 47
rect 25 43 32 45
rect 16 37 23 39
rect 16 35 19 37
rect 21 35 23 37
rect 16 33 23 35
rect 16 30 18 33
rect 27 30 29 43
rect 37 39 39 52
rect 37 37 46 39
rect 37 35 42 37
rect 44 35 46 37
rect 37 33 46 35
rect 37 30 39 33
rect 9 18 11 23
rect 16 18 18 23
rect 27 19 29 24
rect 37 19 39 24
<< ndif >>
rect 2 27 9 30
rect 2 25 4 27
rect 6 25 9 27
rect 2 23 9 25
rect 11 23 16 30
rect 18 28 27 30
rect 18 26 21 28
rect 23 26 27 28
rect 18 24 27 26
rect 29 28 37 30
rect 29 26 32 28
rect 34 26 37 28
rect 29 24 37 26
rect 39 24 46 30
rect 18 23 25 24
rect 41 13 46 24
rect 40 11 46 13
rect 40 9 42 11
rect 44 9 46 11
rect 40 7 46 9
<< pdif >>
rect 2 71 8 73
rect 2 69 4 71
rect 6 69 8 71
rect 2 67 8 69
rect 2 60 7 67
rect 23 61 30 67
rect 23 60 25 61
rect 2 52 9 60
rect 11 56 19 60
rect 11 54 14 56
rect 16 54 19 56
rect 11 52 19 54
rect 21 59 25 60
rect 27 59 30 61
rect 21 52 30 59
rect 32 52 37 67
rect 39 58 44 67
rect 39 56 46 58
rect 39 54 42 56
rect 44 54 46 56
rect 39 52 46 54
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 71 50 79
rect -2 69 4 71
rect 6 69 50 71
rect -2 68 50 69
rect 2 56 18 57
rect 2 54 14 56
rect 16 54 18 56
rect 34 55 38 63
rect 2 53 18 54
rect 2 28 6 53
rect 26 49 38 55
rect 10 47 14 49
rect 26 47 30 49
rect 10 45 11 47
rect 13 45 22 47
rect 10 41 22 45
rect 26 45 27 47
rect 29 45 30 47
rect 26 41 30 45
rect 10 33 14 41
rect 41 37 46 39
rect 41 35 42 37
rect 44 35 46 37
rect 2 27 14 28
rect 2 25 4 27
rect 6 25 14 27
rect 2 24 14 25
rect 10 17 14 24
rect 41 33 46 35
rect 42 22 46 33
rect 33 17 46 22
rect -2 11 50 12
rect -2 9 42 11
rect 44 9 50 11
rect -2 1 50 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 9 23 11 30
rect 16 23 18 30
rect 27 24 29 30
rect 37 24 39 30
<< pmos >>
rect 9 52 11 60
rect 19 52 21 60
rect 30 52 32 67
rect 37 52 39 67
<< polyct0 >>
rect 19 35 21 37
<< polyct1 >>
rect 11 45 13 47
rect 27 45 29 47
rect 42 35 44 37
<< ndifct0 >>
rect 21 26 23 28
rect 32 26 34 28
<< ndifct1 >>
rect 4 25 6 27
rect 42 9 44 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 25 59 27 61
rect 42 54 44 56
<< pdifct1 >>
rect 4 69 6 71
rect 14 54 16 56
<< alu0 >>
rect 23 61 29 68
rect 23 59 25 61
rect 27 59 29 61
rect 23 58 29 59
rect 41 56 45 58
rect 41 54 42 56
rect 44 54 45 56
rect 41 46 45 54
rect 34 42 45 46
rect 34 38 38 42
rect 17 37 38 38
rect 17 35 19 37
rect 21 35 38 37
rect 17 34 38 35
rect 20 28 24 30
rect 20 26 21 28
rect 23 26 24 28
rect 20 12 24 26
rect 30 28 36 34
rect 30 26 32 28
rect 34 26 36 28
rect 30 25 36 26
<< labels >>
rlabel alu0 33 31 33 31 6 nd
rlabel alu0 27 36 27 36 6 nd
rlabel alu0 43 50 43 50 6 nd
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 44 20 44 6 c
rlabel alu1 12 40 12 40 6 c
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 48 28 48 6 a
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 36 20 36 20 6 b
rlabel alu1 44 28 44 28 6 b
rlabel alu1 36 56 36 56 6 a
<< end >>
