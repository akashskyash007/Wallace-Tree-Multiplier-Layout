magic
tech scmos
timestamp 1199202567
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 9 35 11 42
rect 19 35 21 42
rect 29 35 31 42
rect 39 35 41 42
rect 49 36 51 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 31 35
rect 19 31 27 33
rect 29 31 31 33
rect 19 29 31 31
rect 35 33 41 35
rect 35 31 37 33
rect 39 31 41 33
rect 35 29 41 31
rect 45 34 51 36
rect 45 32 47 34
rect 49 32 51 34
rect 45 30 51 32
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 47 26 49 30
rect 47 7 49 12
rect 12 2 14 6
rect 19 2 21 6
rect 29 2 31 6
rect 36 2 38 6
<< ndif >>
rect 4 10 12 26
rect 4 8 7 10
rect 9 8 12 10
rect 4 6 12 8
rect 14 6 19 26
rect 21 17 29 26
rect 21 15 24 17
rect 26 15 29 17
rect 21 6 29 15
rect 31 6 36 26
rect 38 17 47 26
rect 38 15 41 17
rect 43 15 47 17
rect 38 12 47 15
rect 49 24 56 26
rect 49 22 52 24
rect 54 22 56 24
rect 49 17 56 22
rect 49 15 52 17
rect 54 15 56 17
rect 49 12 56 15
rect 38 10 45 12
rect 38 8 41 10
rect 43 8 45 10
rect 38 6 45 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 42 9 55
rect 11 56 19 66
rect 11 54 14 56
rect 16 54 19 56
rect 11 49 19 54
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 42 29 55
rect 31 56 39 66
rect 31 54 34 56
rect 36 54 39 56
rect 31 49 39 54
rect 31 47 34 49
rect 36 47 39 49
rect 31 42 39 47
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 57 49 62
rect 41 55 44 57
rect 46 55 49 57
rect 41 42 49 55
rect 43 39 49 42
rect 51 52 56 66
rect 51 50 58 52
rect 51 48 54 50
rect 56 48 58 50
rect 51 43 58 48
rect 51 41 54 43
rect 56 41 58 43
rect 51 39 58 41
<< alu1 >>
rect -2 64 66 72
rect 33 56 38 59
rect 33 54 34 56
rect 36 54 38 56
rect 33 50 38 54
rect 2 49 38 50
rect 2 47 14 49
rect 16 47 34 49
rect 36 47 38 49
rect 2 46 38 47
rect 2 18 6 46
rect 42 42 46 51
rect 17 34 23 42
rect 33 38 50 42
rect 46 34 50 38
rect 17 33 31 34
rect 17 31 27 33
rect 29 31 31 33
rect 17 30 31 31
rect 46 32 47 34
rect 49 32 50 34
rect 46 30 50 32
rect 2 17 31 18
rect 2 15 24 17
rect 26 15 31 17
rect 2 14 31 15
rect -2 0 66 8
<< nmos >>
rect 12 6 14 26
rect 19 6 21 26
rect 29 6 31 26
rect 36 6 38 26
rect 47 12 49 26
<< pmos >>
rect 9 42 11 66
rect 19 42 21 66
rect 29 42 31 66
rect 39 42 41 66
rect 49 39 51 66
<< polyct0 >>
rect 11 31 13 33
rect 37 31 39 33
<< polyct1 >>
rect 27 31 29 33
rect 47 32 49 34
<< ndifct0 >>
rect 7 8 9 10
rect 41 15 43 17
rect 52 22 54 24
rect 52 15 54 17
rect 41 8 43 10
<< ndifct1 >>
rect 24 15 26 17
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 54 16 56
rect 24 62 26 64
rect 24 55 26 57
rect 44 62 46 64
rect 44 55 46 57
rect 54 48 56 50
rect 54 41 56 43
<< pdifct1 >>
rect 14 47 16 49
rect 34 54 36 56
rect 34 47 36 49
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 22 62 24 64
rect 26 62 28 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 56 17 58
rect 13 54 14 56
rect 16 54 17 56
rect 22 57 28 62
rect 42 62 44 64
rect 46 62 48 64
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 42 57 48 62
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 13 50 17 54
rect 53 50 57 52
rect 53 48 54 50
rect 56 48 57 50
rect 53 43 57 48
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 35 33 41 34
rect 35 31 37 33
rect 39 31 41 33
rect 35 26 41 31
rect 53 41 54 43
rect 56 41 57 43
rect 53 26 57 41
rect 10 24 57 26
rect 10 22 52 24
rect 54 22 57 24
rect 39 17 45 18
rect 39 15 41 17
rect 43 15 45 17
rect 5 10 11 11
rect 5 8 7 10
rect 9 8 11 10
rect 39 10 45 15
rect 51 17 55 22
rect 51 15 52 17
rect 54 15 55 17
rect 51 13 55 15
rect 39 8 41 10
rect 43 8 45 10
<< labels >>
rlabel alu0 12 28 12 28 6 an
rlabel alu0 53 19 53 19 6 an
rlabel alu0 38 28 38 28 6 an
rlabel alu0 55 37 55 37 6 an
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel polyct1 28 32 28 32 6 b
rlabel alu1 20 36 20 36 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 40 36 40 6 a
rlabel alu1 44 44 44 44 6 a
rlabel alu1 36 56 36 56 6 z
rlabel alu1 32 68 32 68 6 vdd
<< end >>
