magic
tech scmos
timestamp 1199202850
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 32 69 34 74
rect 42 69 44 74
rect 64 53 70 55
rect 64 51 66 53
rect 68 51 70 53
rect 64 49 70 51
rect 54 45 60 47
rect 9 35 11 44
rect 19 41 21 44
rect 32 41 34 44
rect 19 39 25 41
rect 19 37 21 39
rect 23 37 25 39
rect 32 39 38 41
rect 32 37 34 39
rect 36 37 38 39
rect 19 35 25 37
rect 29 35 38 37
rect 42 39 44 44
rect 54 43 56 45
rect 58 43 60 45
rect 54 41 60 43
rect 42 37 49 39
rect 42 35 45 37
rect 47 35 49 37
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 17 31
rect 15 26 17 29
rect 22 26 24 35
rect 29 26 31 35
rect 42 33 49 35
rect 42 31 48 33
rect 54 32 56 41
rect 64 37 66 49
rect 36 29 48 31
rect 36 26 38 29
rect 46 26 48 29
rect 53 29 56 32
rect 60 35 66 37
rect 53 26 55 29
rect 60 26 62 35
rect 72 33 78 35
rect 72 31 74 33
rect 76 31 78 33
rect 67 29 78 31
rect 67 26 69 29
rect 15 6 17 11
rect 22 6 24 11
rect 29 6 31 11
rect 36 6 38 11
rect 46 6 48 11
rect 53 6 55 11
rect 60 6 62 11
rect 67 6 69 11
<< ndif >>
rect 6 11 15 26
rect 17 11 22 26
rect 24 11 29 26
rect 31 11 36 26
rect 38 21 46 26
rect 38 19 41 21
rect 43 19 46 21
rect 38 11 46 19
rect 48 11 53 26
rect 55 11 60 26
rect 62 11 67 26
rect 69 15 77 26
rect 69 13 72 15
rect 74 13 77 15
rect 69 11 77 13
rect 6 9 9 11
rect 11 9 13 11
rect 6 7 13 9
<< pdif >>
rect 24 69 30 71
rect 2 67 9 69
rect 2 65 4 67
rect 6 65 9 67
rect 2 60 9 65
rect 2 58 4 60
rect 6 58 9 60
rect 2 44 9 58
rect 11 61 19 69
rect 11 59 14 61
rect 16 59 19 61
rect 11 53 19 59
rect 11 51 14 53
rect 16 51 19 53
rect 11 44 19 51
rect 21 68 32 69
rect 21 66 26 68
rect 28 66 32 68
rect 21 44 32 66
rect 34 61 42 69
rect 34 59 37 61
rect 39 59 42 61
rect 34 44 42 59
rect 44 67 52 69
rect 44 65 47 67
rect 49 65 52 67
rect 44 60 52 65
rect 44 58 47 60
rect 49 58 52 60
rect 44 44 52 58
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 12 61 41 62
rect 12 59 14 61
rect 16 59 37 61
rect 39 59 41 61
rect 12 58 41 59
rect 12 54 18 58
rect 58 54 62 63
rect 2 53 18 54
rect 2 51 14 53
rect 16 51 18 53
rect 2 50 18 51
rect 24 53 71 54
rect 24 51 66 53
rect 68 51 71 53
rect 24 50 71 51
rect 2 22 6 50
rect 24 46 28 50
rect 17 42 28 46
rect 33 45 60 46
rect 33 43 56 45
rect 58 43 60 45
rect 33 42 60 43
rect 64 42 71 46
rect 20 39 24 42
rect 20 37 21 39
rect 23 37 24 39
rect 20 35 24 37
rect 33 39 39 42
rect 33 37 34 39
rect 36 37 39 39
rect 64 38 68 42
rect 10 33 14 35
rect 33 34 39 37
rect 43 37 68 38
rect 43 35 45 37
rect 47 35 68 37
rect 43 34 68 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 30 14 31
rect 72 33 78 35
rect 72 31 74 33
rect 76 31 78 33
rect 72 30 78 31
rect 10 26 78 30
rect 58 25 78 26
rect 2 21 47 22
rect 2 19 41 21
rect 43 19 47 21
rect 2 18 47 19
rect 58 17 62 25
rect -2 11 82 12
rect -2 9 9 11
rect 11 9 82 11
rect -2 1 82 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 15 11 17 26
rect 22 11 24 26
rect 29 11 31 26
rect 36 11 38 26
rect 46 11 48 26
rect 53 11 55 26
rect 60 11 62 26
rect 67 11 69 26
<< pmos >>
rect 9 44 11 69
rect 19 44 21 69
rect 32 44 34 69
rect 42 44 44 69
<< polyct1 >>
rect 66 51 68 53
rect 21 37 23 39
rect 34 37 36 39
rect 56 43 58 45
rect 45 35 47 37
rect 11 31 13 33
rect 74 31 76 33
<< ndifct0 >>
rect 72 13 74 15
<< ndifct1 >>
rect 41 19 43 21
rect 9 9 11 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 4 65 6 67
rect 4 58 6 60
rect 26 66 28 68
rect 47 65 49 67
rect 47 58 49 60
<< pdifct1 >>
rect 14 59 16 61
rect 14 51 16 53
rect 37 59 39 61
<< alu0 >>
rect 2 67 8 68
rect 2 65 4 67
rect 6 65 8 67
rect 24 66 26 68
rect 28 66 30 68
rect 24 65 30 66
rect 45 67 51 68
rect 45 65 47 67
rect 49 65 51 67
rect 2 60 8 65
rect 2 58 4 60
rect 6 58 8 60
rect 2 57 8 58
rect 45 60 51 65
rect 45 58 47 60
rect 49 58 51 60
rect 45 57 51 58
rect 71 15 75 17
rect 71 13 72 15
rect 74 13 75 15
rect 71 12 75 13
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 28 20 28 6 a
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 20 44 20 44 6 b
rlabel alu1 28 52 28 52 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 36 20 36 20 6 z
rlabel alu1 36 28 36 28 6 a
rlabel alu1 44 20 44 20 6 z
rlabel alu1 44 28 44 28 6 a
rlabel alu1 36 40 36 40 6 c
rlabel alu1 44 44 44 44 6 c
rlabel alu1 36 52 36 52 6 b
rlabel alu1 44 52 44 52 6 b
rlabel alu1 36 60 36 60 6 z
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 52 28 52 28 6 a
rlabel alu1 60 24 60 24 6 a
rlabel alu1 52 36 52 36 6 d
rlabel alu1 52 44 52 44 6 c
rlabel alu1 60 36 60 36 6 d
rlabel alu1 52 52 52 52 6 b
rlabel alu1 60 56 60 56 6 b
rlabel alu1 68 28 68 28 6 a
rlabel alu1 76 28 76 28 6 a
rlabel alu1 68 44 68 44 6 d
rlabel alu1 68 52 68 52 6 b
<< end >>
