magic
tech scmos
timestamp 1199203591
<< ab >>
rect 0 0 136 72
<< nwell >>
rect -5 32 141 77
<< pwell >>
rect -5 -5 141 32
<< poly >>
rect 20 66 22 70
rect 30 66 32 70
rect 45 66 47 70
rect 55 66 57 70
rect 85 66 87 70
rect 95 66 97 70
rect 105 66 107 70
rect 115 66 117 70
rect 125 66 127 70
rect 71 58 77 60
rect 71 56 73 58
rect 75 56 77 58
rect 65 51 67 56
rect 71 54 77 56
rect 75 51 77 54
rect 20 35 22 38
rect 30 35 32 38
rect 45 35 47 38
rect 55 35 57 38
rect 9 33 51 35
rect 9 31 11 33
rect 13 31 21 33
rect 9 29 21 31
rect 9 26 11 29
rect 19 26 21 29
rect 39 26 41 33
rect 49 26 51 33
rect 55 33 61 35
rect 55 31 57 33
rect 59 31 61 33
rect 65 33 67 38
rect 75 33 77 38
rect 85 35 87 38
rect 95 35 97 38
rect 105 35 107 38
rect 85 33 97 35
rect 101 33 107 35
rect 65 31 80 33
rect 55 29 61 31
rect 59 26 61 29
rect 66 26 68 31
rect 78 26 80 31
rect 85 31 87 33
rect 89 31 91 33
rect 85 29 91 31
rect 101 31 103 33
rect 105 31 107 33
rect 101 29 107 31
rect 115 35 117 38
rect 125 35 127 38
rect 115 33 127 35
rect 115 31 123 33
rect 125 31 127 33
rect 115 29 127 31
rect 85 26 87 29
rect 115 26 117 29
rect 125 26 127 29
rect 9 11 11 15
rect 19 4 21 9
rect 39 7 41 12
rect 49 7 51 12
rect 115 8 117 12
rect 125 8 127 12
rect 59 2 61 7
rect 66 2 68 7
rect 78 2 80 7
rect 85 2 87 7
<< ndif >>
rect 2 19 9 26
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 15 19 22
rect 14 9 19 15
rect 21 13 28 26
rect 21 11 24 13
rect 26 11 28 13
rect 32 24 39 26
rect 32 22 34 24
rect 36 22 39 24
rect 32 17 39 22
rect 32 15 34 17
rect 36 15 39 17
rect 32 12 39 15
rect 41 24 49 26
rect 41 22 44 24
rect 46 22 49 24
rect 41 12 49 22
rect 51 24 59 26
rect 51 22 54 24
rect 56 22 59 24
rect 51 17 59 22
rect 51 15 54 17
rect 56 15 59 17
rect 51 12 59 15
rect 21 9 28 11
rect 54 7 59 12
rect 61 7 66 26
rect 68 7 78 26
rect 80 7 85 26
rect 87 19 92 26
rect 87 17 94 19
rect 87 15 90 17
rect 92 15 94 17
rect 87 13 94 15
rect 87 7 92 13
rect 108 16 115 26
rect 108 14 110 16
rect 112 14 115 16
rect 108 12 115 14
rect 117 24 125 26
rect 117 22 120 24
rect 122 22 125 24
rect 117 17 125 22
rect 117 15 120 17
rect 122 15 125 17
rect 117 12 125 15
rect 127 16 134 26
rect 127 14 130 16
rect 132 14 134 16
rect 127 12 134 14
rect 70 5 72 7
rect 74 5 76 7
rect 70 3 76 5
<< pdif >>
rect 13 64 20 66
rect 13 62 15 64
rect 17 62 20 64
rect 13 57 20 62
rect 13 55 15 57
rect 17 55 20 57
rect 13 38 20 55
rect 22 49 30 66
rect 22 47 25 49
rect 27 47 30 49
rect 22 42 30 47
rect 22 40 25 42
rect 27 40 30 42
rect 22 38 30 40
rect 32 64 45 66
rect 32 62 37 64
rect 39 62 45 64
rect 32 57 45 62
rect 32 55 37 57
rect 39 55 45 57
rect 32 38 45 55
rect 47 57 55 66
rect 47 55 50 57
rect 52 55 55 57
rect 47 50 55 55
rect 47 48 50 50
rect 52 48 55 50
rect 47 38 55 48
rect 57 51 62 66
rect 80 51 85 66
rect 57 49 65 51
rect 57 47 60 49
rect 62 47 65 49
rect 57 42 65 47
rect 57 40 60 42
rect 62 40 65 42
rect 57 38 65 40
rect 67 42 75 51
rect 67 40 70 42
rect 72 40 75 42
rect 67 38 75 40
rect 77 49 85 51
rect 77 47 80 49
rect 82 47 85 49
rect 77 38 85 47
rect 87 58 95 66
rect 87 56 90 58
rect 92 56 95 58
rect 87 42 95 56
rect 87 40 90 42
rect 92 40 95 42
rect 87 38 95 40
rect 97 57 105 66
rect 97 55 100 57
rect 102 55 105 57
rect 97 50 105 55
rect 97 48 100 50
rect 102 48 105 50
rect 97 38 105 48
rect 107 49 115 66
rect 107 47 110 49
rect 112 47 115 49
rect 107 42 115 47
rect 107 40 110 42
rect 112 40 115 42
rect 107 38 115 40
rect 117 64 125 66
rect 117 62 120 64
rect 122 62 125 64
rect 117 57 125 62
rect 117 55 120 57
rect 122 55 125 57
rect 117 38 125 55
rect 127 51 132 66
rect 127 49 134 51
rect 127 47 130 49
rect 132 47 134 49
rect 127 42 134 47
rect 127 40 130 42
rect 132 40 134 42
rect 127 38 134 40
<< alu1 >>
rect -2 67 138 72
rect -2 65 5 67
rect 7 65 70 67
rect 72 65 138 67
rect -2 64 138 65
rect 98 57 103 59
rect 98 55 100 57
rect 102 55 103 57
rect 98 50 103 55
rect 58 49 100 50
rect 58 47 60 49
rect 62 47 80 49
rect 82 48 100 49
rect 102 48 103 50
rect 82 47 103 48
rect 58 46 103 47
rect 2 35 6 43
rect 58 42 63 46
rect 34 40 60 42
rect 62 40 63 42
rect 34 38 63 40
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 34 25 38 38
rect 32 24 38 25
rect 32 22 34 24
rect 36 22 38 24
rect 32 18 38 22
rect 121 33 134 35
rect 121 31 123 33
rect 125 31 134 33
rect 121 30 134 31
rect 53 24 57 26
rect 53 22 54 24
rect 56 22 57 24
rect 53 18 57 22
rect 32 17 95 18
rect 32 15 34 17
rect 36 15 54 17
rect 56 15 90 17
rect 92 15 95 17
rect 32 14 95 15
rect 130 21 134 30
rect -2 7 138 8
rect -2 5 5 7
rect 7 5 72 7
rect 74 5 100 7
rect 102 5 138 7
rect -2 0 138 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 98 7 104 24
rect 98 5 100 7
rect 102 5 104 7
rect 98 3 104 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 68 67 74 69
rect 3 40 9 65
rect 68 65 70 67
rect 72 65 74 67
rect 68 63 74 65
<< nmos >>
rect 9 15 11 26
rect 19 9 21 26
rect 39 12 41 26
rect 49 12 51 26
rect 59 7 61 26
rect 66 7 68 26
rect 78 7 80 26
rect 85 7 87 26
rect 115 12 117 26
rect 125 12 127 26
<< pmos >>
rect 20 38 22 66
rect 30 38 32 66
rect 45 38 47 66
rect 55 38 57 66
rect 65 38 67 51
rect 75 38 77 51
rect 85 38 87 66
rect 95 38 97 66
rect 105 38 107 66
rect 115 38 117 66
rect 125 38 127 66
<< polyct0 >>
rect 73 56 75 58
rect 57 31 59 33
rect 87 31 89 33
rect 103 31 105 33
<< polyct1 >>
rect 11 31 13 33
rect 123 31 125 33
<< ndifct0 >>
rect 4 17 6 19
rect 14 22 16 24
rect 24 11 26 13
rect 44 22 46 24
rect 110 14 112 16
rect 120 22 122 24
rect 120 15 122 17
rect 130 14 132 16
<< ndifct1 >>
rect 34 22 36 24
rect 34 15 36 17
rect 54 22 56 24
rect 54 15 56 17
rect 90 15 92 17
rect 72 5 74 7
<< ntiect1 >>
rect 5 65 7 67
rect 70 65 72 67
<< ptiect1 >>
rect 5 5 7 7
rect 100 5 102 7
<< pdifct0 >>
rect 15 62 17 64
rect 15 55 17 57
rect 25 47 27 49
rect 25 40 27 42
rect 37 62 39 64
rect 37 55 39 57
rect 50 55 52 57
rect 50 48 52 50
rect 70 40 72 42
rect 90 56 92 58
rect 90 40 92 42
rect 110 47 112 49
rect 110 40 112 42
rect 120 62 122 64
rect 120 55 122 57
rect 130 47 132 49
rect 130 40 132 42
<< pdifct1 >>
rect 60 47 62 49
rect 60 40 62 42
rect 80 47 82 49
rect 100 55 102 57
rect 100 48 102 50
<< alu0 >>
rect 14 62 15 64
rect 17 62 18 64
rect 14 57 18 62
rect 14 55 15 57
rect 17 55 18 57
rect 14 53 18 55
rect 35 62 37 64
rect 39 62 41 64
rect 35 57 41 62
rect 119 62 120 64
rect 122 62 123 64
rect 35 55 37 57
rect 39 55 41 57
rect 35 54 41 55
rect 49 58 94 59
rect 49 57 73 58
rect 49 55 50 57
rect 52 56 73 57
rect 75 56 90 58
rect 92 56 94 58
rect 52 55 94 56
rect 49 50 53 55
rect 119 57 123 62
rect 119 55 120 57
rect 122 55 123 57
rect 119 53 123 55
rect 23 49 50 50
rect 23 47 25 49
rect 27 48 50 49
rect 52 48 53 50
rect 27 47 53 48
rect 23 46 53 47
rect 108 49 113 51
rect 108 47 110 49
rect 112 47 113 49
rect 23 42 28 46
rect 108 43 113 47
rect 129 49 134 51
rect 129 47 130 49
rect 132 47 134 49
rect 129 43 134 47
rect 23 40 25 42
rect 27 40 28 42
rect 23 38 28 40
rect 68 42 74 43
rect 68 40 70 42
rect 72 40 74 42
rect 23 25 27 38
rect 68 34 74 40
rect 88 42 94 43
rect 108 42 134 43
rect 88 40 90 42
rect 92 40 103 42
rect 88 38 103 40
rect 108 40 110 42
rect 112 40 130 42
rect 132 40 134 42
rect 108 39 134 40
rect 99 34 103 38
rect 12 24 27 25
rect 12 22 14 24
rect 16 22 27 24
rect 12 21 27 22
rect 3 19 7 21
rect 3 17 4 19
rect 6 17 7 19
rect 3 8 7 17
rect 42 33 93 34
rect 42 31 57 33
rect 59 31 87 33
rect 89 31 93 33
rect 42 30 93 31
rect 99 33 107 34
rect 99 31 103 33
rect 105 31 107 33
rect 99 30 107 31
rect 42 24 48 30
rect 89 26 93 30
rect 112 26 116 39
rect 42 22 44 24
rect 46 22 48 24
rect 42 21 48 22
rect 89 24 123 26
rect 89 22 120 24
rect 122 22 123 24
rect 23 13 27 15
rect 109 16 113 18
rect 109 14 110 16
rect 112 14 113 16
rect 23 11 24 13
rect 26 11 27 13
rect 23 8 27 11
rect 109 8 113 14
rect 119 17 123 22
rect 119 15 120 17
rect 122 15 123 17
rect 119 13 123 15
rect 128 16 134 17
rect 128 14 130 16
rect 132 14 134 16
rect 128 8 134 14
<< labels >>
rlabel alu0 19 23 19 23 6 bn
rlabel alu0 25 35 25 35 6 bn
rlabel alu0 45 27 45 27 6 an
rlabel alu0 51 52 51 52 6 bn
rlabel alu0 67 32 67 32 6 an
rlabel alu0 91 40 91 40 6 bn
rlabel alu0 71 36 71 36 6 an
rlabel alu0 71 57 71 57 6 bn
rlabel alu0 121 19 121 19 6 an
rlabel alu0 101 36 101 36 6 bn
rlabel alu0 131 45 131 45 6 an
rlabel alu0 110 45 110 45 6 an
rlabel alu0 121 41 121 41 6 an
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 4 36 4 36 6 b
rlabel alu1 44 16 44 16 6 z
rlabel alu1 60 16 60 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 36 24 36 24 6 z
rlabel alu1 44 40 44 40 6 z
rlabel alu1 52 40 52 40 6 z
rlabel alu1 60 40 60 40 6 z
rlabel alu1 68 4 68 4 6 vss
rlabel alu1 76 16 76 16 6 z
rlabel alu1 92 16 92 16 6 z
rlabel alu1 84 16 84 16 6 z
rlabel alu1 68 16 68 16 6 z
rlabel alu1 68 48 68 48 6 z
rlabel alu1 100 52 100 52 6 z
rlabel alu1 92 48 92 48 6 z
rlabel alu1 84 48 84 48 6 z
rlabel alu1 76 48 76 48 6 z
rlabel alu1 68 68 68 68 6 vdd
rlabel polyct1 124 32 124 32 6 a
rlabel alu1 132 28 132 28 6 a
<< end >>
