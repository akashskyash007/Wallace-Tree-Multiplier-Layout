magic
tech scmos
timestamp 1199541616
<< ab >>
rect 0 0 70 100
<< nwell >>
rect -2 48 72 104
<< pwell >>
rect -2 -4 72 48
<< poly >>
rect 57 95 59 98
rect 11 85 13 88
rect 23 85 25 88
rect 35 85 37 88
rect 47 85 49 88
rect 11 53 13 65
rect 23 63 25 65
rect 35 63 37 65
rect 47 63 49 65
rect 19 61 25 63
rect 31 61 37 63
rect 41 61 49 63
rect 19 53 21 61
rect 31 53 33 61
rect 7 51 13 53
rect 7 49 9 51
rect 11 49 13 51
rect 7 47 13 49
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 11 35 13 47
rect 19 35 21 47
rect 27 35 29 47
rect 41 43 43 61
rect 57 53 59 55
rect 47 51 59 53
rect 47 49 49 51
rect 51 49 59 51
rect 47 47 59 49
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 35 37 43 39
rect 35 35 37 37
rect 57 25 59 47
rect 11 12 13 15
rect 19 12 21 15
rect 27 12 29 15
rect 35 12 37 15
rect 57 2 59 5
<< ndif >>
rect 3 15 11 35
rect 13 15 19 35
rect 21 15 27 35
rect 29 15 35 35
rect 37 23 43 35
rect 37 21 45 23
rect 37 19 41 21
rect 43 19 45 21
rect 37 17 45 19
rect 37 15 43 17
rect 3 11 9 15
rect 51 11 57 25
rect 3 9 5 11
rect 7 9 9 11
rect 49 9 57 11
rect 3 7 9 9
rect 49 7 51 9
rect 53 7 57 9
rect 49 5 57 7
rect 59 21 67 25
rect 59 19 63 21
rect 65 19 67 21
rect 59 5 67 19
<< pdif >>
rect 49 95 55 97
rect 49 93 51 95
rect 53 93 57 95
rect 3 91 9 93
rect 3 89 5 91
rect 7 89 9 91
rect 3 85 9 89
rect 27 91 33 93
rect 49 91 57 93
rect 27 89 29 91
rect 31 89 33 91
rect 27 85 33 89
rect 51 85 57 91
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 65 11 79
rect 13 81 23 85
rect 13 79 17 81
rect 19 79 23 81
rect 13 65 23 79
rect 25 65 35 85
rect 37 81 47 85
rect 37 79 41 81
rect 43 79 47 81
rect 37 65 47 79
rect 49 65 57 85
rect 51 55 57 65
rect 59 81 67 95
rect 59 79 63 81
rect 65 79 67 81
rect 59 71 67 79
rect 59 69 63 71
rect 65 69 67 71
rect 59 61 67 69
rect 59 59 63 61
rect 65 59 67 61
rect 59 55 67 59
<< alu1 >>
rect -2 95 72 100
rect -2 93 51 95
rect 53 93 72 95
rect -2 91 72 93
rect -2 89 5 91
rect 7 89 29 91
rect 31 89 72 91
rect -2 88 72 89
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 78 8 79
rect 16 81 20 82
rect 40 81 44 82
rect 58 81 66 82
rect 16 79 17 81
rect 19 79 41 81
rect 43 79 52 81
rect 16 78 20 79
rect 40 78 44 79
rect 8 51 12 72
rect 8 49 9 51
rect 11 49 12 51
rect 8 18 12 49
rect 18 51 22 72
rect 18 49 19 51
rect 21 49 22 51
rect 18 18 22 49
rect 28 51 32 72
rect 28 49 29 51
rect 31 49 32 51
rect 28 18 32 49
rect 38 41 42 72
rect 50 52 52 79
rect 48 51 52 52
rect 48 49 49 51
rect 51 49 52 51
rect 48 48 52 49
rect 38 39 39 41
rect 41 39 42 41
rect 38 28 42 39
rect 40 21 44 22
rect 50 21 52 48
rect 40 19 41 21
rect 43 19 52 21
rect 58 79 63 81
rect 65 79 66 81
rect 58 78 66 79
rect 58 72 62 78
rect 58 71 66 72
rect 58 69 63 71
rect 65 69 66 71
rect 58 68 66 69
rect 58 62 62 68
rect 58 61 66 62
rect 58 59 63 61
rect 65 59 66 61
rect 58 58 66 59
rect 58 22 62 58
rect 58 21 66 22
rect 58 19 63 21
rect 65 19 66 21
rect 40 18 44 19
rect 58 18 66 19
rect -2 11 72 12
rect -2 9 5 11
rect 7 9 72 11
rect -2 7 51 9
rect 53 7 72 9
rect -2 5 19 7
rect 21 5 35 7
rect 37 5 72 7
rect -2 0 72 5
<< ptie >>
rect 17 7 39 9
rect 17 5 19 7
rect 21 5 35 7
rect 37 5 39 7
rect 17 3 39 5
<< nmos >>
rect 11 15 13 35
rect 19 15 21 35
rect 27 15 29 35
rect 35 15 37 35
rect 57 5 59 25
<< pmos >>
rect 11 65 13 85
rect 23 65 25 85
rect 35 65 37 85
rect 47 65 49 85
rect 57 55 59 95
<< polyct1 >>
rect 9 49 11 51
rect 19 49 21 51
rect 29 49 31 51
rect 49 49 51 51
rect 39 39 41 41
<< ndifct1 >>
rect 41 19 43 21
rect 5 9 7 11
rect 51 7 53 9
rect 63 19 65 21
<< ptiect1 >>
rect 19 5 21 7
rect 35 5 37 7
<< pdifct1 >>
rect 51 93 53 95
rect 5 89 7 91
rect 29 89 31 91
rect 5 79 7 81
rect 17 79 19 81
rect 41 79 43 81
rect 63 79 65 81
rect 63 69 65 71
rect 63 59 65 61
<< labels >>
rlabel alu1 10 45 10 45 6 i0
rlabel alu1 20 45 20 45 6 i1
rlabel alu1 30 45 30 45 6 i2
rlabel alu1 35 6 35 6 6 vss
rlabel alu1 40 50 40 50 6 i3
rlabel alu1 35 94 35 94 6 vdd
rlabel alu1 60 50 60 50 6 q
<< end >>
