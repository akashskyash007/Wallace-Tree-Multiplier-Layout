magic
tech scmos
timestamp 1199202814
<< ab >>
rect 0 0 112 72
<< nwell >>
rect -5 32 117 77
<< pwell >>
rect -5 -5 117 32
<< poly >>
rect 10 58 12 63
rect 20 58 22 63
rect 30 58 32 63
rect 40 58 42 63
rect 50 58 52 63
rect 60 58 62 63
rect 70 58 72 63
rect 80 58 82 63
rect 90 58 92 63
rect 10 35 12 38
rect 20 35 22 38
rect 30 35 32 38
rect 10 33 32 35
rect 10 31 12 33
rect 14 31 19 33
rect 21 31 32 33
rect 10 29 32 31
rect 10 26 12 29
rect 20 26 22 29
rect 30 26 32 29
rect 40 35 42 38
rect 50 35 52 38
rect 60 35 62 38
rect 40 33 62 35
rect 40 31 43 33
rect 45 31 51 33
rect 53 31 62 33
rect 40 29 62 31
rect 40 26 42 29
rect 50 26 52 29
rect 60 26 62 29
rect 70 35 72 38
rect 80 35 82 38
rect 90 35 92 38
rect 70 33 103 35
rect 70 31 99 33
rect 101 31 103 33
rect 70 29 103 31
rect 70 26 72 29
rect 80 26 82 29
rect 90 26 92 29
rect 101 26 103 29
rect 90 11 92 16
rect 101 11 103 16
rect 10 2 12 6
rect 20 2 22 6
rect 30 2 32 6
rect 40 2 42 6
rect 50 2 52 6
rect 60 2 62 6
rect 70 2 72 6
rect 80 2 82 6
<< ndif >>
rect 2 17 10 26
rect 2 15 4 17
rect 6 15 10 17
rect 2 10 10 15
rect 2 8 4 10
rect 6 8 10 10
rect 2 6 10 8
rect 12 24 20 26
rect 12 22 15 24
rect 17 22 20 24
rect 12 17 20 22
rect 12 15 15 17
rect 17 15 20 17
rect 12 6 20 15
rect 22 10 30 26
rect 22 8 25 10
rect 27 8 30 10
rect 22 6 30 8
rect 32 17 40 26
rect 32 15 35 17
rect 37 15 40 17
rect 32 6 40 15
rect 42 24 50 26
rect 42 22 45 24
rect 47 22 50 24
rect 42 6 50 22
rect 52 17 60 26
rect 52 15 55 17
rect 57 15 60 17
rect 52 6 60 15
rect 62 24 70 26
rect 62 22 65 24
rect 67 22 70 24
rect 62 17 70 22
rect 62 15 65 17
rect 67 15 70 17
rect 62 6 70 15
rect 72 24 80 26
rect 72 22 75 24
rect 77 22 80 24
rect 72 6 80 22
rect 82 20 90 26
rect 82 18 85 20
rect 87 18 90 20
rect 82 16 90 18
rect 92 24 101 26
rect 92 22 95 24
rect 97 22 101 24
rect 92 16 101 22
rect 103 22 108 26
rect 103 20 110 22
rect 103 18 106 20
rect 108 18 110 20
rect 103 16 110 18
rect 82 6 87 16
<< pdif >>
rect 2 56 10 58
rect 2 54 4 56
rect 6 54 10 56
rect 2 49 10 54
rect 2 47 4 49
rect 6 47 10 49
rect 2 38 10 47
rect 12 49 20 58
rect 12 47 15 49
rect 17 47 20 49
rect 12 42 20 47
rect 12 40 15 42
rect 17 40 20 42
rect 12 38 20 40
rect 22 56 30 58
rect 22 54 25 56
rect 27 54 30 56
rect 22 49 30 54
rect 22 47 25 49
rect 27 47 30 49
rect 22 38 30 47
rect 32 49 40 58
rect 32 47 35 49
rect 37 47 40 49
rect 32 42 40 47
rect 32 40 35 42
rect 37 40 40 42
rect 32 38 40 40
rect 42 56 50 58
rect 42 54 45 56
rect 47 54 50 56
rect 42 49 50 54
rect 42 47 45 49
rect 47 47 50 49
rect 42 38 50 47
rect 52 49 60 58
rect 52 47 55 49
rect 57 47 60 49
rect 52 42 60 47
rect 52 40 55 42
rect 57 40 60 42
rect 52 38 60 40
rect 62 56 70 58
rect 62 54 65 56
rect 67 54 70 56
rect 62 49 70 54
rect 62 47 65 49
rect 67 47 70 49
rect 62 38 70 47
rect 72 49 80 58
rect 72 47 75 49
rect 77 47 80 49
rect 72 42 80 47
rect 72 40 75 42
rect 77 40 80 42
rect 72 38 80 40
rect 82 56 90 58
rect 82 54 85 56
rect 87 54 90 56
rect 82 49 90 54
rect 82 47 85 49
rect 87 47 90 49
rect 82 38 90 47
rect 92 51 97 58
rect 92 49 99 51
rect 92 47 95 49
rect 97 47 99 49
rect 92 42 99 47
rect 92 40 95 42
rect 97 40 99 42
rect 92 38 99 40
<< alu1 >>
rect -2 67 114 72
rect -2 65 105 67
rect 107 65 114 67
rect -2 64 114 65
rect 14 49 18 51
rect 14 47 15 49
rect 17 47 18 49
rect 2 34 6 43
rect 14 42 18 47
rect 34 49 38 51
rect 34 47 35 49
rect 37 47 38 49
rect 34 42 38 47
rect 54 49 58 51
rect 54 47 55 49
rect 57 47 58 49
rect 54 42 58 47
rect 74 49 78 59
rect 74 47 75 49
rect 77 47 78 49
rect 74 42 78 47
rect 90 42 96 43
rect 14 40 15 42
rect 17 40 35 42
rect 37 40 55 42
rect 57 40 75 42
rect 77 40 95 42
rect 14 39 96 40
rect 14 38 94 39
rect 74 37 94 38
rect 2 33 23 34
rect 2 31 12 33
rect 14 31 19 33
rect 21 31 23 33
rect 2 30 23 31
rect 33 33 55 34
rect 33 31 43 33
rect 45 31 51 33
rect 53 31 55 33
rect 33 30 55 31
rect 2 21 6 30
rect 33 22 39 30
rect 74 24 78 37
rect 74 22 75 24
rect 77 22 78 24
rect 106 35 110 51
rect 98 33 110 35
rect 98 31 99 33
rect 101 31 110 33
rect 98 29 110 31
rect 74 20 78 22
rect -2 7 114 8
rect -2 5 97 7
rect 99 5 105 7
rect 107 5 114 7
rect -2 0 114 5
<< ptie >>
rect 95 7 109 9
rect 95 5 97 7
rect 99 5 105 7
rect 107 5 109 7
rect 95 3 109 5
<< ntie >>
rect 103 67 109 69
rect 103 65 105 67
rect 107 65 109 67
rect 103 63 109 65
<< nmos >>
rect 10 6 12 26
rect 20 6 22 26
rect 30 6 32 26
rect 40 6 42 26
rect 50 6 52 26
rect 60 6 62 26
rect 70 6 72 26
rect 80 6 82 26
rect 90 16 92 26
rect 101 16 103 26
<< pmos >>
rect 10 38 12 58
rect 20 38 22 58
rect 30 38 32 58
rect 40 38 42 58
rect 50 38 52 58
rect 60 38 62 58
rect 70 38 72 58
rect 80 38 82 58
rect 90 38 92 58
<< polyct1 >>
rect 12 31 14 33
rect 19 31 21 33
rect 43 31 45 33
rect 51 31 53 33
rect 99 31 101 33
<< ndifct0 >>
rect 4 15 6 17
rect 4 8 6 10
rect 15 22 17 24
rect 15 15 17 17
rect 25 8 27 10
rect 35 15 37 17
rect 45 22 47 24
rect 55 15 57 17
rect 65 22 67 24
rect 65 15 67 17
rect 85 18 87 20
rect 95 22 97 24
rect 106 18 108 20
<< ndifct1 >>
rect 75 22 77 24
<< ntiect1 >>
rect 105 65 107 67
<< ptiect1 >>
rect 97 5 99 7
rect 105 5 107 7
<< pdifct0 >>
rect 4 54 6 56
rect 4 47 6 49
rect 25 54 27 56
rect 25 47 27 49
rect 45 54 47 56
rect 45 47 47 49
rect 65 54 67 56
rect 65 47 67 49
rect 85 54 87 56
rect 85 47 87 49
rect 95 47 97 49
rect 96 40 97 42
<< pdifct1 >>
rect 15 47 17 49
rect 15 40 17 42
rect 35 47 37 49
rect 35 40 37 42
rect 55 47 57 49
rect 55 40 57 42
rect 75 47 77 49
rect 75 40 77 42
rect 95 40 96 42
<< alu0 >>
rect 2 56 8 64
rect 2 54 4 56
rect 6 54 8 56
rect 2 49 8 54
rect 23 56 29 64
rect 23 54 25 56
rect 27 54 29 56
rect 2 47 4 49
rect 6 47 8 49
rect 2 46 8 47
rect 23 49 29 54
rect 43 56 49 64
rect 43 54 45 56
rect 47 54 49 56
rect 23 47 25 49
rect 27 47 29 49
rect 23 46 29 47
rect 43 49 49 54
rect 63 56 69 64
rect 63 54 65 56
rect 67 54 69 56
rect 43 47 45 49
rect 47 47 49 49
rect 43 46 49 47
rect 63 49 69 54
rect 63 47 65 49
rect 67 47 69 49
rect 63 46 69 47
rect 83 56 89 64
rect 83 54 85 56
rect 87 54 89 56
rect 83 49 89 54
rect 83 47 85 49
rect 87 47 89 49
rect 83 46 89 47
rect 94 49 98 51
rect 94 47 95 49
rect 97 47 98 49
rect 94 43 98 47
rect 96 42 98 43
rect 97 40 98 42
rect 96 39 98 40
rect 94 38 98 39
rect 94 37 95 38
rect 13 24 18 26
rect 13 22 15 24
rect 17 22 18 24
rect 43 24 69 25
rect 43 22 45 24
rect 47 22 65 24
rect 67 22 69 24
rect 13 18 18 22
rect 43 21 69 22
rect 2 17 8 18
rect 2 15 4 17
rect 6 15 8 17
rect 2 10 8 15
rect 13 17 59 18
rect 13 15 15 17
rect 17 15 35 17
rect 37 15 55 17
rect 57 15 59 17
rect 13 14 59 15
rect 64 17 69 21
rect 91 25 95 37
rect 91 24 99 25
rect 91 22 95 24
rect 97 22 99 24
rect 84 20 88 22
rect 91 21 99 22
rect 84 18 85 20
rect 87 18 88 20
rect 84 17 88 18
rect 105 20 109 22
rect 105 18 106 20
rect 108 18 109 20
rect 105 17 109 18
rect 64 15 65 17
rect 67 15 109 17
rect 64 13 109 15
rect 2 8 4 10
rect 6 8 8 10
rect 23 10 29 11
rect 23 8 25 10
rect 27 8 29 10
<< labels >>
rlabel alu0 15 20 15 20 6 n1
rlabel ndifct0 36 16 36 16 6 n1
rlabel alu0 66 19 66 19 6 n2
rlabel alu0 56 23 56 23 6 n2
rlabel alu0 107 17 107 17 6 n2
rlabel alu0 86 17 86 17 6 n2
rlabel polyct1 20 32 20 32 6 a
rlabel alu1 12 32 12 32 6 a
rlabel alu1 4 32 4 32 6 a
rlabel alu1 20 40 20 40 6 z
rlabel polyct1 44 32 44 32 6 b
rlabel polyct1 52 32 52 32 6 b
rlabel alu1 36 28 36 28 6 b
rlabel alu1 44 40 44 40 6 z
rlabel alu1 52 40 52 40 6 z
rlabel alu1 28 40 28 40 6 z
rlabel alu1 36 44 36 44 6 z
rlabel alu1 56 4 56 4 6 vss
rlabel alu1 68 40 68 40 6 z
rlabel alu1 76 40 76 40 6 z
rlabel alu1 60 40 60 40 6 z
rlabel alu1 56 68 56 68 6 vdd
rlabel polyct1 100 32 100 32 6 c
rlabel alu1 92 40 92 40 6 z
rlabel alu1 108 40 108 40 6 c
rlabel alu1 84 40 84 40 6 z
<< end >>
