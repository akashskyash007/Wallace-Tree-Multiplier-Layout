magic
tech scmos
timestamp 1199202409
<< ab >>
rect 0 0 24 72
<< nwell >>
rect -5 32 29 77
<< pwell >>
rect -5 -5 29 32
<< poly >>
rect 9 57 11 61
rect 9 35 11 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 9 24 11 29
rect 9 11 11 15
<< ndif >>
rect 2 22 9 24
rect 2 20 4 22
rect 6 20 9 22
rect 2 18 9 20
rect 4 15 9 18
rect 11 15 20 24
rect 13 7 20 15
rect 13 5 15 7
rect 17 5 20 7
rect 13 3 20 5
<< pdif >>
rect 13 67 20 69
rect 13 65 15 67
rect 17 65 20 67
rect 13 57 20 65
rect 4 52 9 57
rect 2 50 9 52
rect 2 48 4 50
rect 6 48 9 50
rect 2 43 9 48
rect 2 41 4 43
rect 6 41 9 43
rect 2 39 9 41
rect 11 39 20 57
<< alu1 >>
rect -2 67 26 72
rect -2 65 5 67
rect 7 65 15 67
rect 17 65 26 67
rect -2 64 26 65
rect 2 53 14 59
rect 2 50 6 53
rect 2 48 4 50
rect 2 43 6 48
rect 2 41 4 43
rect 2 22 6 41
rect 18 35 22 59
rect 10 33 22 35
rect 10 31 11 33
rect 13 31 22 33
rect 10 29 22 31
rect 2 20 4 22
rect 2 19 6 20
rect 2 13 14 19
rect 18 13 22 29
rect -2 7 26 8
rect -2 5 5 7
rect 7 5 15 7
rect 17 5 26 7
rect -2 0 26 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 15 11 24
<< pmos >>
rect 9 39 11 57
<< polyct1 >>
rect 11 31 13 33
<< ndifct1 >>
rect 4 20 6 22
rect 15 5 17 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct1 >>
rect 15 65 17 67
rect 4 48 6 50
rect 4 41 6 43
<< alu0 >>
rect 6 39 7 53
rect 6 19 7 24
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 4 12 4 6 vss
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 a
rlabel alu1 12 56 12 56 6 z
rlabel alu1 12 68 12 68 6 vdd
rlabel alu1 20 36 20 36 6 a
<< end >>
