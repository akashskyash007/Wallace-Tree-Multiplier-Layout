magic
tech scmos
timestamp 1199544199
<< ab >>
rect 0 0 120 100
<< nwell >>
rect -2 48 122 104
<< pwell >>
rect -2 -4 122 48
<< poly >>
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 59 95 61 98
rect 95 95 97 98
rect 107 95 109 98
rect 11 75 13 78
rect 71 75 73 78
rect 11 53 13 55
rect 23 53 25 55
rect 11 51 25 53
rect 35 53 37 55
rect 35 51 43 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 3 41 9 43
rect 47 41 49 55
rect 59 43 61 55
rect 71 53 73 55
rect 67 51 73 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 95 43 97 55
rect 107 43 109 55
rect 3 39 5 41
rect 7 39 49 41
rect 3 37 9 39
rect 17 31 23 33
rect 17 29 19 31
rect 21 29 23 31
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 11 27 25 29
rect 11 25 13 27
rect 23 25 25 27
rect 35 27 43 29
rect 35 25 37 27
rect 47 25 49 39
rect 57 41 63 43
rect 77 41 83 43
rect 57 39 59 41
rect 61 39 79 41
rect 81 39 83 41
rect 57 37 63 39
rect 77 37 83 39
rect 87 41 109 43
rect 87 39 89 41
rect 91 39 109 41
rect 87 37 109 39
rect 67 31 73 33
rect 67 29 69 31
rect 71 29 73 31
rect 59 27 73 29
rect 59 25 61 27
rect 71 25 73 27
rect 95 25 97 37
rect 107 25 109 37
rect 11 12 13 15
rect 71 12 73 15
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
rect 59 2 61 5
rect 95 2 97 5
rect 107 2 109 5
<< ndif >>
rect 75 31 83 33
rect 75 29 79 31
rect 81 29 83 31
rect 75 27 83 29
rect 75 25 81 27
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 15 11 23 15
rect 15 9 17 11
rect 19 9 23 11
rect 15 5 23 9
rect 25 5 35 25
rect 37 21 47 25
rect 37 19 41 21
rect 43 19 47 21
rect 37 5 47 19
rect 49 5 59 25
rect 61 15 71 25
rect 73 15 81 25
rect 91 21 95 25
rect 61 11 69 15
rect 61 9 65 11
rect 67 9 69 11
rect 61 5 69 9
rect 87 11 95 21
rect 87 9 89 11
rect 91 9 95 11
rect 87 5 95 9
rect 97 21 107 25
rect 97 19 101 21
rect 103 19 107 21
rect 97 5 107 19
rect 109 21 117 25
rect 109 19 113 21
rect 115 19 117 21
rect 109 11 117 19
rect 109 9 113 11
rect 115 9 117 11
rect 109 5 117 9
<< pdif >>
rect 15 91 23 95
rect 15 89 17 91
rect 19 89 23 91
rect 15 75 23 89
rect 3 71 11 75
rect 3 69 5 71
rect 7 69 11 71
rect 3 61 11 69
rect 3 59 5 61
rect 7 59 11 61
rect 3 55 11 59
rect 13 55 23 75
rect 25 81 35 95
rect 25 79 29 81
rect 31 79 35 81
rect 25 71 35 79
rect 25 69 29 71
rect 31 69 35 71
rect 25 55 35 69
rect 37 71 47 95
rect 37 69 41 71
rect 43 69 47 71
rect 37 55 47 69
rect 49 81 59 95
rect 49 79 53 81
rect 55 79 59 81
rect 49 71 59 79
rect 49 69 53 71
rect 55 69 59 71
rect 49 61 59 69
rect 49 59 53 61
rect 55 59 59 61
rect 49 55 59 59
rect 61 91 69 95
rect 61 89 65 91
rect 67 89 69 91
rect 61 75 69 89
rect 87 91 95 95
rect 87 89 89 91
rect 91 89 95 91
rect 87 81 95 89
rect 87 79 89 81
rect 91 79 95 81
rect 61 55 71 75
rect 73 61 81 75
rect 87 71 95 79
rect 87 69 89 71
rect 91 69 95 71
rect 87 67 95 69
rect 73 59 83 61
rect 73 57 79 59
rect 81 57 83 59
rect 73 55 83 57
rect 91 55 95 67
rect 97 81 107 95
rect 97 79 101 81
rect 103 79 107 81
rect 97 71 107 79
rect 97 69 101 71
rect 103 69 107 71
rect 97 61 107 69
rect 97 59 101 61
rect 103 59 107 61
rect 97 55 107 59
rect 109 91 117 95
rect 109 89 113 91
rect 115 89 117 91
rect 109 81 117 89
rect 109 79 113 81
rect 115 79 117 81
rect 109 71 117 79
rect 109 69 113 71
rect 115 69 117 71
rect 109 61 117 69
rect 109 59 113 61
rect 115 59 117 61
rect 109 55 117 59
<< alu1 >>
rect -2 95 122 100
rect -2 93 5 95
rect 7 93 77 95
rect 79 93 122 95
rect -2 91 122 93
rect -2 89 17 91
rect 19 89 65 91
rect 67 89 89 91
rect 91 89 113 91
rect 115 89 122 91
rect -2 88 122 89
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 62 7 68
rect 4 61 8 62
rect 4 59 5 61
rect 7 59 8 61
rect 4 58 8 59
rect 5 42 7 58
rect 18 51 22 82
rect 28 81 32 82
rect 52 81 56 82
rect 28 79 29 81
rect 31 79 53 81
rect 55 79 56 81
rect 28 78 32 79
rect 52 78 56 79
rect 29 72 31 78
rect 53 72 55 78
rect 28 71 32 72
rect 28 69 29 71
rect 31 69 32 71
rect 28 68 32 69
rect 40 71 44 72
rect 40 69 41 71
rect 43 69 44 71
rect 40 68 44 69
rect 52 71 56 72
rect 52 69 53 71
rect 55 69 56 71
rect 52 68 56 69
rect 41 61 43 68
rect 53 62 55 68
rect 18 49 19 51
rect 21 49 22 51
rect 4 41 8 42
rect 4 39 5 41
rect 7 39 8 41
rect 4 38 8 39
rect 5 22 7 38
rect 18 31 22 49
rect 18 29 19 31
rect 21 29 22 31
rect 4 21 8 22
rect 4 19 5 21
rect 7 19 8 21
rect 4 18 8 19
rect 18 18 22 29
rect 29 59 43 61
rect 52 61 56 62
rect 52 59 53 61
rect 55 59 56 61
rect 29 21 31 59
rect 52 58 56 59
rect 38 51 42 52
rect 68 51 72 82
rect 88 81 92 88
rect 88 79 89 81
rect 91 79 92 81
rect 88 71 92 79
rect 88 69 89 71
rect 91 69 92 71
rect 88 68 92 69
rect 98 81 104 82
rect 98 79 101 81
rect 103 79 104 81
rect 98 78 104 79
rect 112 81 116 88
rect 112 79 113 81
rect 115 79 116 81
rect 98 72 102 78
rect 98 71 104 72
rect 98 69 101 71
rect 103 69 104 71
rect 98 68 104 69
rect 112 71 116 79
rect 112 69 113 71
rect 115 69 116 71
rect 98 62 102 68
rect 98 61 104 62
rect 78 59 82 60
rect 78 57 79 59
rect 81 57 82 59
rect 78 56 82 57
rect 98 59 101 61
rect 103 59 104 61
rect 98 58 104 59
rect 112 61 116 69
rect 112 59 113 61
rect 115 59 116 61
rect 112 58 116 59
rect 38 49 39 51
rect 41 49 69 51
rect 71 49 72 51
rect 38 48 42 49
rect 58 41 62 42
rect 49 39 59 41
rect 61 39 62 41
rect 38 31 42 32
rect 49 31 51 39
rect 58 38 62 39
rect 38 29 39 31
rect 41 29 51 31
rect 68 31 72 49
rect 79 42 81 56
rect 78 41 82 42
rect 78 39 79 41
rect 81 39 82 41
rect 78 38 82 39
rect 88 41 92 42
rect 88 39 89 41
rect 91 39 92 41
rect 88 38 92 39
rect 79 32 81 38
rect 68 29 69 31
rect 71 29 72 31
rect 38 28 42 29
rect 68 28 72 29
rect 78 31 82 32
rect 78 29 79 31
rect 81 29 82 31
rect 78 28 82 29
rect 40 21 44 22
rect 89 21 91 38
rect 29 19 41 21
rect 43 19 91 21
rect 98 22 102 58
rect 98 21 104 22
rect 98 19 101 21
rect 103 19 104 21
rect 40 18 44 19
rect 98 18 104 19
rect 112 21 116 22
rect 112 19 113 21
rect 115 19 116 21
rect 112 12 116 19
rect -2 11 122 12
rect -2 9 17 11
rect 19 9 65 11
rect 67 9 89 11
rect 91 9 113 11
rect 115 9 122 11
rect -2 0 122 9
<< ntie >>
rect 3 95 9 97
rect 75 95 81 97
rect 3 93 5 95
rect 7 93 9 95
rect 3 85 9 93
rect 75 93 77 95
rect 79 93 81 95
rect 75 85 81 93
<< nmos >>
rect 11 15 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
rect 59 5 61 25
rect 71 15 73 25
rect 95 5 97 25
rect 107 5 109 25
<< pmos >>
rect 11 55 13 75
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 59 55 61 95
rect 71 55 73 75
rect 95 55 97 95
rect 107 55 109 95
<< polyct1 >>
rect 19 49 21 51
rect 39 49 41 51
rect 69 49 71 51
rect 5 39 7 41
rect 19 29 21 31
rect 39 29 41 31
rect 59 39 61 41
rect 79 39 81 41
rect 89 39 91 41
rect 69 29 71 31
<< ndifct1 >>
rect 79 29 81 31
rect 5 19 7 21
rect 17 9 19 11
rect 41 19 43 21
rect 65 9 67 11
rect 89 9 91 11
rect 101 19 103 21
rect 113 19 115 21
rect 113 9 115 11
<< ntiect1 >>
rect 5 93 7 95
rect 77 93 79 95
<< pdifct1 >>
rect 17 89 19 91
rect 5 69 7 71
rect 5 59 7 61
rect 29 79 31 81
rect 29 69 31 71
rect 41 69 43 71
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
rect 65 89 67 91
rect 89 89 91 91
rect 89 79 91 81
rect 89 69 91 71
rect 79 57 81 59
rect 101 79 103 81
rect 101 69 103 71
rect 101 59 103 61
rect 113 89 115 91
rect 113 79 115 81
rect 113 69 115 71
rect 113 59 115 61
<< labels >>
rlabel polyct1 20 50 20 50 6 i0
rlabel alu1 60 6 60 6 6 vss
rlabel alu1 60 94 60 94 6 vdd
rlabel alu1 70 55 70 55 6 i1
rlabel alu1 100 50 100 50 6 q
<< end >>
