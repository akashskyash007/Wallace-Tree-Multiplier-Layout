magic
tech scmos
timestamp 1199980656
<< ab >>
rect 0 0 64 88
<< nwell >>
rect -8 40 72 97
<< pwell >>
rect -8 -9 72 40
<< poly >>
rect 5 84 14 86
rect 5 82 7 84
rect 9 82 14 84
rect 5 80 14 82
rect 18 80 27 86
rect 37 80 46 86
rect 50 80 59 86
rect 9 77 11 80
rect 21 77 23 80
rect 41 77 43 80
rect 53 77 55 80
rect 9 48 11 51
rect 21 48 23 51
rect 41 48 43 51
rect 53 48 55 51
rect 2 42 11 48
rect 15 46 30 48
rect 15 44 23 46
rect 25 44 30 46
rect 15 42 30 44
rect 34 46 43 48
rect 34 44 36 46
rect 38 44 43 46
rect 34 42 43 44
rect 47 46 62 48
rect 47 44 55 46
rect 57 44 62 46
rect 47 42 62 44
rect 2 32 17 38
rect 21 36 30 38
rect 21 34 23 36
rect 25 34 30 36
rect 21 32 30 34
rect 34 36 49 38
rect 34 34 36 36
rect 38 34 49 36
rect 34 32 49 34
rect 53 36 62 38
rect 53 34 55 36
rect 57 34 62 36
rect 53 32 62 34
rect 9 29 11 32
rect 21 29 23 32
rect 41 29 43 32
rect 53 29 55 32
rect 9 8 11 11
rect 21 8 23 11
rect 41 8 43 11
rect 53 8 55 11
rect 5 6 14 8
rect 5 4 7 6
rect 9 4 14 6
rect 5 2 14 4
rect 18 2 27 8
rect 37 2 46 8
rect 50 2 59 8
<< ndif >>
rect 2 11 9 29
rect 11 23 21 29
rect 11 21 15 23
rect 17 21 21 23
rect 11 16 21 21
rect 11 14 15 16
rect 17 14 21 16
rect 11 11 21 14
rect 23 24 30 29
rect 23 22 26 24
rect 28 22 30 24
rect 23 17 30 22
rect 23 15 26 17
rect 28 15 30 17
rect 23 11 30 15
rect 34 16 41 29
rect 34 14 36 16
rect 38 14 41 16
rect 34 11 41 14
rect 43 11 53 29
rect 55 24 62 29
rect 55 22 58 24
rect 60 22 62 24
rect 55 17 62 22
rect 55 15 58 17
rect 60 15 62 17
rect 55 11 62 15
<< pdif >>
rect 2 51 9 77
rect 11 74 21 77
rect 11 72 15 74
rect 17 72 21 74
rect 11 67 21 72
rect 11 65 15 67
rect 17 65 21 67
rect 11 51 21 65
rect 23 65 30 77
rect 23 63 26 65
rect 28 63 30 65
rect 23 58 30 63
rect 23 56 26 58
rect 28 56 30 58
rect 23 51 30 56
rect 34 74 41 77
rect 34 72 36 74
rect 38 72 41 74
rect 34 67 41 72
rect 34 65 36 67
rect 38 65 41 67
rect 34 51 41 65
rect 43 65 53 77
rect 43 63 47 65
rect 49 63 53 65
rect 43 57 53 63
rect 43 55 47 57
rect 49 55 53 57
rect 43 51 53 55
rect 55 74 62 77
rect 55 72 58 74
rect 60 72 62 74
rect 55 67 62 72
rect 55 65 58 67
rect 60 65 62 67
rect 55 51 62 65
<< alu1 >>
rect -2 85 2 90
rect 30 85 34 90
rect 62 85 66 90
rect -2 83 -1 85
rect 1 84 31 85
rect 1 83 7 84
rect -2 82 7 83
rect 9 83 31 84
rect 33 83 39 85
rect 9 82 39 83
rect -2 81 39 82
rect 14 74 18 81
rect 14 72 15 74
rect 17 72 18 74
rect 14 67 18 72
rect 35 74 39 81
rect 35 72 36 74
rect 38 72 39 74
rect 35 67 39 72
rect 57 83 63 85
rect 65 83 66 85
rect 57 81 66 83
rect 57 74 61 81
rect 57 72 58 74
rect 60 72 61 74
rect 57 67 61 72
rect 14 65 15 67
rect 17 65 18 67
rect 14 63 18 65
rect 35 65 36 67
rect 38 65 39 67
rect 35 63 39 65
rect 46 65 50 67
rect 46 63 47 65
rect 49 63 50 65
rect 57 65 58 67
rect 60 65 61 67
rect 57 63 61 65
rect 22 46 26 51
rect 22 44 23 46
rect 25 44 26 46
rect 22 36 26 44
rect 22 34 23 36
rect 25 34 26 36
rect 22 29 26 34
rect 14 23 18 25
rect 14 21 15 23
rect 17 21 18 23
rect 14 16 18 21
rect 14 14 15 16
rect 17 14 18 16
rect 14 7 18 14
rect 46 57 50 63
rect 46 55 47 57
rect 49 55 50 57
rect 46 26 50 55
rect 54 46 58 59
rect 54 44 55 46
rect 57 44 58 46
rect 54 36 58 44
rect 54 34 55 36
rect 57 34 58 36
rect 54 32 58 34
rect 46 24 61 26
rect 46 22 58 24
rect 60 22 61 24
rect 46 21 61 22
rect 35 16 39 18
rect 35 14 36 16
rect 38 14 39 16
rect 35 7 39 14
rect 54 17 61 21
rect 54 15 58 17
rect 60 15 61 17
rect 54 13 61 15
rect -2 6 39 7
rect -2 5 7 6
rect -2 3 -1 5
rect 1 4 7 5
rect 9 5 39 6
rect 9 4 31 5
rect 1 3 31 4
rect 33 3 39 5
rect 62 5 66 7
rect 62 3 63 5
rect 65 3 66 5
rect -2 -2 2 3
rect 30 -2 34 3
rect 62 -2 66 3
<< alu2 >>
rect -2 85 66 90
rect -2 83 -1 85
rect 1 83 31 85
rect 33 83 63 85
rect 65 83 66 85
rect -2 80 66 83
rect -2 5 66 8
rect -2 3 -1 5
rect 1 3 31 5
rect 33 3 63 5
rect 65 3 66 5
rect -2 -2 66 3
<< ptie >>
rect -3 5 3 7
rect -3 3 -1 5
rect 1 3 3 5
rect -3 0 3 3
rect 29 5 35 7
rect 29 3 31 5
rect 33 3 35 5
rect 29 0 35 3
rect 61 5 67 7
rect 61 3 63 5
rect 65 3 67 5
rect 61 0 67 3
<< ntie >>
rect -3 85 3 88
rect -3 83 -1 85
rect 1 83 3 85
rect -3 81 3 83
rect 29 85 35 88
rect 29 83 31 85
rect 33 83 35 85
rect 29 81 35 83
rect 61 85 67 88
rect 61 83 63 85
rect 65 83 67 85
rect 61 81 67 83
<< nmos >>
rect 9 11 11 29
rect 21 11 23 29
rect 41 11 43 29
rect 53 11 55 29
<< pmos >>
rect 9 51 11 77
rect 21 51 23 77
rect 41 51 43 77
rect 53 51 55 77
<< polyct0 >>
rect 36 44 38 46
rect 36 34 38 36
<< polyct1 >>
rect 7 82 9 84
rect 23 44 25 46
rect 55 44 57 46
rect 23 34 25 36
rect 55 34 57 36
rect 7 4 9 6
<< ndifct0 >>
rect 26 22 28 24
rect 26 15 28 17
<< ndifct1 >>
rect 15 21 17 23
rect 15 14 17 16
rect 36 14 38 16
rect 58 22 60 24
rect 58 15 60 17
<< ntiect1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
<< ptiect1 >>
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< pdifct0 >>
rect 26 63 28 65
rect 26 56 28 58
<< pdifct1 >>
rect 15 72 17 74
rect 15 65 17 67
rect 36 72 38 74
rect 36 65 38 67
rect 47 63 49 65
rect 47 55 49 57
rect 58 72 60 74
rect 58 65 60 67
<< alu0 >>
rect 25 65 29 67
rect 25 63 26 65
rect 28 63 29 65
rect 25 58 29 63
rect 25 56 26 58
rect 28 56 39 58
rect 25 54 39 56
rect 35 46 39 54
rect 35 44 36 46
rect 38 44 39 46
rect 35 36 39 44
rect 35 34 36 36
rect 38 34 39 36
rect 35 26 39 34
rect 25 24 39 26
rect 25 22 26 24
rect 28 22 39 24
rect 25 17 29 22
rect 25 15 26 17
rect 28 15 29 17
rect 25 13 29 15
<< via1 >>
rect -1 83 1 85
rect 31 83 33 85
rect 63 83 65 85
rect -1 3 1 5
rect 31 3 33 5
rect 63 3 65 5
<< labels >>
rlabel alu1 24 40 24 40 6 a
rlabel alu1 56 20 56 20 6 z
rlabel alu1 56 48 56 48 6 b
rlabel alu1 48 44 48 44 6 z
rlabel via1 32 4 32 4 6 vss
rlabel via1 32 84 32 84 6 vdd
<< end >>
