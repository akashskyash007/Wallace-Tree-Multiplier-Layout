magic
tech scmos
timestamp 1199202808
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 10 68 62 70
rect 10 59 12 68
rect 20 59 22 64
rect 30 59 32 64
rect 40 59 42 64
rect 50 59 52 64
rect 60 59 62 68
rect 10 31 12 39
rect 20 35 22 39
rect 30 35 32 39
rect 40 35 42 39
rect 50 35 52 39
rect 60 35 62 39
rect 20 33 26 35
rect 20 31 22 33
rect 24 31 26 33
rect 10 29 16 31
rect 20 29 26 31
rect 30 33 42 35
rect 30 31 35 33
rect 37 31 42 33
rect 30 29 42 31
rect 46 33 52 35
rect 46 31 48 33
rect 50 31 52 33
rect 46 29 52 31
rect 56 33 63 35
rect 56 31 59 33
rect 61 31 63 33
rect 56 29 63 31
rect 14 26 16 29
rect 22 26 24 29
rect 30 26 32 29
rect 40 26 42 29
rect 48 26 50 29
rect 56 26 58 29
rect 14 2 16 6
rect 22 2 24 6
rect 30 2 32 6
rect 40 2 42 6
rect 48 2 50 6
rect 56 2 58 6
<< ndif >>
rect 6 10 14 26
rect 6 8 9 10
rect 11 8 14 10
rect 6 6 14 8
rect 16 6 22 26
rect 24 6 30 26
rect 32 17 40 26
rect 32 15 35 17
rect 37 15 40 17
rect 32 6 40 15
rect 42 6 48 26
rect 50 6 56 26
rect 58 17 66 26
rect 58 15 61 17
rect 63 15 66 17
rect 58 10 66 15
rect 58 8 61 10
rect 63 8 66 10
rect 58 6 66 8
<< pdif >>
rect 2 57 10 59
rect 2 55 4 57
rect 6 55 10 57
rect 2 50 10 55
rect 2 48 4 50
rect 6 48 10 50
rect 2 39 10 48
rect 12 57 20 59
rect 12 55 15 57
rect 17 55 20 57
rect 12 50 20 55
rect 12 48 15 50
rect 17 48 20 50
rect 12 39 20 48
rect 22 57 30 59
rect 22 55 25 57
rect 27 55 30 57
rect 22 39 30 55
rect 32 57 40 59
rect 32 55 35 57
rect 37 55 40 57
rect 32 50 40 55
rect 32 48 35 50
rect 37 48 40 50
rect 32 39 40 48
rect 42 57 50 59
rect 42 55 45 57
rect 47 55 50 57
rect 42 39 50 55
rect 52 57 60 59
rect 52 55 55 57
rect 57 55 60 57
rect 52 50 60 55
rect 52 48 55 50
rect 57 48 60 50
rect 52 39 60 48
rect 62 57 70 59
rect 62 55 66 57
rect 68 55 70 57
rect 62 39 70 55
<< alu1 >>
rect -2 64 74 72
rect 14 57 18 59
rect 14 55 15 57
rect 17 55 18 57
rect 14 51 18 55
rect 34 57 38 59
rect 34 55 35 57
rect 37 55 38 57
rect 10 50 18 51
rect 34 50 38 55
rect 54 57 58 59
rect 54 55 55 57
rect 57 55 58 57
rect 54 50 58 55
rect 10 48 15 50
rect 17 48 35 50
rect 37 48 55 50
rect 57 48 58 50
rect 10 46 58 48
rect 10 18 14 46
rect 22 38 52 42
rect 22 35 26 38
rect 18 33 26 35
rect 18 31 22 33
rect 24 31 26 33
rect 18 29 26 31
rect 33 33 39 34
rect 33 31 35 33
rect 37 31 39 33
rect 33 26 39 31
rect 46 33 52 38
rect 66 35 70 51
rect 46 31 48 33
rect 50 31 52 33
rect 46 30 52 31
rect 58 33 70 35
rect 58 31 59 33
rect 61 31 70 33
rect 58 29 70 31
rect 33 22 47 26
rect 10 17 39 18
rect 10 15 35 17
rect 37 15 39 17
rect 10 14 39 15
rect -2 0 74 8
<< nmos >>
rect 14 6 16 26
rect 22 6 24 26
rect 30 6 32 26
rect 40 6 42 26
rect 48 6 50 26
rect 56 6 58 26
<< pmos >>
rect 10 39 12 59
rect 20 39 22 59
rect 30 39 32 59
rect 40 39 42 59
rect 50 39 52 59
rect 60 39 62 59
<< polyct1 >>
rect 22 31 24 33
rect 35 31 37 33
rect 48 31 50 33
rect 59 31 61 33
<< ndifct0 >>
rect 9 8 11 10
rect 61 15 63 17
rect 61 8 63 10
<< ndifct1 >>
rect 35 15 37 17
<< pdifct0 >>
rect 4 55 6 57
rect 4 48 6 50
rect 25 55 27 57
rect 45 55 47 57
rect 66 55 68 57
<< pdifct1 >>
rect 15 55 17 57
rect 15 48 17 50
rect 35 55 37 57
rect 35 48 37 50
rect 55 55 57 57
rect 55 48 57 50
<< alu0 >>
rect 3 57 7 64
rect 3 55 4 57
rect 6 55 7 57
rect 3 50 7 55
rect 23 57 29 64
rect 23 55 25 57
rect 27 55 29 57
rect 23 54 29 55
rect 3 48 4 50
rect 6 48 7 50
rect 3 46 7 48
rect 43 57 49 64
rect 43 55 45 57
rect 47 55 49 57
rect 43 54 49 55
rect 64 57 70 64
rect 64 55 66 57
rect 68 55 70 57
rect 64 54 70 55
rect 59 17 65 18
rect 59 15 61 17
rect 63 15 65 17
rect 7 10 13 11
rect 7 8 9 10
rect 11 8 13 10
rect 59 10 65 15
rect 59 8 61 10
rect 63 8 65 10
<< labels >>
rlabel alu1 12 36 12 36 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 32 20 32 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel ndifct1 36 16 36 16 6 z
rlabel alu1 36 28 36 28 6 c
rlabel alu1 44 24 44 24 6 c
rlabel alu1 44 40 44 40 6 b
rlabel alu1 36 40 36 40 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel polyct1 60 32 60 32 6 a
rlabel alu1 68 40 68 40 6 a
<< end >>
