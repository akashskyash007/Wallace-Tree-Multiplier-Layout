magic
tech scmos
timestamp 1199201990
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 65 31 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 33 22 35
rect 9 31 18 33
rect 20 31 22 33
rect 9 29 22 31
rect 26 33 32 35
rect 26 31 28 33
rect 30 31 32 33
rect 26 29 32 31
rect 9 26 11 29
rect 19 26 21 29
rect 29 26 31 29
rect 9 7 11 12
rect 19 7 21 12
rect 29 6 31 11
<< ndif >>
rect 2 23 9 26
rect 2 21 4 23
rect 6 21 9 23
rect 2 16 9 21
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 17 19 26
rect 11 15 14 17
rect 16 15 19 17
rect 11 12 19 15
rect 21 16 29 26
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 23 11 29 12
rect 31 24 38 26
rect 31 22 34 24
rect 36 22 38 24
rect 31 17 38 22
rect 31 15 34 17
rect 36 15 38 17
rect 31 13 38 15
rect 31 11 36 13
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 65 27 66
rect 21 63 29 65
rect 21 61 24 63
rect 26 61 29 63
rect 21 56 29 61
rect 21 54 24 56
rect 26 54 29 56
rect 21 38 29 54
rect 31 58 36 65
rect 31 56 38 58
rect 31 54 34 56
rect 36 54 38 56
rect 31 49 38 54
rect 31 47 34 49
rect 36 47 38 49
rect 31 45 38 47
rect 31 38 36 45
<< alu1 >>
rect -2 64 42 72
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 50 17 55
rect 2 48 14 50
rect 16 48 17 50
rect 2 46 17 48
rect 2 33 6 46
rect 17 38 31 42
rect 2 29 14 33
rect 10 19 14 29
rect 26 33 31 38
rect 26 31 28 33
rect 30 31 31 33
rect 26 29 31 31
rect 10 17 17 19
rect 10 15 14 17
rect 16 15 17 17
rect 10 13 17 15
rect -2 0 42 8
<< nmos >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 11 31 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 65
<< polyct0 >>
rect 18 31 20 33
<< polyct1 >>
rect 28 31 30 33
<< ndifct0 >>
rect 4 21 6 23
rect 4 14 6 16
rect 24 14 26 16
rect 34 22 36 24
rect 34 15 36 17
<< ndifct1 >>
rect 14 15 16 17
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 24 61 26 63
rect 24 54 26 56
rect 34 54 36 56
rect 34 47 36 49
<< pdifct1 >>
rect 14 55 16 57
rect 14 48 16 50
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 23 63 27 64
rect 23 61 24 63
rect 26 61 27 63
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 23 56 27 61
rect 23 54 24 56
rect 26 54 27 56
rect 23 52 27 54
rect 33 56 38 58
rect 33 54 34 56
rect 36 54 38 56
rect 33 49 38 54
rect 33 47 34 49
rect 36 47 38 49
rect 33 45 38 47
rect 17 33 21 35
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 16 7 21
rect 3 14 4 16
rect 6 14 7 16
rect 3 8 7 14
rect 17 31 18 33
rect 20 31 21 33
rect 17 26 21 31
rect 34 26 38 45
rect 17 24 38 26
rect 17 22 34 24
rect 36 22 38 24
rect 23 16 27 18
rect 23 14 24 16
rect 26 14 27 16
rect 23 8 27 14
rect 33 17 37 22
rect 33 15 34 17
rect 36 15 37 17
rect 33 13 37 15
<< labels >>
rlabel alu0 19 28 19 28 6 an
rlabel alu0 35 19 35 19 6 an
rlabel alu0 36 40 36 40 6 an
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 28 36 28 36 6 a
rlabel alu1 20 40 20 40 6 a
rlabel alu1 20 68 20 68 6 vdd
<< end >>
