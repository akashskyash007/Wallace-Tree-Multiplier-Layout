magic
tech scmos
timestamp 1199543209
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -2 48 92 104
<< pwell >>
rect -2 -4 92 48
<< poly >>
rect 23 95 25 98
rect 35 95 37 98
rect 47 95 49 98
rect 59 95 61 98
rect 11 85 13 88
rect 11 53 13 65
rect 71 85 73 88
rect 23 53 25 55
rect 11 51 25 53
rect 35 53 37 55
rect 35 51 43 53
rect 17 49 19 51
rect 21 49 23 51
rect 17 47 23 49
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 3 41 9 43
rect 47 41 49 55
rect 59 43 61 55
rect 71 53 73 65
rect 67 51 73 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 3 39 5 41
rect 7 39 49 41
rect 3 37 9 39
rect 17 31 23 33
rect 17 29 19 31
rect 21 29 23 31
rect 37 31 43 33
rect 37 29 39 31
rect 41 29 43 31
rect 11 27 25 29
rect 11 25 13 27
rect 23 25 25 27
rect 35 27 43 29
rect 35 25 37 27
rect 47 25 49 39
rect 57 41 63 43
rect 77 41 83 43
rect 57 39 59 41
rect 61 39 79 41
rect 81 39 83 41
rect 57 37 63 39
rect 77 37 83 39
rect 67 31 73 33
rect 67 29 69 31
rect 71 29 73 31
rect 59 27 73 29
rect 59 25 61 27
rect 71 25 73 27
rect 11 12 13 15
rect 71 12 73 15
rect 23 2 25 5
rect 35 2 37 5
rect 47 2 49 5
rect 59 2 61 5
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 15 11 23 15
rect 15 9 17 11
rect 19 9 23 11
rect 15 5 23 9
rect 25 5 35 25
rect 37 21 47 25
rect 37 19 41 21
rect 43 19 47 21
rect 37 5 47 19
rect 49 5 59 25
rect 61 15 71 25
rect 73 21 83 25
rect 73 19 79 21
rect 81 19 83 21
rect 73 15 83 19
rect 61 11 69 15
rect 61 9 65 11
rect 67 9 69 11
rect 61 5 69 9
<< pdif >>
rect 15 91 23 95
rect 15 89 17 91
rect 19 89 23 91
rect 15 85 23 89
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 65 11 69
rect 13 65 23 85
rect 15 55 23 65
rect 25 81 35 95
rect 25 79 29 81
rect 31 79 35 81
rect 25 55 35 79
rect 37 71 47 95
rect 37 69 41 71
rect 43 69 47 71
rect 37 55 47 69
rect 49 81 59 95
rect 49 79 53 81
rect 55 79 59 81
rect 49 71 59 79
rect 49 69 53 71
rect 55 69 59 71
rect 49 61 59 69
rect 49 59 53 61
rect 55 59 59 61
rect 49 55 59 59
rect 61 91 69 95
rect 61 89 65 91
rect 67 89 69 91
rect 61 85 69 89
rect 61 65 71 85
rect 73 81 83 85
rect 73 79 79 81
rect 81 79 83 81
rect 73 71 83 79
rect 73 69 79 71
rect 81 69 83 71
rect 73 65 83 69
rect 61 55 69 65
<< alu1 >>
rect -2 95 92 100
rect -2 93 77 95
rect 79 93 92 95
rect -2 91 92 93
rect -2 89 17 91
rect 19 89 65 91
rect 67 89 92 91
rect -2 88 92 89
rect 4 81 8 82
rect 4 79 5 81
rect 7 79 8 81
rect 4 78 8 79
rect 5 72 7 78
rect 4 71 8 72
rect 4 69 5 71
rect 7 69 8 71
rect 4 68 8 69
rect 5 42 7 68
rect 18 51 22 82
rect 28 81 32 82
rect 52 81 56 82
rect 28 79 29 81
rect 31 79 53 81
rect 55 79 56 81
rect 28 78 32 79
rect 52 78 56 79
rect 53 72 55 78
rect 18 49 19 51
rect 21 49 22 51
rect 4 41 8 42
rect 4 39 5 41
rect 7 39 8 41
rect 4 38 8 39
rect 5 22 7 38
rect 18 31 22 49
rect 18 29 19 31
rect 21 29 22 31
rect 4 21 8 22
rect 4 19 5 21
rect 7 19 8 21
rect 4 18 8 19
rect 18 18 22 29
rect 28 71 44 72
rect 28 69 41 71
rect 43 69 44 71
rect 28 68 44 69
rect 52 71 56 72
rect 52 69 53 71
rect 55 69 56 71
rect 52 68 56 69
rect 28 22 32 68
rect 53 62 55 68
rect 52 61 56 62
rect 52 59 53 61
rect 55 59 56 61
rect 52 58 56 59
rect 38 51 42 52
rect 68 51 72 82
rect 78 81 82 82
rect 78 79 79 81
rect 81 79 82 81
rect 78 78 82 79
rect 79 72 81 78
rect 78 71 82 72
rect 78 69 79 71
rect 81 69 82 71
rect 78 68 82 69
rect 38 49 39 51
rect 41 49 69 51
rect 71 49 72 51
rect 38 48 42 49
rect 58 41 62 42
rect 49 39 59 41
rect 61 39 62 41
rect 38 31 42 32
rect 49 31 51 39
rect 58 38 62 39
rect 38 29 39 31
rect 41 29 51 31
rect 68 31 72 49
rect 79 42 81 68
rect 78 41 82 42
rect 78 39 79 41
rect 81 39 82 41
rect 78 38 82 39
rect 68 29 69 31
rect 71 29 72 31
rect 38 28 42 29
rect 28 21 44 22
rect 28 19 41 21
rect 43 19 44 21
rect 28 18 44 19
rect 68 18 72 29
rect 79 22 81 38
rect 78 21 82 22
rect 78 19 79 21
rect 81 19 82 21
rect 78 18 82 19
rect -2 11 92 12
rect -2 9 17 11
rect 19 9 65 11
rect 67 9 92 11
rect -2 7 92 9
rect -2 5 77 7
rect 79 5 92 7
rect -2 0 92 5
<< ptie >>
rect 75 7 87 9
rect 75 5 77 7
rect 79 5 87 7
rect 75 3 87 5
<< ntie >>
rect 75 95 87 97
rect 75 93 77 95
rect 79 93 87 95
rect 75 91 87 93
<< nmos >>
rect 11 15 13 25
rect 23 5 25 25
rect 35 5 37 25
rect 47 5 49 25
rect 59 5 61 25
rect 71 15 73 25
<< pmos >>
rect 11 65 13 85
rect 23 55 25 95
rect 35 55 37 95
rect 47 55 49 95
rect 59 55 61 95
rect 71 65 73 85
<< polyct1 >>
rect 19 49 21 51
rect 39 49 41 51
rect 69 49 71 51
rect 5 39 7 41
rect 19 29 21 31
rect 39 29 41 31
rect 59 39 61 41
rect 79 39 81 41
rect 69 29 71 31
<< ndifct1 >>
rect 5 19 7 21
rect 17 9 19 11
rect 41 19 43 21
rect 79 19 81 21
rect 65 9 67 11
<< ntiect1 >>
rect 77 93 79 95
<< ptiect1 >>
rect 77 5 79 7
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 5 69 7 71
rect 29 79 31 81
rect 41 69 43 71
rect 53 79 55 81
rect 53 69 55 71
rect 53 59 55 61
rect 65 89 67 91
rect 79 79 81 81
rect 79 69 81 71
<< labels >>
rlabel alu1 30 45 30 45 6 nq
rlabel polyct1 20 50 20 50 6 i0
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 45 94 45 94 6 vdd
rlabel polyct1 70 50 70 50 6 i1
<< end >>
