magic
tech scmos
timestamp 1199202193
<< ab >>
rect 0 0 168 80
<< nwell >>
rect -5 36 173 88
<< pwell >>
rect -5 -8 173 36
<< poly >>
rect 9 70 11 74
rect 19 70 21 74
rect 29 70 31 74
rect 39 70 41 74
rect 49 70 51 74
rect 59 70 61 74
rect 69 70 71 74
rect 76 70 78 74
rect 89 70 91 74
rect 96 70 98 74
rect 106 70 108 74
rect 113 70 115 74
rect 125 70 127 74
rect 135 70 137 74
rect 145 70 147 74
rect 9 37 11 42
rect 19 37 21 42
rect 29 37 31 42
rect 9 35 31 37
rect 9 30 11 35
rect 19 30 21 35
rect 29 30 31 35
rect 39 39 41 42
rect 49 39 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 76 39 78 42
rect 89 39 91 42
rect 39 37 61 39
rect 39 30 41 37
rect 49 35 57 37
rect 59 35 61 37
rect 49 33 61 35
rect 66 37 72 39
rect 66 35 68 37
rect 70 35 72 37
rect 66 33 72 35
rect 76 37 91 39
rect 76 35 83 37
rect 85 35 91 37
rect 76 33 91 35
rect 49 30 51 33
rect 59 30 61 33
rect 69 30 71 33
rect 76 30 78 33
rect 89 30 91 33
rect 96 39 98 42
rect 106 39 108 42
rect 96 37 108 39
rect 96 35 98 37
rect 100 35 108 37
rect 96 33 108 35
rect 96 30 98 33
rect 106 30 108 33
rect 113 39 115 42
rect 125 39 127 42
rect 135 39 137 42
rect 145 39 147 42
rect 113 37 147 39
rect 113 35 115 37
rect 117 35 128 37
rect 113 33 128 35
rect 113 30 115 33
rect 126 30 128 33
rect 136 30 138 37
rect 9 11 11 16
rect 19 11 21 16
rect 29 8 31 16
rect 39 12 41 16
rect 49 12 51 16
rect 59 12 61 16
rect 69 8 71 16
rect 76 11 78 16
rect 89 11 91 16
rect 96 11 98 16
rect 106 11 108 16
rect 113 11 115 16
rect 29 6 71 8
rect 126 6 128 10
rect 136 6 138 10
<< ndif >>
rect 2 27 9 30
rect 2 25 4 27
rect 6 25 9 27
rect 2 20 9 25
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 21 19 26
rect 11 19 14 21
rect 16 19 19 21
rect 11 16 19 19
rect 21 20 29 30
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 21 39 26
rect 31 19 34 21
rect 36 19 39 21
rect 31 16 39 19
rect 41 28 49 30
rect 41 26 44 28
rect 46 26 49 28
rect 41 16 49 26
rect 51 21 59 30
rect 51 19 54 21
rect 56 19 59 21
rect 51 16 59 19
rect 61 28 69 30
rect 61 26 64 28
rect 66 26 69 28
rect 61 16 69 26
rect 71 16 76 30
rect 78 16 89 30
rect 91 16 96 30
rect 98 28 106 30
rect 98 26 101 28
rect 103 26 106 28
rect 98 16 106 26
rect 108 16 113 30
rect 115 16 126 30
rect 80 11 87 16
rect 117 14 126 16
rect 117 12 119 14
rect 121 12 126 14
rect 80 9 82 11
rect 84 9 87 11
rect 117 10 126 12
rect 128 28 136 30
rect 128 26 131 28
rect 133 26 136 28
rect 128 21 136 26
rect 128 19 131 21
rect 133 19 136 21
rect 128 10 136 19
rect 138 22 146 30
rect 138 20 141 22
rect 143 20 146 22
rect 138 14 146 20
rect 138 12 141 14
rect 143 12 146 14
rect 138 10 146 12
rect 80 7 87 9
<< pdif >>
rect 2 68 9 70
rect 2 66 4 68
rect 6 66 9 68
rect 2 61 9 66
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 42 9 52
rect 11 61 19 70
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 68 29 70
rect 21 66 24 68
rect 26 66 29 68
rect 21 61 29 66
rect 21 59 24 61
rect 26 59 29 61
rect 21 42 29 59
rect 31 61 39 70
rect 31 59 34 61
rect 36 59 39 61
rect 31 54 39 59
rect 31 52 34 54
rect 36 52 39 54
rect 31 42 39 52
rect 41 53 49 70
rect 41 51 44 53
rect 46 51 49 53
rect 41 42 49 51
rect 51 61 59 70
rect 51 59 54 61
rect 56 59 59 61
rect 51 42 59 59
rect 61 53 69 70
rect 61 51 64 53
rect 66 51 69 53
rect 61 42 69 51
rect 71 42 76 70
rect 78 68 89 70
rect 78 66 82 68
rect 84 66 89 68
rect 78 42 89 66
rect 91 42 96 70
rect 98 53 106 70
rect 98 51 101 53
rect 103 51 106 53
rect 98 42 106 51
rect 108 42 113 70
rect 115 68 125 70
rect 115 66 119 68
rect 121 66 125 68
rect 115 42 125 66
rect 127 61 135 70
rect 127 59 130 61
rect 132 59 135 61
rect 127 54 135 59
rect 127 52 130 54
rect 132 52 135 54
rect 127 42 135 52
rect 137 68 145 70
rect 137 66 140 68
rect 142 66 145 68
rect 137 61 145 66
rect 137 59 140 61
rect 142 59 145 61
rect 137 42 145 59
rect 147 55 152 70
rect 147 53 154 55
rect 147 51 150 53
rect 152 51 154 53
rect 147 46 154 51
rect 147 44 150 46
rect 152 44 154 46
rect 147 42 154 44
<< alu1 >>
rect -2 81 170 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 170 81
rect -2 68 170 79
rect 42 53 126 54
rect 42 51 44 53
rect 46 51 64 53
rect 66 51 101 53
rect 103 51 126 53
rect 42 50 126 51
rect 42 29 46 50
rect 57 39 63 46
rect 81 42 118 46
rect 50 37 63 39
rect 50 35 57 37
rect 59 35 63 37
rect 50 33 63 35
rect 67 37 77 39
rect 67 35 68 37
rect 70 35 77 37
rect 67 33 77 35
rect 81 37 87 42
rect 81 35 83 37
rect 85 35 87 37
rect 81 34 87 35
rect 91 37 103 38
rect 91 35 98 37
rect 100 35 103 37
rect 91 34 103 35
rect 114 37 118 42
rect 114 35 115 37
rect 117 35 118 37
rect 73 30 77 33
rect 91 30 95 34
rect 114 33 118 35
rect 42 28 68 29
rect 42 26 44 28
rect 46 26 64 28
rect 66 26 68 28
rect 73 26 95 30
rect 122 29 126 50
rect 99 28 126 29
rect 99 26 101 28
rect 103 26 126 28
rect 42 25 68 26
rect 99 25 126 26
rect -2 11 170 12
rect -2 9 82 11
rect 84 9 170 11
rect -2 1 170 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 170 1
rect -2 -2 170 -1
<< ptie >>
rect 0 1 168 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 168 1
rect 0 -3 168 -1
<< ntie >>
rect 0 81 168 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 168 81
rect 0 77 168 79
<< nmos >>
rect 9 16 11 30
rect 19 16 21 30
rect 29 16 31 30
rect 39 16 41 30
rect 49 16 51 30
rect 59 16 61 30
rect 69 16 71 30
rect 76 16 78 30
rect 89 16 91 30
rect 96 16 98 30
rect 106 16 108 30
rect 113 16 115 30
rect 126 10 128 30
rect 136 10 138 30
<< pmos >>
rect 9 42 11 70
rect 19 42 21 70
rect 29 42 31 70
rect 39 42 41 70
rect 49 42 51 70
rect 59 42 61 70
rect 69 42 71 70
rect 76 42 78 70
rect 89 42 91 70
rect 96 42 98 70
rect 106 42 108 70
rect 113 42 115 70
rect 125 42 127 70
rect 135 42 137 70
rect 145 42 147 70
<< polyct1 >>
rect 57 35 59 37
rect 68 35 70 37
rect 83 35 85 37
rect 98 35 100 37
rect 115 35 117 37
<< ndifct0 >>
rect 4 25 6 27
rect 4 18 6 20
rect 14 26 16 28
rect 14 19 16 21
rect 24 18 26 20
rect 34 26 36 28
rect 34 19 36 21
rect 54 19 56 21
rect 119 12 121 14
rect 131 26 133 28
rect 131 19 133 21
rect 141 20 143 22
rect 141 12 143 14
<< ndifct1 >>
rect 44 26 46 28
rect 64 26 66 28
rect 101 26 103 28
rect 82 9 84 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 4 52 6 54
rect 14 59 16 61
rect 14 52 16 54
rect 24 66 26 68
rect 24 59 26 61
rect 34 59 36 61
rect 34 52 36 54
rect 54 59 56 61
rect 82 66 84 68
rect 119 66 121 68
rect 130 59 132 61
rect 130 52 132 54
rect 140 66 142 68
rect 140 59 142 61
rect 150 51 152 53
rect 150 44 152 46
<< pdifct1 >>
rect 44 51 46 53
rect 64 51 66 53
rect 101 51 103 53
<< alu0 >>
rect 3 66 4 68
rect 6 66 7 68
rect 3 61 7 66
rect 22 66 24 68
rect 26 66 28 68
rect 3 59 4 61
rect 6 59 7 61
rect 3 54 7 59
rect 3 52 4 54
rect 6 52 7 54
rect 3 50 7 52
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 61 28 66
rect 80 66 82 68
rect 84 66 86 68
rect 80 65 86 66
rect 117 66 119 68
rect 121 66 123 68
rect 117 65 123 66
rect 138 66 140 68
rect 142 66 144 68
rect 22 59 24 61
rect 26 59 28 61
rect 22 58 28 59
rect 32 61 134 62
rect 32 59 34 61
rect 36 59 54 61
rect 56 59 130 61
rect 132 59 134 61
rect 32 58 134 59
rect 138 61 144 66
rect 138 59 140 61
rect 142 59 144 61
rect 157 59 161 68
rect 138 58 144 59
rect 32 54 37 58
rect 129 54 134 58
rect 13 52 14 54
rect 16 52 34 54
rect 36 52 37 54
rect 13 50 37 52
rect 129 52 130 54
rect 132 53 154 54
rect 132 52 150 53
rect 129 51 150 52
rect 152 51 154 53
rect 129 50 154 51
rect 3 27 7 29
rect 3 25 4 27
rect 6 25 7 27
rect 3 20 7 25
rect 3 18 4 20
rect 6 18 7 20
rect 3 12 7 18
rect 13 28 37 30
rect 13 26 14 28
rect 16 26 34 28
rect 36 26 37 28
rect 13 21 17 26
rect 32 22 37 26
rect 148 46 154 50
rect 148 44 150 46
rect 152 44 154 46
rect 148 43 154 44
rect 130 28 135 30
rect 130 26 131 28
rect 133 26 135 28
rect 130 22 135 26
rect 13 19 14 21
rect 16 19 17 21
rect 13 17 17 19
rect 23 20 27 22
rect 23 18 24 20
rect 26 18 27 20
rect 32 21 135 22
rect 32 19 34 21
rect 36 19 54 21
rect 56 19 131 21
rect 133 19 135 21
rect 32 18 135 19
rect 140 22 144 24
rect 140 20 141 22
rect 143 20 144 22
rect 23 12 27 18
rect 117 14 123 15
rect 117 12 119 14
rect 121 12 123 14
rect 140 14 144 20
rect 140 12 141 14
rect 143 12 144 14
rect 154 12 158 21
<< labels >>
rlabel alu0 15 23 15 23 6 n3
rlabel alu0 15 56 15 56 6 n1
rlabel alu0 34 24 34 24 6 n3
rlabel alu0 34 56 34 56 6 n1
rlabel alu0 132 24 132 24 6 n3
rlabel alu0 83 20 83 20 6 n3
rlabel alu0 151 48 151 48 6 n1
rlabel alu0 141 52 141 52 6 n1
rlabel alu0 131 56 131 56 6 n1
rlabel alu0 83 60 83 60 6 n1
rlabel alu1 52 36 52 36 6 c
rlabel alu1 60 40 60 40 6 c
rlabel alu1 44 36 44 36 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 84 6 84 6 6 vss
rlabel alu1 76 28 76 28 6 b
rlabel alu1 84 28 84 28 6 b
rlabel alu1 92 28 92 28 6 b
rlabel alu1 84 40 84 40 6 a
rlabel alu1 92 44 92 44 6 a
rlabel alu1 76 52 76 52 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 92 52 92 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 84 74 84 74 6 vdd
rlabel alu1 100 36 100 36 6 b
rlabel alu1 100 44 100 44 6 a
rlabel alu1 108 44 108 44 6 a
rlabel polyct1 116 36 116 36 6 a
rlabel alu1 124 36 124 36 6 z
rlabel alu1 108 52 108 52 6 z
rlabel alu1 116 52 116 52 6 z
rlabel alu1 100 52 100 52 6 z
<< end >>
