magic
tech scmos
timestamp 1199203492
<< ab >>
rect 0 0 168 80
<< nwell >>
rect -5 36 173 88
<< pwell >>
rect -5 -8 173 36
<< poly >>
rect 9 70 11 74
rect 16 70 18 74
rect 26 70 28 74
rect 33 70 35 74
rect 43 70 45 74
rect 50 70 52 74
rect 60 70 62 74
rect 67 70 69 74
rect 77 70 79 74
rect 87 70 89 74
rect 117 70 119 74
rect 127 70 129 74
rect 137 70 139 74
rect 147 70 149 74
rect 97 61 99 65
rect 107 61 109 65
rect 157 61 159 65
rect 9 39 11 42
rect 16 39 18 42
rect 26 39 28 42
rect 33 39 35 42
rect 43 39 45 42
rect 5 37 11 39
rect 5 35 7 37
rect 9 35 11 37
rect 5 33 11 35
rect 15 37 28 39
rect 32 37 45 39
rect 50 39 52 42
rect 60 39 62 42
rect 67 39 69 42
rect 77 39 79 42
rect 87 39 89 42
rect 97 39 99 42
rect 50 37 62 39
rect 66 37 72 39
rect 15 22 17 37
rect 32 35 34 37
rect 36 35 38 37
rect 32 33 38 35
rect 26 29 28 33
rect 36 29 38 33
rect 46 29 48 33
rect 56 29 58 37
rect 66 35 68 37
rect 70 35 72 37
rect 66 33 72 35
rect 76 37 99 39
rect 66 29 68 33
rect 76 29 78 37
rect 88 35 95 37
rect 97 35 99 37
rect 88 33 99 35
rect 107 39 109 42
rect 117 39 119 42
rect 127 39 129 42
rect 137 39 139 42
rect 147 39 149 42
rect 157 39 159 42
rect 107 37 129 39
rect 107 35 123 37
rect 125 35 129 37
rect 107 33 129 35
rect 133 37 159 39
rect 133 35 135 37
rect 137 35 139 37
rect 133 33 139 35
rect 88 29 90 33
rect 109 30 111 33
rect 119 30 121 33
rect 11 20 17 22
rect 11 18 13 20
rect 15 18 17 20
rect 11 16 17 18
rect 15 8 17 16
rect 26 15 28 18
rect 36 15 38 18
rect 26 13 38 15
rect 46 8 48 11
rect 56 8 58 11
rect 66 8 68 13
rect 15 6 58 8
rect 76 6 78 10
rect 88 6 90 10
rect 109 6 111 11
rect 119 6 121 11
<< ndif >>
rect 19 27 26 29
rect 19 25 21 27
rect 23 25 26 27
rect 19 23 26 25
rect 21 18 26 23
rect 28 22 36 29
rect 28 20 31 22
rect 33 20 36 22
rect 28 18 36 20
rect 38 27 46 29
rect 38 25 41 27
rect 43 25 46 27
rect 38 18 46 25
rect 41 11 46 18
rect 48 27 56 29
rect 48 25 51 27
rect 53 25 56 27
rect 48 11 56 25
rect 58 27 66 29
rect 58 25 61 27
rect 63 25 66 27
rect 58 13 66 25
rect 68 20 76 29
rect 68 18 71 20
rect 73 18 76 20
rect 68 13 76 18
rect 58 11 63 13
rect 71 10 76 13
rect 78 11 88 29
rect 78 10 82 11
rect 80 9 82 10
rect 84 10 88 11
rect 90 22 95 29
rect 90 20 97 22
rect 90 18 93 20
rect 95 18 97 20
rect 90 16 97 18
rect 90 10 95 16
rect 101 11 109 30
rect 111 28 119 30
rect 111 26 114 28
rect 116 26 119 28
rect 111 11 119 26
rect 121 11 129 30
rect 84 9 86 10
rect 80 7 86 9
rect 101 9 103 11
rect 105 9 107 11
rect 101 7 107 9
rect 123 9 125 11
rect 127 9 129 11
rect 123 7 129 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 42 16 70
rect 18 68 26 70
rect 18 66 21 68
rect 23 66 26 68
rect 18 42 26 66
rect 28 42 33 70
rect 35 61 43 70
rect 35 59 38 61
rect 40 59 43 61
rect 35 46 43 59
rect 35 44 38 46
rect 40 44 43 46
rect 35 42 43 44
rect 45 42 50 70
rect 52 68 60 70
rect 52 66 55 68
rect 57 66 60 68
rect 52 42 60 66
rect 62 42 67 70
rect 69 61 77 70
rect 69 59 72 61
rect 74 59 77 61
rect 69 46 77 59
rect 69 44 72 46
rect 74 44 77 46
rect 69 42 77 44
rect 79 53 87 70
rect 79 51 82 53
rect 84 51 87 53
rect 79 46 87 51
rect 79 44 82 46
rect 84 44 87 46
rect 79 42 87 44
rect 89 61 94 70
rect 112 61 117 70
rect 89 59 97 61
rect 89 57 92 59
rect 94 57 97 59
rect 89 42 97 57
rect 99 53 107 61
rect 99 51 102 53
rect 104 51 107 53
rect 99 46 107 51
rect 99 44 102 46
rect 104 44 107 46
rect 99 42 107 44
rect 109 59 117 61
rect 109 57 112 59
rect 114 57 117 59
rect 109 42 117 57
rect 119 60 127 70
rect 119 58 122 60
rect 124 58 127 60
rect 119 53 127 58
rect 119 51 122 53
rect 124 51 127 53
rect 119 42 127 51
rect 129 68 137 70
rect 129 66 132 68
rect 134 66 137 68
rect 129 61 137 66
rect 129 59 132 61
rect 134 59 137 61
rect 129 42 137 59
rect 139 53 147 70
rect 139 51 142 53
rect 144 51 147 53
rect 139 46 147 51
rect 139 44 142 46
rect 144 44 147 46
rect 139 42 147 44
rect 149 61 154 70
rect 149 59 157 61
rect 149 57 152 59
rect 154 57 157 59
rect 149 42 157 57
rect 159 55 164 61
rect 159 53 166 55
rect 159 51 162 53
rect 164 51 166 53
rect 159 46 166 51
rect 159 44 162 46
rect 164 44 166 46
rect 159 42 166 44
<< alu1 >>
rect -2 81 170 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 170 81
rect -2 68 170 79
rect 17 61 95 62
rect 17 59 38 61
rect 40 59 72 61
rect 74 59 95 61
rect 17 58 92 59
rect 17 54 23 58
rect 91 57 92 58
rect 94 57 95 59
rect 91 55 95 57
rect 2 53 23 54
rect 2 51 4 53
rect 6 51 23 53
rect 2 50 23 51
rect 2 46 7 50
rect 2 44 4 46
rect 6 44 7 46
rect 2 41 7 44
rect 113 42 135 46
rect 113 38 117 42
rect 131 38 135 42
rect 93 37 117 38
rect 93 35 95 37
rect 97 35 117 37
rect 93 34 117 35
rect 121 37 127 38
rect 121 35 123 37
rect 125 35 127 37
rect 121 30 127 35
rect 131 37 139 38
rect 131 35 135 37
rect 137 35 139 37
rect 131 34 139 35
rect 121 26 135 30
rect -2 11 170 12
rect -2 9 82 11
rect 84 9 103 11
rect 105 9 125 11
rect 127 9 170 11
rect -2 1 170 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 170 1
rect -2 -2 170 -1
<< ptie >>
rect 0 1 168 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 168 1
rect 0 -3 168 -1
<< ntie >>
rect 0 81 168 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 168 81
rect 0 77 168 79
<< nmos >>
rect 26 18 28 29
rect 36 18 38 29
rect 46 11 48 29
rect 56 11 58 29
rect 66 13 68 29
rect 76 10 78 29
rect 88 10 90 29
rect 109 11 111 30
rect 119 11 121 30
<< pmos >>
rect 9 42 11 70
rect 16 42 18 70
rect 26 42 28 70
rect 33 42 35 70
rect 43 42 45 70
rect 50 42 52 70
rect 60 42 62 70
rect 67 42 69 70
rect 77 42 79 70
rect 87 42 89 70
rect 97 42 99 61
rect 107 42 109 61
rect 117 42 119 70
rect 127 42 129 70
rect 137 42 139 70
rect 147 42 149 70
rect 157 42 159 61
<< polyct0 >>
rect 7 35 9 37
rect 34 35 36 37
rect 68 35 70 37
rect 13 18 15 20
<< polyct1 >>
rect 95 35 97 37
rect 123 35 125 37
rect 135 35 137 37
<< ndifct0 >>
rect 21 25 23 27
rect 31 20 33 22
rect 41 25 43 27
rect 51 25 53 27
rect 61 25 63 27
rect 71 18 73 20
rect 93 18 95 20
rect 114 26 116 28
<< ndifct1 >>
rect 82 9 84 11
rect 103 9 105 11
rect 125 9 127 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
<< pdifct0 >>
rect 21 66 23 68
rect 38 44 40 46
rect 55 66 57 68
rect 72 44 74 46
rect 82 51 84 53
rect 82 44 84 46
rect 102 51 104 53
rect 102 44 104 46
rect 112 57 114 59
rect 122 58 124 60
rect 122 51 124 53
rect 132 66 134 68
rect 132 59 134 61
rect 142 51 144 53
rect 142 44 144 46
rect 152 57 154 59
rect 162 51 164 53
rect 162 44 164 46
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 38 59 40 61
rect 72 59 74 61
rect 92 57 94 59
<< alu0 >>
rect 19 66 21 68
rect 23 66 25 68
rect 19 65 25 66
rect 53 66 55 68
rect 57 66 59 68
rect 53 65 59 66
rect 110 59 116 68
rect 131 66 132 68
rect 134 66 135 68
rect 110 57 112 59
rect 114 57 116 59
rect 110 56 116 57
rect 121 60 125 62
rect 121 58 122 60
rect 124 58 125 60
rect 28 53 86 54
rect 28 51 82 53
rect 84 51 86 53
rect 28 50 86 51
rect 28 38 32 50
rect 36 46 45 47
rect 36 44 38 46
rect 40 44 45 46
rect 36 43 45 44
rect 5 37 38 38
rect 5 35 7 37
rect 9 35 34 37
rect 36 35 38 37
rect 5 34 38 35
rect 41 30 45 43
rect 19 27 45 30
rect 19 25 21 27
rect 23 26 41 27
rect 23 25 25 26
rect 19 24 25 25
rect 39 25 41 26
rect 43 25 45 27
rect 39 24 45 25
rect 49 28 53 50
rect 59 46 76 47
rect 59 44 72 46
rect 74 44 76 46
rect 59 43 76 44
rect 81 46 86 50
rect 101 53 105 55
rect 121 53 125 58
rect 131 61 135 66
rect 131 59 132 61
rect 134 59 135 61
rect 131 57 135 59
rect 151 59 155 68
rect 151 57 152 59
rect 154 57 155 59
rect 151 55 155 57
rect 101 51 102 53
rect 104 51 122 53
rect 124 51 125 53
rect 101 49 125 51
rect 141 53 145 55
rect 141 51 142 53
rect 144 51 145 53
rect 101 46 105 49
rect 141 46 145 51
rect 161 53 165 55
rect 161 51 162 53
rect 164 51 165 53
rect 161 46 165 51
rect 81 44 82 46
rect 84 44 102 46
rect 104 44 105 46
rect 59 28 63 43
rect 81 42 105 44
rect 141 44 142 46
rect 144 44 162 46
rect 164 44 165 46
rect 141 42 165 44
rect 81 38 85 42
rect 66 37 85 38
rect 66 35 68 37
rect 70 35 85 37
rect 66 34 85 35
rect 81 29 85 34
rect 81 28 118 29
rect 49 27 55 28
rect 49 25 51 27
rect 53 25 55 27
rect 49 24 55 25
rect 59 27 65 28
rect 59 25 61 27
rect 63 25 65 27
rect 81 26 114 28
rect 116 26 118 28
rect 81 25 118 26
rect 59 24 65 25
rect 29 22 35 23
rect 29 21 31 22
rect 11 20 31 21
rect 33 21 35 22
rect 143 21 147 42
rect 33 20 147 21
rect 11 18 13 20
rect 15 18 71 20
rect 73 18 93 20
rect 95 18 147 20
rect 11 17 147 18
<< labels >>
rlabel alu0 21 36 21 36 6 an
rlabel alu0 51 39 51 39 6 an
rlabel alu0 75 36 75 36 6 an
rlabel alu0 83 39 83 39 6 an
rlabel alu0 99 27 99 27 6 an
rlabel alu0 123 55 123 55 6 an
rlabel alu0 103 48 103 48 6 an
rlabel alu0 79 19 79 19 6 bn
rlabel alu0 163 48 163 48 6 bn
rlabel alu0 143 48 143 48 6 bn
rlabel alu1 4 44 4 44 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 60 28 60 6 z
rlabel alu1 36 60 36 60 6 z
rlabel alu1 52 60 52 60 6 z
rlabel alu1 60 60 60 60 6 z
rlabel alu1 68 60 68 60 6 z
rlabel alu1 76 60 76 60 6 z
rlabel alu1 44 60 44 60 6 z
rlabel alu1 84 6 84 6 6 vss
rlabel alu1 108 36 108 36 6 b
rlabel alu1 100 36 100 36 6 b
rlabel alu1 124 32 124 32 6 a
rlabel alu1 116 44 116 44 6 b
rlabel alu1 124 44 124 44 6 b
rlabel alu1 92 60 92 60 6 z
rlabel alu1 84 60 84 60 6 z
rlabel alu1 84 74 84 74 6 vdd
rlabel alu1 132 28 132 28 6 a
rlabel alu1 132 44 132 44 6 b
<< end >>
