magic
tech scmos
timestamp 1199543130
<< ab >>
rect 0 0 90 100
<< nwell >>
rect -5 48 95 105
<< pwell >>
rect -5 -5 95 48
<< poly >>
rect 45 94 47 98
rect 57 94 59 98
rect 67 94 69 98
rect 77 94 79 98
rect 11 85 13 89
rect 23 85 25 89
rect 33 85 35 89
rect 11 43 13 55
rect 23 53 25 56
rect 33 53 35 56
rect 45 53 47 56
rect 21 51 25 53
rect 31 51 35 53
rect 43 51 47 53
rect 57 53 59 56
rect 67 53 69 56
rect 57 51 63 53
rect 21 43 23 51
rect 31 43 33 51
rect 43 43 45 51
rect 57 49 59 51
rect 61 49 63 51
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 37 41 45 43
rect 37 39 39 41
rect 41 39 45 41
rect 37 37 45 39
rect 11 34 13 37
rect 21 34 23 37
rect 31 34 33 37
rect 43 34 45 37
rect 55 47 63 49
rect 67 51 73 53
rect 67 49 69 51
rect 71 49 73 51
rect 67 47 73 49
rect 55 35 57 47
rect 67 39 69 47
rect 65 37 69 39
rect 77 43 79 55
rect 77 41 83 43
rect 77 39 79 41
rect 81 39 83 41
rect 77 37 83 39
rect 65 34 67 37
rect 77 34 79 37
rect 43 12 45 16
rect 55 13 57 17
rect 65 13 67 17
rect 77 13 79 17
rect 11 6 13 10
rect 21 6 23 10
rect 31 6 33 10
<< ndif >>
rect 50 34 55 35
rect 3 11 11 34
rect 3 9 5 11
rect 7 10 11 11
rect 13 10 21 34
rect 23 10 31 34
rect 33 21 43 34
rect 33 19 37 21
rect 39 19 43 21
rect 33 16 43 19
rect 45 21 55 34
rect 45 19 49 21
rect 51 19 55 21
rect 45 17 55 19
rect 57 34 62 35
rect 57 17 65 34
rect 67 21 77 34
rect 67 19 71 21
rect 73 19 77 21
rect 67 17 77 19
rect 79 21 87 34
rect 79 19 83 21
rect 85 19 87 21
rect 79 17 87 19
rect 45 16 52 17
rect 33 10 40 16
rect 59 11 63 17
rect 7 9 9 10
rect 3 7 9 9
rect 58 9 64 11
rect 58 7 60 9
rect 62 7 64 9
rect 58 5 64 7
<< pdif >>
rect 26 95 32 97
rect 26 93 28 95
rect 30 93 32 95
rect 26 91 32 93
rect 27 85 31 91
rect 40 85 45 94
rect 3 81 11 85
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 81 23 85
rect 13 79 17 81
rect 19 79 23 81
rect 13 56 23 79
rect 25 56 33 85
rect 35 81 45 85
rect 35 79 39 81
rect 41 79 45 81
rect 35 56 45 79
rect 47 71 57 94
rect 47 69 51 71
rect 53 69 57 71
rect 47 56 57 69
rect 59 56 67 94
rect 69 56 77 94
rect 13 55 18 56
rect 72 55 77 56
rect 79 81 87 94
rect 79 79 83 81
rect 85 79 87 81
rect 79 55 87 79
<< alu1 >>
rect -2 95 92 100
rect -2 93 8 95
rect 10 93 16 95
rect 18 93 28 95
rect 30 93 92 95
rect -2 88 92 93
rect 4 81 8 88
rect 4 79 5 81
rect 7 79 8 81
rect 4 77 8 79
rect 15 81 87 82
rect 15 79 17 81
rect 19 79 39 81
rect 41 79 83 81
rect 85 79 87 81
rect 15 78 87 79
rect 8 41 12 73
rect 8 39 9 41
rect 11 39 12 41
rect 8 17 12 39
rect 18 41 22 73
rect 18 39 19 41
rect 21 39 22 41
rect 18 17 22 39
rect 28 41 32 73
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 41 42 73
rect 38 39 39 41
rect 41 39 42 41
rect 38 37 42 39
rect 48 72 52 73
rect 48 71 55 72
rect 48 69 51 71
rect 53 69 55 71
rect 48 68 55 69
rect 38 32 42 33
rect 48 32 52 68
rect 38 28 52 32
rect 38 22 42 28
rect 48 27 52 28
rect 58 51 62 63
rect 58 49 59 51
rect 61 49 62 51
rect 58 27 62 49
rect 68 51 72 73
rect 68 49 69 51
rect 71 49 72 51
rect 68 27 72 49
rect 78 41 82 73
rect 78 39 79 41
rect 81 39 82 41
rect 78 27 82 39
rect 35 21 42 22
rect 35 19 37 21
rect 39 19 42 21
rect 35 18 42 19
rect 47 21 75 22
rect 47 19 49 21
rect 51 19 71 21
rect 73 19 75 21
rect 47 18 75 19
rect 82 21 86 23
rect 82 19 83 21
rect 85 19 86 21
rect 38 17 42 18
rect 82 12 86 19
rect -2 11 92 12
rect -2 9 5 11
rect 7 9 92 11
rect -2 7 60 9
rect 62 7 73 9
rect 75 7 81 9
rect 83 7 92 9
rect -2 0 92 7
<< ptie >>
rect 71 9 85 11
rect 71 7 73 9
rect 75 7 81 9
rect 83 7 85 9
rect 71 5 85 7
<< ntie >>
rect 6 95 20 97
rect 6 93 8 95
rect 10 93 16 95
rect 18 93 20 95
rect 6 91 20 93
<< nmos >>
rect 11 10 13 34
rect 21 10 23 34
rect 31 10 33 34
rect 43 16 45 34
rect 55 17 57 35
rect 65 17 67 34
rect 77 17 79 34
<< pmos >>
rect 11 55 13 85
rect 23 56 25 85
rect 33 56 35 85
rect 45 56 47 94
rect 57 56 59 94
rect 67 56 69 94
rect 77 55 79 94
<< polyct1 >>
rect 59 49 61 51
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 39 39 41 41
rect 69 49 71 51
rect 79 39 81 41
<< ndifct1 >>
rect 5 9 7 11
rect 37 19 39 21
rect 49 19 51 21
rect 71 19 73 21
rect 83 19 85 21
rect 60 7 62 9
<< ntiect1 >>
rect 8 93 10 95
rect 16 93 18 95
<< ptiect1 >>
rect 73 7 75 9
rect 81 7 83 9
<< pdifct1 >>
rect 28 93 30 95
rect 5 79 7 81
rect 17 79 19 81
rect 39 79 41 81
rect 51 69 53 71
rect 83 79 85 81
<< labels >>
rlabel alu1 10 45 10 45 6 i0
rlabel alu1 40 25 40 25 6 nq
rlabel alu1 20 45 20 45 6 i1
rlabel alu1 30 50 30 50 6 i2
rlabel alu1 40 55 40 55 6 i6
rlabel alu1 45 6 45 6 6 vss
rlabel alu1 60 45 60 45 6 i3
rlabel alu1 50 50 50 50 6 nq
rlabel alu1 45 94 45 94 6 vdd
rlabel alu1 80 50 80 50 6 i5
rlabel polyct1 70 50 70 50 6 i4
<< end >>
