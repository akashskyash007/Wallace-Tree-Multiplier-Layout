magic
tech scmos
timestamp 1199202412
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 9 61 11 65
rect 9 39 11 43
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 28 11 33
rect 9 15 11 19
<< ndif >>
rect 2 26 9 28
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 4 19 9 22
rect 11 19 20 28
rect 13 11 20 19
rect 13 9 15 11
rect 17 9 20 11
rect 13 7 20 9
<< pdif >>
rect 13 71 20 73
rect 13 69 15 71
rect 17 69 20 71
rect 13 61 20 69
rect 4 56 9 61
rect 2 54 9 56
rect 2 52 4 54
rect 6 52 9 54
rect 2 47 9 52
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 43 20 61
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 71 26 79
rect -2 69 15 71
rect 17 69 26 71
rect -2 68 26 69
rect 2 57 14 63
rect 2 54 6 57
rect 2 52 4 54
rect 2 47 6 52
rect 2 45 4 47
rect 2 26 6 45
rect 18 39 22 63
rect 10 37 22 39
rect 10 35 11 37
rect 13 35 22 37
rect 10 33 22 35
rect 2 24 4 26
rect 2 23 6 24
rect 2 17 14 23
rect 18 17 22 33
rect -2 11 26 12
rect -2 9 15 11
rect 17 9 26 11
rect -2 1 26 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 9 19 11 28
<< pmos >>
rect 9 43 11 61
<< polyct1 >>
rect 11 35 13 37
<< ndifct1 >>
rect 4 24 6 26
rect 15 9 17 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct1 >>
rect 15 69 17 71
rect 4 52 6 54
rect 4 45 6 47
<< alu0 >>
rect 6 43 7 57
rect 6 23 7 28
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 12 60 12 60 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 40 20 40 6 a
<< end >>
