magic
tech scmos
timestamp 1199542834
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 11 43 13 55
rect 23 43 25 55
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 25 43
rect 17 39 19 41
rect 21 39 25 41
rect 17 37 25 39
rect 11 25 13 37
rect 23 25 25 37
rect 35 43 37 55
rect 35 41 43 43
rect 35 39 39 41
rect 41 39 43 41
rect 35 37 43 39
rect 35 25 37 37
rect 11 2 13 6
rect 23 2 25 6
rect 35 2 37 6
<< ndif >>
rect 3 11 11 25
rect 3 9 5 11
rect 7 9 11 11
rect 3 6 11 9
rect 13 6 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 6 35 19
rect 37 11 45 25
rect 37 9 41 11
rect 43 9 45 11
rect 37 6 45 9
<< pdif >>
rect 3 81 11 94
rect 3 79 5 81
rect 7 79 11 81
rect 3 71 11 79
rect 3 69 5 71
rect 7 69 11 71
rect 3 55 11 69
rect 13 71 23 94
rect 13 69 17 71
rect 19 69 23 71
rect 13 55 23 69
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 55 35 79
rect 37 91 45 94
rect 37 89 41 91
rect 43 89 45 91
rect 37 55 45 89
<< alu1 >>
rect -2 95 62 100
rect -2 93 53 95
rect 55 93 62 95
rect -2 91 62 93
rect -2 89 41 91
rect 43 89 62 91
rect -2 88 62 89
rect 4 82 8 83
rect 4 81 33 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 33 81
rect 4 78 33 79
rect 4 71 8 78
rect 28 72 32 73
rect 4 69 5 71
rect 7 69 8 71
rect 4 67 8 69
rect 15 71 32 72
rect 15 69 17 71
rect 19 69 32 71
rect 15 68 32 69
rect 8 41 12 63
rect 8 39 9 41
rect 11 39 12 41
rect 8 17 12 39
rect 18 41 22 63
rect 18 39 19 41
rect 21 39 22 41
rect 18 17 22 39
rect 28 21 32 68
rect 28 19 29 21
rect 31 19 32 21
rect 28 17 32 19
rect 38 41 42 83
rect 52 59 56 88
rect 52 57 53 59
rect 55 57 56 59
rect 52 55 56 57
rect 38 39 39 41
rect 41 39 42 41
rect 38 17 42 39
rect 52 35 56 37
rect 52 33 53 35
rect 55 33 56 35
rect 52 12 56 33
rect -2 11 62 12
rect -2 9 5 11
rect 7 9 41 11
rect 43 9 62 11
rect -2 7 62 9
rect -2 5 53 7
rect 55 5 62 7
rect -2 0 62 5
<< ptie >>
rect 51 35 57 37
rect 51 33 53 35
rect 55 33 57 35
rect 51 26 57 33
rect 51 7 57 14
rect 51 5 53 7
rect 55 5 57 7
rect 51 3 57 5
<< ntie >>
rect 51 95 57 97
rect 51 93 53 95
rect 55 93 57 95
rect 51 86 57 93
rect 51 59 57 66
rect 51 57 53 59
rect 55 57 57 59
rect 51 55 57 57
<< nmos >>
rect 11 6 13 25
rect 23 6 25 25
rect 35 6 37 25
<< pmos >>
rect 11 55 13 94
rect 23 55 25 94
rect 35 55 37 94
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 39 39 41 41
<< ndifct1 >>
rect 5 9 7 11
rect 29 19 31 21
rect 41 9 43 11
<< ntiect1 >>
rect 53 93 55 95
rect 53 57 55 59
<< ptiect1 >>
rect 53 33 55 35
rect 53 5 55 7
<< pdifct1 >>
rect 5 79 7 81
rect 5 69 7 71
rect 17 69 19 71
rect 29 79 31 81
rect 41 89 43 91
<< labels >>
rlabel polyct1 10 40 10 40 6 i0
rlabel polyct1 20 40 20 40 6 i1
rlabel alu1 20 70 20 70 6 nq
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 30 45 30 45 6 nq
rlabel alu1 40 50 40 50 6 i2
rlabel alu1 30 94 30 94 6 vdd
<< end >>
