magic
tech scmos
timestamp 1199202157
<< ab >>
rect 0 0 128 72
<< nwell >>
rect -5 32 133 77
<< pwell >>
rect -5 -5 133 32
<< poly >>
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 71 66 73 70
rect 78 66 80 70
rect 88 66 90 70
rect 95 66 97 70
rect 107 66 109 70
rect 117 66 119 70
rect 9 54 11 59
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 33 21 35
rect 9 31 11 33
rect 13 31 21 33
rect 9 29 21 31
rect 25 33 31 35
rect 25 31 27 33
rect 29 31 31 33
rect 25 29 31 31
rect 9 26 11 29
rect 19 23 21 29
rect 29 26 31 29
rect 39 35 41 38
rect 49 35 51 38
rect 39 33 51 35
rect 39 31 41 33
rect 43 31 51 33
rect 39 29 51 31
rect 39 26 41 29
rect 49 26 51 29
rect 59 35 61 38
rect 71 35 73 38
rect 59 33 73 35
rect 59 31 63 33
rect 65 31 73 33
rect 59 29 73 31
rect 59 26 61 29
rect 71 26 73 29
rect 78 35 80 38
rect 88 35 90 38
rect 78 33 90 35
rect 78 31 86 33
rect 88 31 90 33
rect 78 29 90 31
rect 78 26 80 29
rect 88 26 90 29
rect 95 35 97 38
rect 107 35 109 38
rect 117 35 119 38
rect 95 33 103 35
rect 95 31 99 33
rect 101 31 103 33
rect 95 29 103 31
rect 107 33 119 35
rect 107 31 115 33
rect 117 31 119 33
rect 107 29 119 31
rect 95 26 97 29
rect 107 26 109 29
rect 117 26 119 29
rect 9 11 11 15
rect 19 7 21 12
rect 29 7 31 12
rect 39 7 41 12
rect 49 7 51 12
rect 59 7 61 12
rect 88 11 90 15
rect 95 11 97 15
rect 71 4 73 9
rect 78 4 80 9
rect 107 7 109 12
rect 117 7 119 12
<< ndif >>
rect 2 19 9 26
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 23 16 26
rect 23 23 29 26
rect 11 21 19 23
rect 11 19 14 21
rect 16 19 19 21
rect 11 15 19 19
rect 14 12 19 15
rect 21 16 29 23
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 31 16 39 26
rect 31 14 34 16
rect 36 14 39 16
rect 31 12 39 14
rect 41 24 49 26
rect 41 22 44 24
rect 46 22 49 24
rect 41 12 49 22
rect 51 16 59 26
rect 51 14 54 16
rect 56 14 59 16
rect 51 12 59 14
rect 61 12 71 26
rect 63 9 71 12
rect 73 9 78 26
rect 80 24 88 26
rect 80 22 83 24
rect 85 22 88 24
rect 80 15 88 22
rect 90 15 95 26
rect 97 15 107 26
rect 80 9 85 15
rect 99 12 107 15
rect 109 16 117 26
rect 109 14 112 16
rect 114 14 117 16
rect 109 12 117 14
rect 119 23 126 26
rect 119 21 122 23
rect 124 21 126 23
rect 119 16 126 21
rect 119 14 122 16
rect 124 14 126 16
rect 119 12 126 14
rect 63 7 69 9
rect 63 5 65 7
rect 67 5 69 7
rect 63 3 69 5
rect 99 7 105 12
rect 99 5 101 7
rect 103 5 105 7
rect 99 3 105 5
<< pdif >>
rect 14 54 19 66
rect 2 52 9 54
rect 2 50 4 52
rect 6 50 9 52
rect 2 38 9 50
rect 11 49 19 54
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 57 39 66
rect 31 55 34 57
rect 36 55 39 57
rect 31 38 39 55
rect 41 42 49 66
rect 41 40 44 42
rect 46 40 49 42
rect 41 38 49 40
rect 51 57 59 66
rect 51 55 54 57
rect 56 55 59 57
rect 51 38 59 55
rect 61 64 71 66
rect 61 62 65 64
rect 67 62 71 64
rect 61 38 71 62
rect 73 38 78 66
rect 80 42 88 66
rect 80 40 83 42
rect 85 40 88 42
rect 80 38 88 40
rect 90 38 95 66
rect 97 64 107 66
rect 97 62 101 64
rect 103 62 107 64
rect 97 38 107 62
rect 109 57 117 66
rect 109 55 112 57
rect 114 55 117 57
rect 109 50 117 55
rect 109 48 112 50
rect 114 48 117 50
rect 109 38 117 48
rect 119 64 126 66
rect 119 62 122 64
rect 124 62 126 64
rect 119 56 126 62
rect 119 54 122 56
rect 124 54 126 56
rect 119 38 126 54
<< alu1 >>
rect -2 67 130 72
rect -2 65 5 67
rect 7 65 130 67
rect -2 64 130 65
rect 2 35 6 43
rect 26 46 103 50
rect 2 33 14 35
rect 2 31 11 33
rect 13 31 14 33
rect 2 29 14 31
rect 26 33 30 46
rect 41 40 44 42
rect 46 40 55 42
rect 41 38 55 40
rect 26 31 27 33
rect 29 31 30 33
rect 26 29 30 31
rect 50 26 55 38
rect 73 40 83 42
rect 85 40 87 42
rect 73 38 87 40
rect 97 38 103 46
rect 73 26 78 38
rect 84 33 95 34
rect 84 31 86 33
rect 88 31 95 33
rect 84 30 95 31
rect 89 26 95 30
rect 114 33 118 35
rect 114 31 115 33
rect 117 31 118 33
rect 114 26 118 31
rect 41 24 78 26
rect 41 22 44 24
rect 46 22 78 24
rect 89 22 118 26
rect -2 7 130 8
rect -2 5 5 7
rect 7 5 65 7
rect 67 5 91 7
rect 93 5 101 7
rect 103 5 130 7
rect -2 0 130 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
rect 89 7 95 9
rect 89 5 91 7
rect 93 5 95 7
rect 89 3 95 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 15 11 26
rect 19 12 21 23
rect 29 12 31 26
rect 39 12 41 26
rect 49 12 51 26
rect 59 12 61 26
rect 71 9 73 26
rect 78 9 80 26
rect 88 15 90 26
rect 95 15 97 26
rect 107 12 109 26
rect 117 12 119 26
<< pmos >>
rect 9 38 11 54
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 66
rect 59 38 61 66
rect 71 38 73 66
rect 78 38 80 66
rect 88 38 90 66
rect 95 38 97 66
rect 107 38 109 66
rect 117 38 119 66
<< polyct0 >>
rect 41 31 43 33
rect 63 31 65 33
rect 99 31 101 33
<< polyct1 >>
rect 11 31 13 33
rect 27 31 29 33
rect 86 31 88 33
rect 115 31 117 33
<< ndifct0 >>
rect 4 17 6 19
rect 14 19 16 21
rect 24 14 26 16
rect 34 14 36 16
rect 54 14 56 16
rect 83 22 85 24
rect 112 14 114 16
rect 122 21 124 23
rect 122 14 124 16
<< ndifct1 >>
rect 44 22 46 24
rect 65 5 67 7
rect 101 5 103 7
<< ntiect1 >>
rect 5 65 7 67
<< ptiect1 >>
rect 5 5 7 7
rect 91 5 93 7
<< pdifct0 >>
rect 4 50 6 52
rect 14 47 16 49
rect 14 40 16 42
rect 24 62 26 64
rect 24 55 26 57
rect 34 55 36 57
rect 54 55 56 57
rect 65 62 67 64
rect 101 62 103 64
rect 112 55 114 57
rect 112 48 114 50
rect 122 62 124 64
rect 122 54 124 56
<< pdifct1 >>
rect 44 40 46 42
rect 83 40 85 42
<< alu0 >>
rect 3 52 7 64
rect 23 62 24 64
rect 26 62 27 64
rect 23 57 27 62
rect 63 62 65 64
rect 67 62 69 64
rect 63 61 69 62
rect 99 62 101 64
rect 103 62 105 64
rect 99 61 105 62
rect 121 62 122 64
rect 124 62 125 64
rect 23 55 24 57
rect 26 55 27 57
rect 23 53 27 55
rect 32 57 116 58
rect 32 55 34 57
rect 36 55 54 57
rect 56 55 112 57
rect 114 55 116 57
rect 32 54 116 55
rect 3 50 4 52
rect 6 50 7 52
rect 3 48 7 50
rect 13 49 17 51
rect 111 50 116 54
rect 121 56 125 62
rect 121 54 122 56
rect 124 54 125 56
rect 121 52 125 54
rect 13 47 14 49
rect 16 47 17 49
rect 13 42 17 47
rect 111 48 112 50
rect 114 48 116 50
rect 111 46 116 48
rect 13 40 14 42
rect 16 40 22 42
rect 13 38 22 40
rect 18 25 22 38
rect 42 42 48 43
rect 34 33 45 34
rect 34 31 41 33
rect 43 31 45 33
rect 34 30 45 31
rect 34 25 38 30
rect 62 33 66 46
rect 81 42 87 43
rect 62 31 63 33
rect 65 31 66 33
rect 62 29 66 31
rect 98 33 102 38
rect 98 31 99 33
rect 101 31 102 33
rect 98 29 102 31
rect 13 21 38 25
rect 78 24 86 26
rect 78 22 83 24
rect 85 22 86 24
rect 121 23 125 25
rect 42 21 48 22
rect 3 19 7 21
rect 3 17 4 19
rect 6 17 7 19
rect 13 19 14 21
rect 16 19 17 21
rect 73 20 86 22
rect 121 21 122 23
rect 124 21 125 23
rect 13 17 17 19
rect 3 8 7 17
rect 23 16 27 18
rect 23 14 24 16
rect 26 14 27 16
rect 23 8 27 14
rect 32 16 116 17
rect 32 14 34 16
rect 36 14 54 16
rect 56 14 112 16
rect 114 14 116 16
rect 32 13 116 14
rect 121 16 125 21
rect 121 14 122 16
rect 124 14 125 16
rect 121 8 125 14
<< labels >>
rlabel alu0 15 44 15 44 6 cn
rlabel alu0 39 32 39 32 6 cn
rlabel alu0 25 23 25 23 6 cn
rlabel alu0 74 15 74 15 6 n3
rlabel alu0 113 52 113 52 6 n1
rlabel alu0 74 56 74 56 6 n1
rlabel polyct1 12 32 12 32 6 c
rlabel alu1 4 36 4 36 6 c
rlabel alu1 44 24 44 24 6 z
rlabel alu1 44 40 44 40 6 z
rlabel alu1 28 36 28 36 6 a
rlabel alu1 36 48 36 48 6 a
rlabel alu1 44 48 44 48 6 a
rlabel alu1 64 4 64 4 6 vss
rlabel alu1 60 24 60 24 6 z
rlabel alu1 68 24 68 24 6 z
rlabel alu1 52 32 52 32 6 z
rlabel alu1 52 48 52 48 6 a
rlabel alu1 60 48 60 48 6 a
rlabel alu1 68 48 68 48 6 a
rlabel alu1 64 68 64 68 6 vdd
rlabel alu1 100 24 100 24 6 b
rlabel alu1 92 28 92 28 6 b
rlabel alu1 76 32 76 32 6 z
rlabel alu1 84 40 84 40 6 z
rlabel alu1 100 44 100 44 6 a
rlabel alu1 76 48 76 48 6 a
rlabel alu1 84 48 84 48 6 a
rlabel alu1 92 48 92 48 6 a
rlabel alu1 108 24 108 24 6 b
rlabel polyct1 116 32 116 32 6 b
<< end >>
