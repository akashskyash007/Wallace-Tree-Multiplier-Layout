magic
tech scmos
timestamp 1199203702
<< ab >>
rect 0 0 120 80
<< nwell >>
rect -5 36 125 88
<< pwell >>
rect -5 -8 125 36
<< poly >>
rect 17 67 19 72
rect 29 67 31 72
rect 39 67 41 72
rect 49 67 51 72
rect 77 70 79 74
rect 2 53 8 55
rect 2 51 4 53
rect 6 51 8 53
rect 2 49 8 51
rect 6 45 8 49
rect 89 65 91 70
rect 99 65 101 70
rect 109 65 111 70
rect 77 51 79 54
rect 65 49 79 51
rect 17 45 19 48
rect 6 43 19 45
rect 9 25 11 43
rect 29 38 31 48
rect 39 39 41 48
rect 49 45 51 48
rect 65 47 67 49
rect 69 47 71 49
rect 65 45 71 47
rect 45 43 51 45
rect 45 41 47 43
rect 49 41 51 43
rect 89 41 91 49
rect 45 39 51 41
rect 55 39 91 41
rect 99 40 101 49
rect 17 36 31 38
rect 35 37 41 39
rect 17 34 19 36
rect 21 34 23 36
rect 17 32 23 34
rect 35 35 37 37
rect 39 35 41 37
rect 35 33 41 35
rect 20 25 22 32
rect 39 31 41 33
rect 30 25 32 29
rect 39 28 42 31
rect 40 25 42 28
rect 47 25 49 39
rect 55 37 57 39
rect 59 37 61 39
rect 55 35 61 37
rect 65 33 71 35
rect 65 31 67 33
rect 69 31 71 33
rect 65 29 71 31
rect 69 26 71 29
rect 81 23 83 39
rect 95 38 101 40
rect 109 39 111 49
rect 95 36 97 38
rect 99 36 101 38
rect 95 34 101 36
rect 99 29 101 34
rect 105 37 111 39
rect 105 35 107 37
rect 109 35 111 37
rect 105 33 111 35
rect 91 23 93 28
rect 99 26 103 29
rect 101 23 103 26
rect 108 23 110 33
rect 9 8 11 16
rect 20 12 22 16
rect 30 8 32 16
rect 40 11 42 16
rect 47 11 49 16
rect 9 6 32 8
rect 69 8 71 19
rect 81 12 83 16
rect 91 8 93 16
rect 101 11 103 16
rect 108 11 110 16
rect 69 6 93 8
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 4 16 9 19
rect 11 20 20 25
rect 11 18 15 20
rect 17 18 20 20
rect 11 16 20 18
rect 22 20 30 25
rect 22 18 25 20
rect 27 18 30 20
rect 22 16 30 18
rect 32 21 40 25
rect 32 19 35 21
rect 37 19 40 21
rect 32 16 40 19
rect 42 16 47 25
rect 49 16 57 25
rect 62 24 69 26
rect 62 22 64 24
rect 66 22 69 24
rect 62 19 69 22
rect 71 23 79 26
rect 71 19 81 23
rect 51 14 57 16
rect 51 12 53 14
rect 55 12 57 14
rect 51 10 57 12
rect 73 16 81 19
rect 83 21 91 23
rect 83 19 86 21
rect 88 19 91 21
rect 83 16 91 19
rect 93 21 101 23
rect 93 19 96 21
rect 98 19 101 21
rect 93 16 101 19
rect 103 16 108 23
rect 110 16 118 23
rect 73 14 75 16
rect 77 14 79 16
rect 73 12 79 14
rect 112 11 118 16
rect 112 9 114 11
rect 116 9 118 11
rect 112 7 118 9
<< pdif >>
rect 21 71 27 73
rect 21 69 23 71
rect 25 69 27 71
rect 21 67 27 69
rect 81 71 87 73
rect 81 70 83 71
rect 12 54 17 67
rect 10 52 17 54
rect 10 50 12 52
rect 14 50 17 52
rect 10 48 17 50
rect 19 48 29 67
rect 31 52 39 67
rect 31 50 34 52
rect 36 50 39 52
rect 31 48 39 50
rect 41 53 49 67
rect 41 51 44 53
rect 46 51 49 53
rect 41 48 49 51
rect 51 63 56 67
rect 72 64 77 70
rect 51 61 58 63
rect 51 59 54 61
rect 56 59 58 61
rect 51 57 58 59
rect 70 62 77 64
rect 70 60 72 62
rect 74 60 77 62
rect 70 58 77 60
rect 51 48 56 57
rect 72 54 77 58
rect 79 69 83 70
rect 85 69 87 71
rect 79 65 87 69
rect 79 54 89 65
rect 81 49 89 54
rect 91 53 99 65
rect 91 51 94 53
rect 96 51 99 53
rect 91 49 99 51
rect 101 54 109 65
rect 101 52 104 54
rect 106 52 109 54
rect 101 49 109 52
rect 111 62 118 65
rect 111 60 114 62
rect 116 60 118 62
rect 111 58 118 60
rect 111 49 116 58
<< alu1 >>
rect -2 81 122 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 122 81
rect -2 71 122 79
rect -2 69 23 71
rect 25 69 83 71
rect 85 69 122 71
rect -2 68 122 69
rect 2 58 15 63
rect 2 53 7 58
rect 2 51 4 53
rect 6 51 7 53
rect 2 49 7 51
rect 18 36 22 39
rect 18 34 19 36
rect 21 34 22 36
rect 18 31 22 34
rect 10 25 22 31
rect 66 49 70 55
rect 66 47 67 49
rect 69 47 70 49
rect 66 46 70 47
rect 66 42 79 46
rect 66 33 70 42
rect 102 54 118 55
rect 102 52 104 54
rect 106 52 118 54
rect 102 51 118 52
rect 66 31 67 33
rect 69 31 70 33
rect 66 29 70 31
rect 114 22 118 51
rect 94 21 118 22
rect 94 19 96 21
rect 98 19 118 21
rect 94 18 118 19
rect -2 11 122 12
rect -2 9 114 11
rect 116 9 122 11
rect -2 1 122 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 122 1
rect -2 -2 122 -1
<< ptie >>
rect 0 1 120 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 120 1
rect 0 -3 120 -1
<< ntie >>
rect 0 81 120 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 120 81
rect 0 77 120 79
<< nmos >>
rect 9 16 11 25
rect 20 16 22 25
rect 30 16 32 25
rect 40 16 42 25
rect 47 16 49 25
rect 69 19 71 26
rect 81 16 83 23
rect 91 16 93 23
rect 101 16 103 23
rect 108 16 110 23
<< pmos >>
rect 17 48 19 67
rect 29 48 31 67
rect 39 48 41 67
rect 49 48 51 67
rect 77 54 79 70
rect 89 49 91 65
rect 99 49 101 65
rect 109 49 111 65
<< polyct0 >>
rect 47 41 49 43
rect 37 35 39 37
rect 57 37 59 39
rect 97 36 99 38
rect 107 35 109 37
<< polyct1 >>
rect 4 51 6 53
rect 67 47 69 49
rect 19 34 21 36
rect 67 31 69 33
<< ndifct0 >>
rect 4 21 6 23
rect 15 18 17 20
rect 25 18 27 20
rect 35 19 37 21
rect 64 22 66 24
rect 53 12 55 14
rect 86 19 88 21
rect 75 14 77 16
<< ndifct1 >>
rect 96 19 98 21
rect 114 9 116 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
<< pdifct0 >>
rect 12 50 14 52
rect 34 50 36 52
rect 44 51 46 53
rect 54 59 56 61
rect 72 60 74 62
rect 94 51 96 53
rect 114 60 116 62
<< pdifct1 >>
rect 23 69 25 71
rect 83 69 85 71
rect 104 52 106 54
<< alu0 >>
rect 70 62 118 63
rect 26 61 58 62
rect 26 59 54 61
rect 56 59 58 61
rect 70 60 72 62
rect 74 60 114 62
rect 116 60 118 62
rect 70 59 118 60
rect 26 58 58 59
rect 26 54 30 58
rect 11 52 30 54
rect 11 50 12 52
rect 14 50 30 52
rect 11 43 15 50
rect 3 39 15 43
rect 3 23 7 39
rect 26 38 30 50
rect 33 52 37 54
rect 33 50 34 52
rect 36 50 37 52
rect 42 53 58 54
rect 42 51 44 53
rect 46 51 58 53
rect 42 50 58 51
rect 33 46 37 50
rect 33 43 50 46
rect 33 42 47 43
rect 46 41 47 42
rect 49 41 50 43
rect 26 37 41 38
rect 26 35 37 37
rect 39 35 41 37
rect 26 34 41 35
rect 46 30 50 41
rect 26 26 50 30
rect 54 40 58 50
rect 54 39 61 40
rect 54 37 57 39
rect 59 37 61 39
rect 54 36 61 37
rect 3 21 4 23
rect 6 21 7 23
rect 26 21 30 26
rect 54 22 58 36
rect 84 39 88 59
rect 93 53 97 55
rect 93 51 94 53
rect 96 51 97 53
rect 93 47 97 51
rect 93 43 110 47
rect 76 38 101 39
rect 76 36 97 38
rect 99 36 101 38
rect 76 35 101 36
rect 106 37 110 43
rect 106 35 107 37
rect 109 35 110 37
rect 76 25 80 35
rect 106 31 110 35
rect 3 19 7 21
rect 13 20 19 21
rect 13 18 15 20
rect 17 18 19 20
rect 13 12 19 18
rect 23 20 30 21
rect 23 18 25 20
rect 27 18 30 20
rect 33 21 58 22
rect 62 24 80 25
rect 62 22 64 24
rect 66 22 80 24
rect 62 21 80 22
rect 85 27 110 31
rect 85 21 89 27
rect 33 19 35 21
rect 37 19 58 21
rect 33 18 58 19
rect 85 19 86 21
rect 88 19 89 21
rect 23 17 30 18
rect 85 17 89 19
rect 73 16 79 17
rect 51 14 57 15
rect 51 12 53 14
rect 55 12 57 14
rect 73 14 75 16
rect 77 14 79 16
rect 73 12 79 14
<< labels >>
rlabel alu0 5 31 5 31 6 bn
rlabel alu0 13 46 13 46 6 bn
rlabel ndifct0 26 19 26 19 6 an
rlabel alu0 33 36 33 36 6 bn
rlabel alu0 35 48 35 48 6 an
rlabel alu0 45 20 45 20 6 iz
rlabel alu0 48 36 48 36 6 an
rlabel alu0 50 52 50 52 6 iz
rlabel alu0 56 36 56 36 6 iz
rlabel alu0 42 60 42 60 6 bn
rlabel alu0 71 23 71 23 6 cn
rlabel alu0 87 24 87 24 6 zn
rlabel alu0 108 37 108 37 6 zn
rlabel alu0 88 37 88 37 6 cn
rlabel alu0 95 49 95 49 6 zn
rlabel alu0 94 61 94 61 6 cn
rlabel alu1 12 28 12 28 6 a
rlabel alu1 20 32 20 32 6 a
rlabel alu1 4 56 4 56 6 b
rlabel alu1 12 60 12 60 6 b
rlabel alu1 60 6 60 6 6 vss
rlabel alu1 68 44 68 44 6 c
rlabel alu1 76 44 76 44 6 c
rlabel alu1 60 74 60 74 6 vdd
rlabel alu1 100 20 100 20 6 z
rlabel alu1 108 20 108 20 6 z
rlabel alu1 116 40 116 40 6 z
<< end >>
