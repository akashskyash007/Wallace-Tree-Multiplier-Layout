magic
tech scmos
timestamp 1199543546
<< ab >>
rect 0 0 130 100
<< nwell >>
rect -5 48 135 105
<< pwell >>
rect -5 -5 135 48
<< poly >>
rect 11 94 13 98
rect 23 94 25 98
rect 35 94 37 98
rect 47 94 49 98
rect 79 94 81 98
rect 91 94 93 98
rect 103 94 105 98
rect 115 94 117 98
rect 11 53 13 56
rect 23 53 25 56
rect 35 53 37 56
rect 47 53 49 56
rect 79 53 81 56
rect 91 53 93 56
rect 11 51 19 53
rect 23 51 29 53
rect 35 51 43 53
rect 17 43 19 51
rect 27 43 29 51
rect 37 49 39 51
rect 41 49 43 51
rect 37 47 43 49
rect 47 51 53 53
rect 47 49 49 51
rect 51 49 53 51
rect 47 47 53 49
rect 77 51 83 53
rect 77 49 79 51
rect 81 49 83 51
rect 77 47 83 49
rect 87 51 93 53
rect 87 49 89 51
rect 91 49 93 51
rect 87 47 93 49
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 27 37 33 39
rect 17 29 19 37
rect 27 29 29 37
rect 37 29 39 47
rect 47 29 49 47
rect 15 27 19 29
rect 23 27 29 29
rect 35 27 39 29
rect 43 27 49 29
rect 79 29 81 47
rect 79 27 85 29
rect 15 24 17 27
rect 23 24 25 27
rect 35 24 37 27
rect 43 24 45 27
rect 83 24 85 27
rect 91 24 93 47
rect 103 43 105 55
rect 97 41 105 43
rect 115 41 117 55
rect 97 39 99 41
rect 101 39 117 41
rect 97 37 105 39
rect 103 25 105 37
rect 115 25 117 39
rect 15 2 17 6
rect 23 2 25 6
rect 35 2 37 6
rect 43 2 45 6
rect 83 2 85 6
rect 91 2 93 6
rect 103 2 105 6
rect 115 2 117 6
<< ndif >>
rect 98 24 103 25
rect 7 11 15 24
rect 7 9 9 11
rect 11 9 15 11
rect 7 6 15 9
rect 17 6 23 24
rect 25 21 35 24
rect 25 19 29 21
rect 31 19 35 21
rect 25 6 35 19
rect 37 6 43 24
rect 45 11 53 24
rect 75 21 83 24
rect 75 19 77 21
rect 79 19 83 21
rect 45 9 49 11
rect 51 9 53 11
rect 45 6 53 9
rect 75 6 83 19
rect 85 6 91 24
rect 93 11 103 24
rect 93 9 97 11
rect 99 9 103 11
rect 93 6 103 9
rect 105 21 115 25
rect 105 19 109 21
rect 111 19 115 21
rect 105 6 115 19
rect 117 21 125 25
rect 117 19 121 21
rect 123 19 125 21
rect 117 11 125 19
rect 117 9 121 11
rect 123 9 125 11
rect 117 6 125 9
<< pdif >>
rect 3 81 11 94
rect 3 79 5 81
rect 7 79 11 81
rect 3 56 11 79
rect 13 71 23 94
rect 13 69 17 71
rect 19 69 23 71
rect 13 56 23 69
rect 25 81 35 94
rect 25 79 29 81
rect 31 79 35 81
rect 25 56 35 79
rect 37 71 47 94
rect 37 69 41 71
rect 43 69 47 71
rect 37 56 47 69
rect 49 81 57 94
rect 49 79 53 81
rect 55 79 57 81
rect 49 56 57 79
rect 71 91 79 94
rect 71 89 73 91
rect 75 89 79 91
rect 71 81 79 89
rect 71 79 73 81
rect 75 79 79 81
rect 71 56 79 79
rect 81 81 91 94
rect 81 79 85 81
rect 87 79 91 81
rect 81 56 91 79
rect 93 91 103 94
rect 93 89 97 91
rect 99 89 103 91
rect 93 81 103 89
rect 93 79 97 81
rect 99 79 103 81
rect 93 71 103 79
rect 93 69 97 71
rect 99 69 103 71
rect 93 56 103 69
rect 98 55 103 56
rect 105 81 115 94
rect 105 79 109 81
rect 111 79 115 81
rect 105 71 115 79
rect 105 69 109 71
rect 111 69 115 71
rect 105 61 115 69
rect 105 59 109 61
rect 111 59 115 61
rect 105 55 115 59
rect 117 91 125 94
rect 117 89 121 91
rect 123 89 125 91
rect 117 81 125 89
rect 117 79 121 81
rect 123 79 125 81
rect 117 71 125 79
rect 117 69 121 71
rect 123 69 125 71
rect 117 55 125 69
<< alu1 >>
rect -2 91 132 100
rect -2 89 73 91
rect 75 89 97 91
rect 99 89 121 91
rect 123 89 132 91
rect -2 88 132 89
rect 3 81 57 82
rect 3 79 5 81
rect 7 79 29 81
rect 31 79 53 81
rect 55 79 57 81
rect 3 78 57 79
rect 72 81 76 88
rect 72 79 73 81
rect 75 79 76 81
rect 72 77 76 79
rect 84 81 88 83
rect 84 79 85 81
rect 87 79 88 81
rect 15 71 21 72
rect 8 69 17 71
rect 19 69 21 71
rect 8 68 21 69
rect 8 67 20 68
rect 8 22 12 67
rect 18 41 22 63
rect 18 39 19 41
rect 21 39 22 41
rect 18 27 22 39
rect 28 41 32 73
rect 84 72 88 79
rect 39 71 88 72
rect 39 69 41 71
rect 43 69 88 71
rect 39 68 88 69
rect 96 81 100 88
rect 96 79 97 81
rect 99 79 100 81
rect 96 71 100 79
rect 96 69 97 71
rect 99 69 100 71
rect 96 67 100 69
rect 108 81 112 83
rect 108 79 109 81
rect 111 79 112 81
rect 108 71 112 79
rect 108 69 109 71
rect 111 69 112 71
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 51 42 63
rect 38 49 39 51
rect 41 49 42 51
rect 38 27 42 49
rect 48 51 52 63
rect 48 49 49 51
rect 51 49 52 51
rect 48 27 52 49
rect 78 51 82 63
rect 78 49 79 51
rect 81 49 82 51
rect 78 27 82 49
rect 88 51 92 63
rect 88 49 89 51
rect 91 49 92 51
rect 88 27 92 49
rect 108 61 112 69
rect 120 81 124 88
rect 120 79 121 81
rect 123 79 124 81
rect 120 71 124 79
rect 120 69 121 71
rect 123 69 124 71
rect 120 67 124 69
rect 108 59 109 61
rect 111 59 112 61
rect 98 41 102 43
rect 98 39 99 41
rect 101 39 102 41
rect 98 22 102 39
rect 8 21 102 22
rect 8 19 29 21
rect 31 19 77 21
rect 79 19 102 21
rect 8 18 102 19
rect 108 21 112 59
rect 108 19 109 21
rect 111 19 112 21
rect 108 17 112 19
rect 120 21 124 23
rect 120 19 121 21
rect 123 19 124 21
rect 120 12 124 19
rect -2 11 132 12
rect -2 9 9 11
rect 11 9 49 11
rect 51 9 97 11
rect 99 9 121 11
rect 123 9 132 11
rect -2 7 63 9
rect 65 7 132 9
rect -2 0 132 7
<< ptie >>
rect 61 9 67 16
rect 61 7 63 9
rect 65 7 67 9
rect 61 5 67 7
<< nmos >>
rect 15 6 17 24
rect 23 6 25 24
rect 35 6 37 24
rect 43 6 45 24
rect 83 6 85 24
rect 91 6 93 24
rect 103 6 105 25
rect 115 6 117 25
<< pmos >>
rect 11 56 13 94
rect 23 56 25 94
rect 35 56 37 94
rect 47 56 49 94
rect 79 56 81 94
rect 91 56 93 94
rect 103 55 105 94
rect 115 55 117 94
<< polyct1 >>
rect 39 49 41 51
rect 49 49 51 51
rect 79 49 81 51
rect 89 49 91 51
rect 19 39 21 41
rect 29 39 31 41
rect 99 39 101 41
<< ndifct1 >>
rect 9 9 11 11
rect 29 19 31 21
rect 77 19 79 21
rect 49 9 51 11
rect 97 9 99 11
rect 109 19 111 21
rect 121 19 123 21
rect 121 9 123 11
<< ptiect1 >>
rect 63 7 65 9
<< pdifct1 >>
rect 5 79 7 81
rect 17 69 19 71
rect 29 79 31 81
rect 41 69 43 71
rect 53 79 55 81
rect 73 89 75 91
rect 73 79 75 81
rect 85 79 87 81
rect 97 89 99 91
rect 97 79 99 81
rect 97 69 99 71
rect 109 79 111 81
rect 109 69 111 71
rect 109 59 111 61
rect 121 89 123 91
rect 121 79 123 81
rect 121 69 123 71
<< labels >>
rlabel alu1 20 45 20 45 6 i5
rlabel alu1 40 45 40 45 6 i3
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 30 50 30 50 6 i4
rlabel alu1 65 6 65 6 6 vss
rlabel alu1 90 45 90 45 6 i0
rlabel alu1 80 45 80 45 6 i1
rlabel alu1 65 94 65 94 6 vdd
rlabel alu1 110 50 110 50 6 q
<< end >>
