magic
tech scmos
timestamp 1199202352
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 19 68 21 73
rect 29 68 31 73
rect 9 58 11 63
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 9 37 31 39
rect 9 35 17 37
rect 19 35 21 37
rect 9 33 21 35
rect 9 30 11 33
rect 9 8 11 13
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 4 13 9 17
rect 11 25 19 30
rect 11 23 14 25
rect 16 23 19 25
rect 11 17 19 23
rect 11 15 14 17
rect 16 15 19 17
rect 11 13 19 15
<< pdif >>
rect 13 58 19 68
rect 4 55 9 58
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 56 19 58
rect 11 54 14 56
rect 16 54 19 56
rect 11 42 19 54
rect 21 53 29 68
rect 21 51 24 53
rect 26 51 29 53
rect 21 46 29 51
rect 21 44 24 46
rect 26 44 29 46
rect 21 42 29 44
rect 31 66 38 68
rect 31 64 34 66
rect 36 64 38 66
rect 31 58 38 64
rect 31 56 34 58
rect 36 56 38 58
rect 31 42 38 56
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 24 46
rect 26 44 31 46
rect 2 42 31 44
rect 2 30 6 42
rect 15 37 31 38
rect 15 35 17 37
rect 19 35 31 37
rect 15 34 31 35
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect 25 26 31 34
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 9 13 11 30
<< pmos >>
rect 9 42 11 58
rect 19 42 21 68
rect 29 42 31 68
<< polyct1 >>
rect 17 35 19 37
<< ndifct0 >>
rect 14 23 16 25
rect 14 15 16 17
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 54 16 56
rect 24 51 26 53
rect 34 64 36 66
rect 34 56 36 58
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
rect 24 44 26 46
<< alu0 >>
rect 13 56 17 68
rect 13 54 14 56
rect 16 54 17 56
rect 33 66 37 68
rect 33 64 34 66
rect 36 64 37 66
rect 33 58 37 64
rect 33 56 34 58
rect 36 56 37 58
rect 13 52 17 54
rect 23 53 27 55
rect 33 54 37 56
rect 23 51 24 53
rect 26 51 27 53
rect 23 46 27 51
rect 13 25 17 27
rect 13 23 14 25
rect 16 23 17 25
rect 13 17 17 23
rect 13 15 14 17
rect 16 15 17 17
rect 13 12 17 15
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 44 12 44 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 36 20 36 6 a
rlabel alu1 28 32 28 32 6 a
rlabel alu1 28 44 28 44 6 z
rlabel alu1 20 44 20 44 6 z
rlabel alu1 20 74 20 74 6 vdd
<< end >>
