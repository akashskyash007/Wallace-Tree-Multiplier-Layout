magic
tech scmos
timestamp 1199621495
<< ab >>
rect -11 0 307 88
<< alu1 >>
rect -10 69 -6 90
rect -10 67 -9 69
rect -7 67 -6 69
rect -10 53 -6 67
rect -10 51 -9 53
rect -7 51 -6 53
rect -10 37 -6 51
rect -10 35 -9 37
rect -7 35 -6 37
rect -10 21 -6 35
rect -10 19 -9 21
rect -7 19 -6 21
rect -10 2 -6 19
rect -10 -2 306 2
<< alu2 >>
rect -11 69 307 70
rect -11 67 -9 69
rect -7 67 307 69
rect -11 66 307 67
rect -11 53 307 54
rect -11 51 -9 53
rect -7 51 307 53
rect -11 50 307 51
rect -11 37 307 38
rect -11 35 -9 37
rect -7 35 307 37
rect -11 34 307 35
rect -11 21 307 22
rect -11 19 -9 21
rect -7 19 7 21
rect 9 19 23 21
rect 25 19 39 21
rect 41 19 55 21
rect 57 19 71 21
rect 73 19 87 21
rect 89 19 103 21
rect 105 19 119 21
rect 121 19 135 21
rect 137 19 151 21
rect 153 19 167 21
rect 169 19 183 21
rect 185 19 199 21
rect 201 19 215 21
rect 217 19 231 21
rect 233 19 247 21
rect 249 19 263 21
rect 265 19 279 21
rect 281 19 295 21
rect 297 19 307 21
rect -11 18 307 19
<< alu3 >>
rect 6 77 10 90
rect 6 75 7 77
rect 9 75 10 77
rect 6 61 10 75
rect 6 59 7 61
rect 9 59 10 61
rect 6 45 10 59
rect 6 43 7 45
rect 9 43 10 45
rect 6 29 10 43
rect 6 27 7 29
rect 9 27 10 29
rect 6 21 10 27
rect 6 19 7 21
rect 9 19 10 21
rect 6 13 10 19
rect 6 11 7 13
rect 9 11 10 13
rect 6 -2 10 11
rect 22 21 26 90
rect 22 19 23 21
rect 25 19 26 21
rect 22 -2 26 19
rect 38 21 42 90
rect 38 19 39 21
rect 41 19 42 21
rect 38 -2 42 19
rect 54 21 58 90
rect 54 19 55 21
rect 57 19 58 21
rect 54 -2 58 19
rect 70 21 74 90
rect 70 19 71 21
rect 73 19 74 21
rect 70 -2 74 19
rect 86 21 90 90
rect 86 19 87 21
rect 89 19 90 21
rect 86 -2 90 19
rect 102 21 106 90
rect 102 19 103 21
rect 105 19 106 21
rect 102 -2 106 19
rect 118 21 122 90
rect 118 19 119 21
rect 121 19 122 21
rect 118 -2 122 19
rect 134 21 138 90
rect 134 19 135 21
rect 137 19 138 21
rect 134 -2 138 19
rect 150 21 154 90
rect 150 19 151 21
rect 153 19 154 21
rect 150 -2 154 19
rect 166 21 170 90
rect 166 19 167 21
rect 169 19 170 21
rect 166 -2 170 19
rect 182 21 186 90
rect 182 19 183 21
rect 185 19 186 21
rect 182 -2 186 19
rect 198 21 202 90
rect 198 19 199 21
rect 201 19 202 21
rect 198 -2 202 19
rect 214 21 218 90
rect 214 19 215 21
rect 217 19 218 21
rect 214 -2 218 19
rect 230 21 234 90
rect 230 19 231 21
rect 233 19 234 21
rect 230 -2 234 19
rect 246 21 250 90
rect 246 19 247 21
rect 249 19 250 21
rect 246 -2 250 19
rect 262 21 266 90
rect 262 19 263 21
rect 265 19 266 21
rect 262 -2 266 19
rect 278 21 282 90
rect 278 19 279 21
rect 281 19 282 21
rect 278 -2 282 19
rect 294 21 298 90
rect 294 19 295 21
rect 297 19 298 21
rect 294 -2 298 19
<< alu4 >>
rect -11 77 307 78
rect -11 75 7 77
rect 9 75 307 77
rect -11 74 307 75
rect -11 61 307 62
rect -11 59 7 61
rect 9 59 307 61
rect -11 58 307 59
rect -11 45 307 46
rect -11 43 7 45
rect 9 43 307 45
rect -11 42 307 43
rect -11 29 307 30
rect -11 27 7 29
rect 9 27 307 29
rect -11 26 307 27
rect -11 13 307 14
rect -11 11 -1 13
rect 1 11 7 13
rect 9 11 15 13
rect 17 11 31 13
rect 33 11 47 13
rect 49 11 63 13
rect 65 11 79 13
rect 81 11 95 13
rect 97 11 111 13
rect 113 11 127 13
rect 129 11 143 13
rect 145 11 159 13
rect 161 11 175 13
rect 177 11 191 13
rect 193 11 207 13
rect 209 11 223 13
rect 225 11 239 13
rect 241 11 255 13
rect 257 11 271 13
rect 273 11 287 13
rect 289 11 303 13
rect 305 11 307 13
rect -11 10 307 11
<< alu5 >>
rect -2 13 2 90
rect -2 11 -1 13
rect 1 11 2 13
rect -2 -2 2 11
rect 14 13 18 90
rect 14 11 15 13
rect 17 11 18 13
rect 14 -2 18 11
rect 30 13 34 90
rect 30 11 31 13
rect 33 11 34 13
rect 30 -2 34 11
rect 46 13 50 90
rect 46 11 47 13
rect 49 11 50 13
rect 46 -2 50 11
rect 62 13 66 90
rect 62 11 63 13
rect 65 11 66 13
rect 62 -2 66 11
rect 78 13 82 90
rect 78 11 79 13
rect 81 11 82 13
rect 78 -2 82 11
rect 94 13 98 90
rect 94 11 95 13
rect 97 11 98 13
rect 94 -2 98 11
rect 110 13 114 90
rect 110 11 111 13
rect 113 11 114 13
rect 110 -2 114 11
rect 126 13 130 90
rect 126 11 127 13
rect 129 11 130 13
rect 126 -2 130 11
rect 142 13 146 90
rect 142 11 143 13
rect 145 11 146 13
rect 142 -2 146 11
rect 158 13 162 90
rect 158 11 159 13
rect 161 11 162 13
rect 158 -2 162 11
rect 174 13 178 90
rect 174 11 175 13
rect 177 11 178 13
rect 174 -2 178 11
rect 190 13 194 90
rect 190 11 191 13
rect 193 11 194 13
rect 190 -2 194 11
rect 206 13 210 90
rect 206 11 207 13
rect 209 11 210 13
rect 206 -2 210 11
rect 222 13 226 90
rect 222 11 223 13
rect 225 11 226 13
rect 222 -2 226 11
rect 238 13 242 90
rect 238 11 239 13
rect 241 11 242 13
rect 238 -2 242 11
rect 254 13 258 90
rect 254 11 255 13
rect 257 11 258 13
rect 254 -2 258 11
rect 270 13 274 90
rect 270 11 271 13
rect 273 11 274 13
rect 270 -2 274 11
rect 286 13 290 90
rect 286 11 287 13
rect 289 11 290 13
rect 286 -2 290 11
rect 302 13 306 90
rect 302 11 303 13
rect 305 11 306 13
rect 302 -2 306 11
<< via1 >>
rect -9 67 -7 69
rect -9 51 -7 53
rect -9 35 -7 37
rect -9 19 -7 21
<< via2 >>
rect 7 19 9 21
rect 23 19 25 21
rect 39 19 41 21
rect 55 19 57 21
rect 71 19 73 21
rect 87 19 89 21
rect 103 19 105 21
rect 119 19 121 21
rect 135 19 137 21
rect 151 19 153 21
rect 167 19 169 21
rect 183 19 185 21
rect 199 19 201 21
rect 215 19 217 21
rect 231 19 233 21
rect 247 19 249 21
rect 263 19 265 21
rect 279 19 281 21
rect 295 19 297 21
<< via3 >>
rect 7 75 9 77
rect 7 59 9 61
rect 7 43 9 45
rect 7 27 9 29
rect 7 11 9 13
<< via4 >>
rect -1 11 1 13
rect 15 11 17 13
rect 31 11 33 13
rect 47 11 49 13
rect 63 11 65 13
rect 79 11 81 13
rect 95 11 97 13
rect 111 11 113 13
rect 127 11 129 13
rect 143 11 145 13
rect 159 11 161 13
rect 175 11 177 13
rect 191 11 193 13
rect 207 11 209 13
rect 223 11 225 13
rect 239 11 241 13
rect 255 11 257 13
rect 271 11 273 13
rect 287 11 289 13
rect 303 11 305 13
<< end >>
