magic
tech scmos
timestamp 1199203171
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 23 66 25 70
rect 30 66 32 70
rect 37 66 39 70
rect 13 57 15 62
rect 13 35 15 46
rect 23 36 25 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 34 26 36
rect 19 32 22 34
rect 24 32 26 34
rect 19 30 26 32
rect 9 19 11 29
rect 19 19 21 30
rect 30 28 32 39
rect 37 36 39 39
rect 37 34 47 36
rect 41 32 43 34
rect 45 32 47 34
rect 41 30 47 32
rect 30 26 37 28
rect 30 24 33 26
rect 35 24 37 26
rect 30 22 37 24
rect 31 19 33 22
rect 41 19 43 30
rect 9 5 11 10
rect 19 5 21 10
rect 31 5 33 10
rect 41 5 43 10
<< ndif >>
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 10 9 13
rect 11 16 19 19
rect 11 14 14 16
rect 16 14 19 16
rect 11 10 19 14
rect 21 10 31 19
rect 33 16 41 19
rect 33 14 36 16
rect 38 14 41 16
rect 33 10 41 14
rect 43 14 50 19
rect 43 12 46 14
rect 48 12 50 14
rect 43 10 50 12
rect 23 7 29 10
rect 23 5 25 7
rect 27 5 29 7
rect 23 3 29 5
<< pdif >>
rect 5 57 11 59
rect 18 57 23 66
rect 5 55 7 57
rect 9 55 13 57
rect 5 46 13 55
rect 15 50 23 57
rect 15 48 18 50
rect 20 48 23 50
rect 15 46 23 48
rect 18 39 23 46
rect 25 39 30 66
rect 32 39 37 66
rect 39 64 48 66
rect 39 62 43 64
rect 45 62 48 64
rect 39 57 48 62
rect 39 55 43 57
rect 45 55 48 57
rect 39 39 48 55
<< alu1 >>
rect -2 67 58 72
rect -2 65 5 67
rect 7 65 58 67
rect -2 64 58 65
rect 2 50 22 51
rect 2 48 18 50
rect 20 48 22 50
rect 2 47 22 48
rect 2 45 14 47
rect 2 17 6 45
rect 26 43 30 59
rect 34 45 47 51
rect 18 37 30 43
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 34 26 38 35
rect 42 34 47 45
rect 42 32 43 34
rect 45 32 47 34
rect 42 30 47 32
rect 10 22 23 26
rect 35 24 47 26
rect 34 21 47 24
rect 2 15 4 17
rect 2 13 6 15
rect -2 7 58 8
rect -2 5 25 7
rect 27 5 58 7
rect -2 0 58 5
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 9 10 11 19
rect 19 10 21 19
rect 31 10 33 19
rect 41 10 43 19
<< pmos >>
rect 13 46 15 57
rect 23 39 25 66
rect 30 39 32 66
rect 37 39 39 66
<< polyct0 >>
rect 22 32 24 34
rect 33 24 34 26
<< polyct1 >>
rect 11 31 13 33
rect 43 32 45 34
rect 34 24 35 26
<< ndifct0 >>
rect 14 14 16 16
rect 36 14 38 16
rect 46 12 48 14
<< ndifct1 >>
rect 4 15 6 17
rect 25 5 27 7
<< ntiect1 >>
rect 5 65 7 67
<< pdifct0 >>
rect 7 55 9 57
rect 43 62 45 64
rect 43 55 45 57
<< pdifct1 >>
rect 18 48 20 50
<< alu0 >>
rect 5 57 11 64
rect 41 62 43 64
rect 45 62 47 64
rect 5 55 7 57
rect 9 55 11 57
rect 5 54 11 55
rect 41 57 47 62
rect 41 55 43 57
rect 45 55 47 57
rect 41 54 47 55
rect 20 34 26 37
rect 20 32 22 34
rect 24 32 26 34
rect 20 31 26 32
rect 32 26 34 28
rect 32 24 33 26
rect 32 22 34 24
rect 6 13 7 19
rect 12 16 40 17
rect 12 14 14 16
rect 16 14 36 16
rect 38 14 40 16
rect 12 13 40 14
rect 45 14 49 16
rect 45 12 46 14
rect 48 12 49 14
rect 45 8 49 12
<< labels >>
rlabel alu0 26 15 26 15 6 n3
rlabel alu1 4 32 4 32 6 z
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 20 24 20 24 6 b
rlabel alu1 20 40 20 40 6 a3
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 28 48 28 48 6 a3
rlabel alu1 36 48 36 48 6 a1
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 24 44 24 6 a2
rlabel alu1 44 44 44 44 6 a1
<< end >>
