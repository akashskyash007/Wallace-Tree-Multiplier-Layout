magic
tech scmos
timestamp 1199203298
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 28 70 30 74
rect 35 70 37 74
rect 42 70 44 74
rect 49 70 51 74
rect 9 61 11 65
rect 9 40 11 49
rect 28 40 30 43
rect 9 38 15 40
rect 9 36 11 38
rect 13 36 15 38
rect 9 34 15 36
rect 19 38 30 40
rect 19 36 21 38
rect 23 36 25 38
rect 19 34 25 36
rect 35 34 37 43
rect 9 25 11 34
rect 19 25 21 34
rect 29 32 37 34
rect 29 30 33 32
rect 35 30 37 32
rect 29 28 37 30
rect 42 31 44 43
rect 49 40 51 43
rect 49 38 58 40
rect 52 36 54 38
rect 56 36 58 38
rect 52 34 58 36
rect 42 29 48 31
rect 29 25 31 28
rect 42 27 44 29
rect 46 27 48 29
rect 42 25 48 27
rect 42 22 44 25
rect 52 22 54 34
rect 9 15 11 19
rect 19 15 21 19
rect 29 14 31 19
rect 42 11 44 16
rect 52 11 54 16
<< ndif >>
rect 2 23 9 25
rect 2 21 4 23
rect 6 21 9 23
rect 2 19 9 21
rect 11 19 19 25
rect 21 23 29 25
rect 21 21 24 23
rect 26 21 29 23
rect 21 19 29 21
rect 31 22 40 25
rect 31 19 42 22
rect 13 13 17 19
rect 33 16 42 19
rect 44 20 52 22
rect 44 18 47 20
rect 49 18 52 20
rect 44 16 52 18
rect 54 16 62 22
rect 13 11 19 13
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
rect 33 11 40 16
rect 56 11 62 16
rect 33 9 35 11
rect 37 9 40 11
rect 33 7 40 9
rect 56 9 58 11
rect 60 9 62 11
rect 56 7 62 9
<< pdif >>
rect 13 63 19 65
rect 13 61 15 63
rect 17 61 19 63
rect 4 55 9 61
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 49 9 51
rect 11 59 19 61
rect 11 49 17 59
rect 23 55 28 70
rect 21 53 28 55
rect 21 51 23 53
rect 25 51 28 53
rect 21 49 28 51
rect 23 43 28 49
rect 30 43 35 70
rect 37 43 42 70
rect 44 43 49 70
rect 51 68 59 70
rect 51 66 54 68
rect 56 66 59 68
rect 51 61 59 66
rect 51 59 54 61
rect 56 59 59 61
rect 51 43 59 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 49 7 51
rect 2 23 6 49
rect 34 46 38 63
rect 20 42 38 46
rect 42 46 46 55
rect 42 42 57 46
rect 20 38 24 42
rect 53 38 57 42
rect 20 36 21 38
rect 23 36 24 38
rect 20 34 24 36
rect 32 34 47 38
rect 53 36 54 38
rect 56 36 57 38
rect 53 34 57 36
rect 32 32 38 34
rect 32 30 33 32
rect 35 30 38 32
rect 2 21 4 23
rect 32 25 38 30
rect 42 29 62 30
rect 42 27 44 29
rect 46 27 62 29
rect 42 26 62 27
rect 6 21 16 22
rect 2 17 16 21
rect 58 17 62 26
rect -2 11 66 12
rect -2 9 15 11
rect 17 9 35 11
rect 37 9 58 11
rect 60 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 19 11 25
rect 19 19 21 25
rect 29 19 31 25
rect 42 16 44 22
rect 52 16 54 22
<< pmos >>
rect 9 49 11 61
rect 28 43 30 70
rect 35 43 37 70
rect 42 43 44 70
rect 49 43 51 70
<< polyct0 >>
rect 11 36 13 38
<< polyct1 >>
rect 21 36 23 38
rect 33 30 35 32
rect 54 36 56 38
rect 44 27 46 29
<< ndifct0 >>
rect 24 21 26 23
rect 47 18 49 20
<< ndifct1 >>
rect 4 21 6 23
rect 15 9 17 11
rect 35 9 37 11
rect 58 9 60 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 15 61 17 63
rect 23 51 25 53
rect 54 66 56 68
rect 54 59 56 61
<< pdifct1 >>
rect 4 51 6 53
<< alu0 >>
rect 14 63 18 68
rect 52 66 54 68
rect 56 66 58 68
rect 14 61 15 63
rect 17 61 18 63
rect 14 59 18 61
rect 11 53 27 54
rect 11 51 23 53
rect 25 51 27 53
rect 11 50 27 51
rect 11 40 15 50
rect 52 61 58 66
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
rect 10 38 15 40
rect 10 36 11 38
rect 13 36 15 38
rect 10 34 15 36
rect 11 30 15 34
rect 11 26 27 30
rect 6 22 7 25
rect 23 23 27 26
rect 23 21 24 23
rect 26 21 27 23
rect 23 20 51 21
rect 23 18 47 20
rect 49 18 51 20
rect 23 17 51 18
<< labels >>
rlabel alu0 13 40 13 40 6 zn
rlabel alu0 25 23 25 23 6 zn
rlabel alu0 19 52 19 52 6 zn
rlabel alu0 37 19 37 19 6 zn
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 28 44 28 44 6 d
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 36 32 36 32 6 c
rlabel alu1 44 36 44 36 6 c
rlabel alu1 36 56 36 56 6 d
rlabel alu1 44 52 44 52 6 a
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 60 20 60 20 6 b
rlabel alu1 52 28 52 28 6 b
rlabel alu1 52 44 52 44 6 a
<< end >>
