magic
tech scmos
timestamp 1199542332
<< ab >>
rect 0 0 40 100
<< nwell >>
rect -5 48 45 105
<< pwell >>
rect -5 -5 45 48
<< poly >>
rect 13 86 15 90
rect 25 85 27 89
rect 13 63 15 66
rect 7 61 15 63
rect 7 59 9 61
rect 11 59 15 61
rect 7 57 15 59
rect 13 34 15 57
rect 25 43 27 65
rect 25 41 33 43
rect 25 39 29 41
rect 31 39 33 41
rect 21 37 33 39
rect 21 34 23 37
rect 13 11 15 15
rect 21 11 23 15
<< ndif >>
rect 5 15 13 34
rect 15 15 21 34
rect 23 21 31 34
rect 23 19 27 21
rect 29 19 31 21
rect 23 15 31 19
rect 5 11 11 15
rect 5 9 7 11
rect 9 9 11 11
rect 5 7 11 9
<< pdif >>
rect 5 91 11 93
rect 5 89 7 91
rect 9 89 11 91
rect 29 91 35 93
rect 5 86 11 89
rect 29 89 31 91
rect 33 89 35 91
rect 5 66 13 86
rect 15 85 23 86
rect 29 85 35 89
rect 15 81 25 85
rect 15 79 19 81
rect 21 79 25 81
rect 15 71 25 79
rect 15 69 19 71
rect 21 69 25 71
rect 15 66 25 69
rect 20 65 25 66
rect 27 65 35 85
<< alu1 >>
rect -2 91 42 100
rect -2 89 7 91
rect 9 89 31 91
rect 33 89 42 91
rect -2 88 42 89
rect 8 61 12 83
rect 8 59 9 61
rect 11 59 12 61
rect 8 17 12 59
rect 18 81 22 83
rect 18 79 19 81
rect 21 79 22 81
rect 18 71 22 79
rect 18 69 19 71
rect 21 69 22 71
rect 18 22 22 69
rect 28 41 32 83
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 18 21 31 22
rect 18 19 27 21
rect 29 19 31 21
rect 18 18 31 19
rect 18 17 22 18
rect -2 11 42 12
rect -2 9 7 11
rect 9 9 42 11
rect -2 7 42 9
rect -2 5 24 7
rect 26 5 42 7
rect -2 0 42 5
<< ptie >>
rect 22 7 34 9
rect 22 5 24 7
rect 26 5 34 7
rect 22 3 34 5
<< nmos >>
rect 13 15 15 34
rect 21 15 23 34
<< pmos >>
rect 13 66 15 86
rect 25 65 27 85
<< polyct1 >>
rect 9 59 11 61
rect 29 39 31 41
<< ndifct1 >>
rect 27 19 29 21
rect 7 9 9 11
<< ptiect1 >>
rect 24 5 26 7
<< pdifct1 >>
rect 7 89 9 91
rect 31 89 33 91
rect 19 79 21 81
rect 19 69 21 71
<< labels >>
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 10 50 10 50 6 i0
rlabel alu1 20 50 20 50 6 nq
rlabel alu1 20 94 20 94 6 vdd
rlabel alu1 30 55 30 55 6 i1
<< end >>
