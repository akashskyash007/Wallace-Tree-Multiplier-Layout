magic
tech scmos
timestamp 1199542750
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -2 48 82 104
<< pwell >>
rect -2 -4 82 48
<< poly >>
rect 11 95 13 98
rect 19 95 21 98
rect 27 95 29 98
rect 43 95 45 98
rect 55 95 57 98
rect 67 75 69 78
rect 11 33 13 55
rect 19 43 21 55
rect 27 53 29 55
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 37 49
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 7 31 13 33
rect 7 29 9 31
rect 11 29 13 31
rect 7 27 13 29
rect 19 29 21 37
rect 19 27 25 29
rect 11 25 13 27
rect 23 25 25 27
rect 35 25 37 47
rect 43 43 45 55
rect 55 43 57 55
rect 67 53 69 55
rect 61 51 69 53
rect 61 49 63 51
rect 65 49 69 51
rect 61 47 69 49
rect 43 41 63 43
rect 43 39 59 41
rect 61 39 63 41
rect 43 37 63 39
rect 45 25 47 37
rect 57 25 59 37
rect 67 25 69 47
rect 11 12 13 15
rect 23 12 25 15
rect 35 12 37 15
rect 67 12 69 15
rect 45 2 47 5
rect 57 2 59 5
<< ndif >>
rect 3 21 11 25
rect 3 19 5 21
rect 7 19 11 21
rect 3 15 11 19
rect 13 15 23 25
rect 25 21 35 25
rect 25 19 29 21
rect 31 19 35 21
rect 25 15 35 19
rect 37 15 45 25
rect 15 11 21 15
rect 15 9 17 11
rect 19 9 21 11
rect 39 9 45 15
rect 15 7 21 9
rect 37 7 45 9
rect 37 5 39 7
rect 41 5 45 7
rect 47 21 57 25
rect 47 19 51 21
rect 53 19 57 21
rect 47 5 57 19
rect 59 15 67 25
rect 69 21 77 25
rect 69 19 73 21
rect 75 19 77 21
rect 69 15 77 19
rect 59 9 65 15
rect 59 7 67 9
rect 59 5 63 7
rect 65 5 67 7
rect 37 3 43 5
rect 61 3 67 5
<< pdif >>
rect 3 81 11 95
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 55 19 95
rect 21 55 27 95
rect 29 91 43 95
rect 29 89 37 91
rect 39 89 43 91
rect 29 55 43 89
rect 45 71 55 95
rect 45 69 49 71
rect 51 69 55 71
rect 45 61 55 69
rect 45 59 49 61
rect 51 59 55 61
rect 45 55 55 59
rect 57 91 65 95
rect 57 89 61 91
rect 63 89 65 91
rect 57 75 65 89
rect 57 55 67 75
rect 69 61 77 75
rect 69 59 73 61
rect 75 59 77 61
rect 69 55 77 59
<< alu1 >>
rect -2 95 82 100
rect -2 93 73 95
rect 75 93 82 95
rect -2 91 82 93
rect -2 89 37 91
rect 39 89 61 91
rect 63 89 82 91
rect -2 88 82 89
rect 4 81 8 82
rect 4 79 5 81
rect 7 79 65 81
rect 4 78 8 79
rect 8 31 12 72
rect 8 29 9 31
rect 11 29 12 31
rect 8 28 12 29
rect 18 41 22 72
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 28 51 32 72
rect 28 49 29 51
rect 31 49 32 51
rect 28 28 32 49
rect 4 21 8 22
rect 28 21 32 22
rect 39 21 41 79
rect 4 19 5 21
rect 7 19 29 21
rect 31 19 41 21
rect 48 71 52 72
rect 48 69 49 71
rect 51 69 52 71
rect 48 61 52 69
rect 48 59 49 61
rect 51 59 52 61
rect 48 22 52 59
rect 63 52 65 79
rect 72 61 76 62
rect 72 59 73 61
rect 75 59 76 61
rect 72 58 76 59
rect 62 51 66 52
rect 62 49 63 51
rect 65 49 66 51
rect 62 48 66 49
rect 58 41 62 42
rect 73 41 75 58
rect 58 39 59 41
rect 61 39 75 41
rect 58 38 62 39
rect 73 22 75 39
rect 48 21 54 22
rect 48 19 51 21
rect 53 19 54 21
rect 4 18 8 19
rect 28 18 32 19
rect 48 18 54 19
rect 72 21 76 22
rect 72 19 73 21
rect 75 19 76 21
rect 72 18 76 19
rect -2 11 82 12
rect -2 9 17 11
rect 19 9 82 11
rect -2 7 82 9
rect -2 5 39 7
rect 41 5 63 7
rect 65 5 82 7
rect -2 0 82 5
<< ntie >>
rect 71 95 77 97
rect 71 93 73 95
rect 75 93 77 95
rect 71 85 77 93
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 35 15 37 25
rect 45 5 47 25
rect 57 5 59 25
rect 67 15 69 25
<< pmos >>
rect 11 55 13 95
rect 19 55 21 95
rect 27 55 29 95
rect 43 55 45 95
rect 55 55 57 95
rect 67 55 69 75
<< polyct1 >>
rect 29 49 31 51
rect 19 39 21 41
rect 9 29 11 31
rect 63 49 65 51
rect 59 39 61 41
<< ndifct1 >>
rect 5 19 7 21
rect 29 19 31 21
rect 17 9 19 11
rect 39 5 41 7
rect 51 19 53 21
rect 73 19 75 21
rect 63 5 65 7
<< ntiect1 >>
rect 73 93 75 95
<< pdifct1 >>
rect 5 79 7 81
rect 37 89 39 91
rect 49 69 51 71
rect 49 59 51 61
rect 61 89 63 91
rect 73 59 75 61
<< labels >>
rlabel alu1 10 50 10 50 6 i2
rlabel polyct1 30 50 30 50 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel ndifct1 40 6 40 6 6 vss
rlabel alu1 50 45 50 45 6 nq
rlabel alu1 40 94 40 94 6 vdd
<< end >>
