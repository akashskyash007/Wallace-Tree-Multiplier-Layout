magic
tech scmos
timestamp 1199202441
<< ab >>
rect 0 0 80 80
<< nwell >>
rect -5 36 85 88
<< pwell >>
rect -5 -8 85 36
<< poly >>
rect 42 72 71 74
rect 9 60 11 65
rect 35 64 37 69
rect 42 64 44 72
rect 52 64 54 68
rect 59 64 61 68
rect 69 64 71 72
rect 19 54 21 59
rect 35 55 37 58
rect 31 53 37 55
rect 31 51 33 53
rect 35 51 37 53
rect 31 49 37 51
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 31 39
rect 10 20 12 37
rect 24 35 27 37
rect 29 35 31 37
rect 24 33 31 35
rect 24 30 26 33
rect 35 24 37 49
rect 42 39 44 58
rect 52 49 54 52
rect 48 47 54 49
rect 59 47 61 52
rect 48 45 50 47
rect 52 45 54 47
rect 48 43 54 45
rect 58 45 64 47
rect 58 43 60 45
rect 62 43 64 45
rect 58 41 64 43
rect 42 37 54 39
rect 41 31 47 33
rect 41 29 43 31
rect 45 29 47 31
rect 41 27 47 29
rect 42 24 44 27
rect 52 24 54 37
rect 59 24 61 41
rect 69 37 71 52
rect 65 35 71 37
rect 65 33 67 35
rect 69 33 71 35
rect 65 31 71 33
rect 69 28 71 31
rect 24 19 26 24
rect 35 13 37 18
rect 42 13 44 18
rect 52 13 54 18
rect 59 13 61 18
rect 69 17 71 22
rect 10 6 12 11
<< ndif >>
rect 2 20 8 22
rect 17 28 24 30
rect 17 26 19 28
rect 21 26 24 28
rect 17 24 24 26
rect 26 28 33 30
rect 26 26 29 28
rect 31 26 33 28
rect 26 24 33 26
rect 63 24 69 28
rect 2 18 4 20
rect 6 18 10 20
rect 2 16 10 18
rect 5 11 10 16
rect 12 15 19 20
rect 28 18 35 24
rect 37 18 42 24
rect 44 22 52 24
rect 44 20 47 22
rect 49 20 52 22
rect 44 18 52 20
rect 54 18 59 24
rect 61 22 69 24
rect 71 26 78 28
rect 71 24 74 26
rect 76 24 78 26
rect 71 22 78 24
rect 61 18 67 22
rect 12 13 15 15
rect 17 13 19 15
rect 63 15 67 18
rect 12 11 19 13
rect 63 11 69 15
rect 63 9 65 11
rect 67 9 69 11
rect 63 7 69 9
<< pdif >>
rect 28 62 35 64
rect 28 60 30 62
rect 32 60 35 62
rect 4 55 9 60
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 54 17 60
rect 28 58 35 60
rect 37 58 42 64
rect 44 62 52 64
rect 44 60 47 62
rect 49 60 52 62
rect 44 58 52 60
rect 11 52 19 54
rect 11 50 14 52
rect 16 50 19 52
rect 11 42 19 50
rect 21 52 28 54
rect 21 50 24 52
rect 26 50 28 52
rect 21 48 28 50
rect 21 42 26 48
rect 47 52 52 58
rect 54 52 59 64
rect 61 62 69 64
rect 61 60 64 62
rect 66 60 69 62
rect 61 52 69 60
rect 71 58 76 64
rect 71 56 78 58
rect 71 54 74 56
rect 76 54 78 56
rect 71 52 78 54
<< alu1 >>
rect -2 81 82 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 82 81
rect -2 68 82 79
rect 2 53 7 55
rect 2 51 4 53
rect 6 51 7 53
rect 2 46 7 51
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 2 31 6 42
rect 2 25 14 31
rect 2 20 8 25
rect 2 18 4 20
rect 6 18 8 20
rect 2 17 8 18
rect 58 45 63 47
rect 58 43 60 45
rect 62 43 63 45
rect 58 41 63 43
rect 58 30 62 41
rect 49 26 62 30
rect 66 35 70 37
rect 66 33 67 35
rect 69 33 70 35
rect 66 22 70 33
rect 57 18 70 22
rect -2 11 82 12
rect -2 9 65 11
rect 67 9 82 11
rect -2 1 82 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 82 1
rect -2 -2 82 -1
<< ptie >>
rect 0 1 80 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 80 1
rect 0 -3 80 -1
<< ntie >>
rect 0 81 80 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 80 81
rect 0 77 80 79
<< nmos >>
rect 24 24 26 30
rect 10 11 12 20
rect 35 18 37 24
rect 42 18 44 24
rect 52 18 54 24
rect 59 18 61 24
rect 69 22 71 28
<< pmos >>
rect 9 42 11 60
rect 35 58 37 64
rect 42 58 44 64
rect 19 42 21 54
rect 52 52 54 64
rect 59 52 61 64
rect 69 52 71 64
<< polyct0 >>
rect 33 51 35 53
rect 27 35 29 37
rect 50 45 52 47
rect 43 29 45 31
<< polyct1 >>
rect 60 43 62 45
rect 67 33 69 35
<< ndifct0 >>
rect 19 26 21 28
rect 29 26 31 28
rect 47 20 49 22
rect 74 24 76 26
rect 15 13 17 15
<< ndifct1 >>
rect 4 18 6 20
rect 65 9 67 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
<< pdifct0 >>
rect 30 60 32 62
rect 47 60 49 62
rect 14 50 16 52
rect 24 50 26 52
rect 64 60 66 62
rect 74 54 76 56
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 12 52 18 68
rect 29 62 33 68
rect 29 60 30 62
rect 32 60 33 62
rect 29 58 33 60
rect 41 62 51 63
rect 41 60 47 62
rect 49 60 51 62
rect 41 59 51 60
rect 63 62 67 68
rect 63 60 64 62
rect 66 60 67 62
rect 12 50 14 52
rect 16 50 18 52
rect 12 49 18 50
rect 23 53 37 54
rect 23 52 33 53
rect 23 50 24 52
rect 26 51 33 52
rect 35 51 37 53
rect 26 50 37 51
rect 23 46 27 50
rect 41 46 45 59
rect 63 58 67 60
rect 73 56 77 58
rect 73 54 74 56
rect 76 54 77 56
rect 18 42 27 46
rect 35 42 45 46
rect 49 50 78 54
rect 49 47 53 50
rect 49 45 50 47
rect 52 45 53 47
rect 18 28 22 42
rect 35 38 39 42
rect 49 38 53 45
rect 25 37 39 38
rect 25 35 27 37
rect 29 35 39 37
rect 25 34 39 35
rect 18 26 19 28
rect 21 26 22 28
rect 18 24 22 26
rect 28 28 32 30
rect 28 26 29 28
rect 31 26 32 28
rect 14 15 18 17
rect 14 13 15 15
rect 17 13 18 15
rect 14 12 18 13
rect 28 12 32 26
rect 35 23 39 34
rect 42 34 53 38
rect 42 31 46 34
rect 42 29 43 31
rect 45 29 46 31
rect 42 27 46 29
rect 35 22 51 23
rect 74 28 78 50
rect 73 26 78 28
rect 73 24 74 26
rect 76 24 78 26
rect 73 22 78 24
rect 35 20 47 22
rect 49 20 51 22
rect 35 19 51 20
<< labels >>
rlabel alu0 32 36 32 36 6 n1
rlabel alu0 25 48 25 48 6 n2
rlabel alu0 20 35 20 35 6 n2
rlabel alu0 30 52 30 52 6 n2
rlabel alu0 43 21 43 21 6 n1
rlabel alu0 44 32 44 32 6 en
rlabel alu0 51 44 51 44 6 en
rlabel alu0 46 61 46 61 6 n1
rlabel alu0 76 38 76 38 6 en
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 52 28 52 28 6 d
rlabel alu1 40 74 40 74 6 vdd
rlabel alu1 60 20 60 20 6 e
rlabel alu1 68 28 68 28 6 e
rlabel alu1 60 40 60 40 6 d
<< end >>
