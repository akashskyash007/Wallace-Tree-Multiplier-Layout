magic
tech scmos
timestamp 1199203194
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 9 68 11 73
rect 16 68 18 73
rect 29 68 31 73
rect 36 68 38 73
rect 9 39 11 48
rect 16 45 18 48
rect 29 45 31 48
rect 16 43 21 45
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 9 23 11 33
rect 19 32 21 43
rect 25 43 31 45
rect 36 45 38 48
rect 36 43 41 45
rect 25 41 27 43
rect 29 41 31 43
rect 25 39 31 41
rect 19 30 25 32
rect 19 28 21 30
rect 23 28 25 30
rect 19 26 25 28
rect 19 23 21 26
rect 29 23 31 39
rect 39 32 41 43
rect 39 30 48 32
rect 39 28 44 30
rect 46 28 48 30
rect 39 26 48 28
rect 39 23 41 26
rect 9 12 11 17
rect 19 12 21 17
rect 29 12 31 17
rect 39 12 41 17
<< ndif >>
rect 2 21 9 23
rect 2 19 4 21
rect 6 19 9 21
rect 2 17 9 19
rect 11 21 19 23
rect 11 19 14 21
rect 16 19 19 21
rect 11 17 19 19
rect 21 21 29 23
rect 21 19 24 21
rect 26 19 29 21
rect 21 17 29 19
rect 31 21 39 23
rect 31 19 34 21
rect 36 19 39 21
rect 31 17 39 19
rect 41 21 48 23
rect 41 19 44 21
rect 46 19 48 21
rect 41 17 48 19
<< pdif >>
rect 4 63 9 68
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 48 9 50
rect 11 48 16 68
rect 18 65 29 68
rect 18 63 23 65
rect 25 63 29 65
rect 18 48 29 63
rect 31 48 36 68
rect 38 61 43 68
rect 38 59 47 61
rect 38 57 43 59
rect 45 57 47 59
rect 38 52 47 57
rect 38 50 43 52
rect 45 50 47 52
rect 38 48 47 50
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 2 61 14 63
rect 2 59 4 61
rect 6 59 14 61
rect 2 57 14 59
rect 2 54 6 57
rect 2 52 4 54
rect 2 29 6 52
rect 26 49 38 55
rect 18 42 22 47
rect 10 38 22 42
rect 26 43 30 49
rect 26 41 27 43
rect 29 41 30 43
rect 26 39 30 41
rect 10 37 14 38
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 50 31 54 39
rect 2 25 15 29
rect 42 30 54 31
rect 42 28 44 30
rect 46 28 54 30
rect 11 22 15 25
rect 11 21 18 22
rect 11 19 14 21
rect 16 19 18 21
rect 11 18 18 19
rect 42 25 54 28
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 17 11 23
rect 19 17 21 23
rect 29 17 31 23
rect 39 17 41 23
<< pmos >>
rect 9 48 11 68
rect 16 48 18 68
rect 29 48 31 68
rect 36 48 38 68
<< polyct0 >>
rect 21 28 23 30
<< polyct1 >>
rect 11 35 13 37
rect 27 41 29 43
rect 44 28 46 30
<< ndifct0 >>
rect 4 19 6 21
rect 24 19 26 21
rect 34 19 36 21
rect 44 19 46 21
<< ndifct1 >>
rect 14 19 16 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 23 63 25 65
rect 43 57 45 59
rect 43 50 45 52
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
<< alu0 >>
rect 22 65 26 68
rect 22 63 23 65
rect 25 63 26 65
rect 22 61 26 63
rect 42 59 46 61
rect 42 57 43 59
rect 45 57 46 59
rect 6 50 7 57
rect 42 52 46 57
rect 42 50 43 52
rect 45 50 46 52
rect 42 42 46 50
rect 34 38 46 42
rect 34 31 38 38
rect 19 30 38 31
rect 19 28 21 30
rect 23 28 38 30
rect 19 27 38 28
rect 2 21 8 22
rect 2 19 4 21
rect 6 19 8 21
rect 2 12 8 19
rect 23 21 27 23
rect 23 19 24 21
rect 26 19 27 21
rect 23 12 27 19
rect 33 21 37 27
rect 33 19 34 21
rect 36 19 37 21
rect 33 17 37 19
rect 42 21 48 22
rect 42 19 44 21
rect 46 19 48 21
rect 42 12 48 19
<< labels >>
rlabel alu0 35 24 35 24 6 an
rlabel alu0 28 29 28 29 6 an
rlabel alu0 44 49 44 49 6 an
rlabel alu1 4 44 4 44 6 z
rlabel polyct1 12 36 12 36 6 b
rlabel alu1 20 44 20 44 6 b
rlabel alu1 12 60 12 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 48 28 48 6 a1
rlabel alu1 36 52 36 52 6 a1
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 28 44 28 6 a2
rlabel alu1 52 32 52 32 6 a2
<< end >>
