magic
tech scmos
timestamp 1199201957
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 31 64 33 69
rect 41 64 43 69
rect 53 64 55 69
rect 9 54 11 59
rect 9 39 11 42
rect 31 39 33 48
rect 41 39 43 48
rect 53 45 55 48
rect 53 43 62 45
rect 53 41 58 43
rect 60 41 62 43
rect 53 39 62 41
rect 9 37 19 39
rect 13 35 15 37
rect 17 35 19 37
rect 13 33 19 35
rect 31 37 37 39
rect 31 35 33 37
rect 35 35 37 37
rect 31 33 37 35
rect 41 37 47 39
rect 41 35 43 37
rect 45 35 47 37
rect 41 33 47 35
rect 13 30 15 33
rect 13 19 15 24
rect 31 23 33 33
rect 41 23 43 33
rect 53 28 55 39
rect 48 26 55 28
rect 48 23 50 26
rect 31 12 33 17
rect 41 11 43 16
rect 48 11 50 16
<< ndif >>
rect 6 28 13 30
rect 6 26 8 28
rect 10 26 13 28
rect 6 24 13 26
rect 15 28 23 30
rect 15 26 19 28
rect 21 26 23 28
rect 15 24 23 26
rect 17 23 23 24
rect 17 21 31 23
rect 17 19 19 21
rect 21 19 26 21
rect 28 19 31 21
rect 17 17 31 19
rect 33 21 41 23
rect 33 19 36 21
rect 38 19 41 21
rect 33 17 41 19
rect 36 16 41 17
rect 43 16 48 23
rect 50 20 57 23
rect 50 18 53 20
rect 55 18 57 20
rect 50 16 57 18
<< pdif >>
rect 45 71 51 73
rect 45 69 47 71
rect 49 69 51 71
rect 45 64 51 69
rect 26 61 31 64
rect 24 59 31 61
rect 24 57 26 59
rect 28 57 31 59
rect 4 48 9 54
rect 2 46 9 48
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 52 18 54
rect 11 50 14 52
rect 16 50 18 52
rect 11 42 18 50
rect 24 52 31 57
rect 24 50 26 52
rect 28 50 31 52
rect 24 48 31 50
rect 33 62 41 64
rect 33 60 36 62
rect 38 60 41 62
rect 33 48 41 60
rect 43 48 53 64
rect 55 62 62 64
rect 55 60 58 62
rect 60 60 62 62
rect 55 58 62 60
rect 55 48 60 58
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 71 66 79
rect -2 69 47 71
rect 49 69 66 71
rect -2 68 66 69
rect 2 46 7 48
rect 2 44 4 46
rect 6 44 7 46
rect 2 42 7 44
rect 2 31 6 42
rect 34 49 46 55
rect 50 49 62 55
rect 34 39 38 49
rect 57 43 62 49
rect 57 41 58 43
rect 60 41 62 43
rect 57 39 62 41
rect 2 28 14 31
rect 32 37 38 39
rect 32 35 33 37
rect 35 35 38 37
rect 32 33 38 35
rect 42 37 46 39
rect 42 35 43 37
rect 45 35 46 37
rect 42 30 46 35
rect 2 26 8 28
rect 10 26 14 28
rect 2 25 14 26
rect 42 26 55 30
rect 2 17 6 25
rect -2 1 66 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 13 24 15 30
rect 31 17 33 23
rect 41 16 43 23
rect 48 16 50 23
<< pmos >>
rect 9 42 11 54
rect 31 48 33 64
rect 41 48 43 64
rect 53 48 55 64
<< polyct0 >>
rect 15 35 17 37
<< polyct1 >>
rect 58 41 60 43
rect 33 35 35 37
rect 43 35 45 37
<< ndifct0 >>
rect 19 26 21 28
rect 19 19 21 21
rect 26 19 28 21
rect 36 19 38 21
rect 53 18 55 20
<< ndifct1 >>
rect 8 26 10 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 26 57 28 59
rect 14 50 16 52
rect 26 50 28 52
rect 36 60 38 62
rect 58 60 60 62
<< pdifct1 >>
rect 47 69 49 71
rect 4 44 6 46
<< alu0 >>
rect 13 52 17 68
rect 34 62 62 63
rect 13 50 14 52
rect 16 50 17 52
rect 13 48 17 50
rect 25 59 29 61
rect 34 60 36 62
rect 38 60 58 62
rect 60 60 62 62
rect 34 59 62 60
rect 25 57 26 59
rect 28 57 29 59
rect 25 52 29 57
rect 25 50 26 52
rect 28 50 29 52
rect 25 38 29 50
rect 13 37 29 38
rect 13 35 15 37
rect 17 35 29 37
rect 13 34 29 35
rect 25 30 29 34
rect 18 28 22 30
rect 18 26 19 28
rect 21 26 22 28
rect 25 26 39 30
rect 18 22 22 26
rect 18 21 30 22
rect 18 19 19 21
rect 21 19 26 21
rect 28 19 30 21
rect 18 18 30 19
rect 35 21 39 26
rect 35 19 36 21
rect 38 19 39 21
rect 18 12 22 18
rect 35 17 39 19
rect 52 20 56 22
rect 52 18 53 20
rect 55 18 56 20
rect 52 12 56 18
<< labels >>
rlabel alu0 48 61 48 61 6 n1
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 28 12 28 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel polyct1 44 36 44 36 6 a2
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 52 44 52 6 b
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 a2
rlabel alu1 52 52 52 52 6 a1
rlabel alu1 60 48 60 48 6 a1
<< end >>
