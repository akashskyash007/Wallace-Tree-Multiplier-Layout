magic
tech scmos
timestamp 1199202554
<< ab >>
rect 0 0 48 72
<< nwell >>
rect -5 32 53 77
<< pwell >>
rect -5 -5 53 32
<< poly >>
rect 10 62 12 67
rect 20 62 22 67
rect 32 56 34 61
rect 10 34 12 38
rect 20 34 22 38
rect 32 35 34 38
rect 9 32 15 34
rect 9 30 11 32
rect 13 30 15 32
rect 9 28 15 30
rect 19 32 25 34
rect 19 30 21 32
rect 23 30 25 32
rect 19 28 25 30
rect 32 33 39 35
rect 32 31 35 33
rect 37 31 39 33
rect 32 29 39 31
rect 12 25 14 28
rect 19 25 21 28
rect 33 25 35 29
rect 33 11 35 16
rect 12 2 14 6
rect 19 2 21 6
<< ndif >>
rect 7 18 12 25
rect 5 16 12 18
rect 5 14 7 16
rect 9 14 12 16
rect 5 12 12 14
rect 7 6 12 12
rect 14 6 19 25
rect 21 17 33 25
rect 21 15 27 17
rect 29 16 33 17
rect 35 23 42 25
rect 35 21 38 23
rect 40 21 42 23
rect 35 19 42 21
rect 35 16 40 19
rect 29 15 31 16
rect 21 10 31 15
rect 21 8 27 10
rect 29 8 31 10
rect 21 6 31 8
<< pdif >>
rect 2 59 10 62
rect 2 57 4 59
rect 6 57 10 59
rect 2 38 10 57
rect 12 58 20 62
rect 12 56 15 58
rect 17 56 20 58
rect 12 38 20 56
rect 22 59 30 62
rect 22 57 26 59
rect 28 57 30 59
rect 22 56 30 57
rect 22 38 32 56
rect 34 52 39 56
rect 34 50 41 52
rect 34 48 37 50
rect 39 48 41 50
rect 34 46 41 48
rect 34 38 39 46
<< alu1 >>
rect -2 67 50 72
rect -2 65 36 67
rect 38 65 50 67
rect -2 64 50 65
rect 10 58 19 59
rect 10 56 15 58
rect 17 56 19 58
rect 10 55 19 56
rect 10 51 14 55
rect 2 45 14 51
rect 2 17 6 45
rect 10 32 14 35
rect 10 30 11 32
rect 13 30 14 32
rect 10 25 14 30
rect 26 37 38 43
rect 34 33 38 37
rect 34 31 35 33
rect 37 31 38 33
rect 34 29 38 31
rect 10 21 22 25
rect 2 16 11 17
rect 2 14 7 16
rect 9 14 11 16
rect 2 13 11 14
rect 18 13 22 21
rect -2 7 50 8
rect -2 5 37 7
rect 39 5 50 7
rect -2 0 50 5
<< ptie >>
rect 35 7 41 9
rect 35 5 37 7
rect 39 5 41 7
rect 35 3 41 5
<< ntie >>
rect 34 67 40 69
rect 34 65 36 67
rect 38 65 40 67
rect 34 63 40 65
<< nmos >>
rect 12 6 14 25
rect 19 6 21 25
rect 33 16 35 25
<< pmos >>
rect 10 38 12 62
rect 20 38 22 62
rect 32 38 34 56
<< polyct0 >>
rect 21 30 23 32
<< polyct1 >>
rect 11 30 13 32
rect 35 31 37 33
<< ndifct0 >>
rect 27 15 29 17
rect 38 21 40 23
rect 27 8 29 10
<< ndifct1 >>
rect 7 14 9 16
<< ntiect1 >>
rect 36 65 38 67
<< ptiect1 >>
rect 37 5 39 7
<< pdifct0 >>
rect 4 57 6 59
rect 26 57 28 59
rect 37 48 39 50
<< pdifct1 >>
rect 15 56 17 58
<< alu0 >>
rect 3 59 7 64
rect 25 59 29 64
rect 3 57 4 59
rect 6 57 7 59
rect 3 55 7 57
rect 25 57 26 59
rect 28 57 29 59
rect 25 55 29 57
rect 18 50 41 51
rect 18 48 37 50
rect 39 48 41 50
rect 18 47 41 48
rect 18 33 22 47
rect 18 32 30 33
rect 18 30 21 32
rect 23 30 30 32
rect 18 29 30 30
rect 26 25 30 29
rect 26 23 42 25
rect 26 21 38 23
rect 40 21 42 23
rect 36 20 42 21
rect 25 17 31 18
rect 25 15 27 17
rect 29 15 31 17
rect 25 10 31 15
rect 25 8 27 10
rect 29 8 31 10
<< labels >>
rlabel alu0 34 23 34 23 6 an
rlabel alu0 24 31 24 31 6 an
rlabel alu0 29 49 29 49 6 an
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 16 20 16 6 b
rlabel alu1 12 28 12 28 6 b
rlabel alu1 12 52 12 52 6 z
rlabel alu1 24 4 24 4 6 vss
rlabel alu1 28 40 28 40 6 a
rlabel alu1 24 68 24 68 6 vdd
rlabel alu1 36 36 36 36 6 a
<< end >>
