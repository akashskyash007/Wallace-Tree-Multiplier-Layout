magic
tech scmos
timestamp 1199202766
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 68
rect 9 36 11 53
rect 19 47 21 53
rect 19 45 25 47
rect 19 43 21 45
rect 23 43 25 45
rect 19 41 25 43
rect 9 34 17 36
rect 9 32 11 34
rect 13 32 17 34
rect 9 30 17 32
rect 15 27 17 30
rect 22 27 24 41
rect 29 39 31 53
rect 29 37 35 39
rect 29 35 31 37
rect 33 35 35 37
rect 29 33 35 35
rect 29 27 31 33
rect 15 12 17 17
rect 22 12 24 17
rect 29 12 31 17
<< ndif >>
rect 10 23 15 27
rect 8 21 15 23
rect 8 19 10 21
rect 12 19 15 21
rect 8 17 15 19
rect 17 17 22 27
rect 24 17 29 27
rect 31 21 38 27
rect 31 19 34 21
rect 36 19 38 21
rect 31 17 38 19
<< pdif >>
rect 4 59 9 63
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 53 9 55
rect 11 61 19 63
rect 11 59 14 61
rect 16 59 19 61
rect 11 53 19 59
rect 21 57 29 63
rect 21 55 24 57
rect 26 55 29 57
rect 21 53 29 55
rect 31 61 38 63
rect 31 59 34 61
rect 36 59 38 61
rect 31 53 38 59
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 57 7 63
rect 2 55 4 57
rect 6 55 7 57
rect 2 54 7 55
rect 23 57 27 59
rect 23 55 24 57
rect 26 55 27 57
rect 23 54 27 55
rect 2 50 27 54
rect 2 17 6 50
rect 34 46 38 55
rect 17 45 38 46
rect 17 43 21 45
rect 23 43 38 45
rect 17 42 38 43
rect 25 37 38 38
rect 10 34 14 36
rect 25 35 31 37
rect 33 35 38 37
rect 25 34 38 35
rect 10 32 11 34
rect 13 32 14 34
rect 10 30 14 32
rect 10 25 23 30
rect 34 25 38 34
rect 18 17 23 25
rect -2 1 42 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 15 17 17 27
rect 22 17 24 27
rect 29 17 31 27
<< pmos >>
rect 9 53 11 63
rect 19 53 21 63
rect 29 53 31 63
<< polyct1 >>
rect 21 43 23 45
rect 11 32 13 34
rect 31 35 33 37
<< ndifct0 >>
rect 10 19 12 21
rect 34 19 36 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 59 16 61
rect 34 59 36 61
<< pdifct1 >>
rect 4 55 6 57
rect 24 55 26 57
<< alu0 >>
rect 12 61 18 68
rect 12 59 14 61
rect 16 59 18 61
rect 32 61 38 68
rect 32 59 34 61
rect 36 59 38 61
rect 12 58 18 59
rect 32 58 38 59
rect 6 21 14 22
rect 6 19 10 21
rect 12 19 14 21
rect 6 18 14 19
rect 32 21 38 22
rect 32 19 34 21
rect 36 19 38 21
rect 32 12 38 19
<< labels >>
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 28 12 28 6 c
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 24 20 24 6 c
rlabel alu1 28 36 28 36 6 a
rlabel alu1 28 44 28 44 6 b
rlabel alu1 20 44 20 44 6 b
rlabel alu1 20 52 20 52 6 z
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 52 36 52 6 b
<< end >>
