magic
tech scmos
timestamp 1199201940
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 68
rect 39 63 41 68
rect 49 63 51 68
rect 59 63 61 68
rect 9 35 11 46
rect 19 43 21 46
rect 29 43 31 46
rect 19 41 31 43
rect 25 39 27 41
rect 29 39 31 41
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 25 33 31 39
rect 39 35 41 46
rect 49 35 51 38
rect 25 31 27 33
rect 29 31 31 33
rect 9 29 15 31
rect 19 29 31 31
rect 35 33 41 35
rect 35 31 37 33
rect 39 31 41 33
rect 35 29 41 31
rect 45 33 51 35
rect 45 31 47 33
rect 49 31 51 33
rect 59 31 61 38
rect 45 29 51 31
rect 55 29 70 31
rect 12 26 14 29
rect 19 26 21 29
rect 29 26 31 29
rect 36 26 38 29
rect 48 26 50 29
rect 55 26 57 29
rect 64 27 66 29
rect 68 27 70 29
rect 12 11 14 15
rect 19 11 21 15
rect 29 4 31 9
rect 36 4 38 9
rect 64 25 70 27
rect 48 2 50 6
rect 55 2 57 6
<< ndif >>
rect 3 15 12 26
rect 14 15 19 26
rect 21 19 29 26
rect 21 17 24 19
rect 26 17 29 19
rect 21 15 29 17
rect 3 7 10 15
rect 24 9 29 15
rect 31 9 36 26
rect 38 10 48 26
rect 38 9 42 10
rect 3 5 6 7
rect 8 5 10 7
rect 3 3 10 5
rect 40 8 42 9
rect 44 8 48 10
rect 40 6 48 8
rect 50 6 55 26
rect 57 19 62 26
rect 57 17 64 19
rect 57 15 60 17
rect 62 15 64 17
rect 57 13 64 15
rect 57 6 62 13
<< pdif >>
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 46 9 59
rect 11 57 19 63
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 46 19 48
rect 21 61 29 63
rect 21 59 24 61
rect 26 59 29 61
rect 21 46 29 59
rect 31 57 39 63
rect 31 55 34 57
rect 36 55 39 57
rect 31 50 39 55
rect 31 48 34 50
rect 36 48 39 50
rect 31 46 39 48
rect 41 61 49 63
rect 41 59 44 61
rect 46 59 49 61
rect 41 46 49 59
rect 43 38 49 46
rect 51 57 59 63
rect 51 55 54 57
rect 56 55 59 57
rect 51 50 59 55
rect 51 48 54 50
rect 56 48 59 50
rect 51 38 59 48
rect 61 61 69 63
rect 61 59 64 61
rect 66 59 69 61
rect 61 53 69 59
rect 61 51 64 53
rect 66 51 69 53
rect 61 38 69 51
<< alu1 >>
rect -2 64 74 72
rect 13 57 17 59
rect 33 57 38 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 51 17 55
rect 2 50 17 51
rect 33 55 34 57
rect 36 55 38 57
rect 33 50 38 55
rect 2 48 14 50
rect 16 48 34 50
rect 36 48 38 50
rect 2 46 38 48
rect 2 18 6 46
rect 17 41 31 42
rect 17 39 27 41
rect 29 39 31 41
rect 17 38 31 39
rect 25 33 31 38
rect 25 31 27 33
rect 29 31 31 33
rect 25 30 31 31
rect 50 37 62 43
rect 22 19 28 20
rect 22 18 24 19
rect 2 17 24 18
rect 26 17 28 19
rect 2 14 28 17
rect 50 21 54 37
rect 66 29 70 35
rect 68 27 70 29
rect 58 21 70 27
rect -2 7 74 8
rect -2 5 6 7
rect 8 5 16 7
rect 18 5 74 7
rect -2 0 74 5
<< ptie >>
rect 14 7 20 9
rect 14 5 16 7
rect 18 5 20 7
rect 14 3 20 5
<< nmos >>
rect 12 15 14 26
rect 19 15 21 26
rect 29 9 31 26
rect 36 9 38 26
rect 48 6 50 26
rect 55 6 57 26
<< pmos >>
rect 9 46 11 63
rect 19 46 21 63
rect 29 46 31 63
rect 39 46 41 63
rect 49 38 51 63
rect 59 38 61 63
<< polyct0 >>
rect 11 31 13 33
rect 37 31 39 33
rect 47 31 49 33
<< polyct1 >>
rect 27 39 29 41
rect 27 31 29 33
rect 66 27 68 29
<< ndifct0 >>
rect 42 8 44 10
rect 60 15 62 17
<< ndifct1 >>
rect 24 17 26 19
rect 6 5 8 7
<< ptiect1 >>
rect 16 5 18 7
<< pdifct0 >>
rect 4 59 6 61
rect 24 59 26 61
rect 44 59 46 61
rect 54 55 56 57
rect 54 48 56 50
rect 64 59 66 61
rect 64 51 66 53
<< pdifct1 >>
rect 14 55 16 57
rect 14 48 16 50
rect 34 55 36 57
rect 34 48 36 50
<< alu0 >>
rect 3 61 7 64
rect 3 59 4 61
rect 6 59 7 61
rect 23 61 27 64
rect 23 59 24 61
rect 26 59 27 61
rect 43 61 47 64
rect 43 59 44 61
rect 46 59 47 61
rect 63 61 67 64
rect 63 59 64 61
rect 66 59 67 61
rect 3 57 7 59
rect 23 57 27 59
rect 43 57 47 59
rect 53 57 57 59
rect 53 55 54 57
rect 56 55 57 57
rect 53 50 57 55
rect 42 48 54 50
rect 56 48 57 50
rect 63 53 67 59
rect 63 51 64 53
rect 66 51 67 53
rect 63 49 67 51
rect 42 46 57 48
rect 42 42 46 46
rect 10 33 14 35
rect 10 31 11 33
rect 13 31 14 33
rect 10 27 14 31
rect 36 38 46 42
rect 36 33 40 38
rect 36 31 37 33
rect 39 31 40 33
rect 36 27 40 31
rect 45 33 50 34
rect 45 31 47 33
rect 49 31 50 33
rect 45 30 50 31
rect 10 23 40 27
rect 36 18 40 23
rect 65 27 66 31
rect 36 17 64 18
rect 36 15 60 17
rect 62 15 64 17
rect 36 14 64 15
rect 40 10 46 11
rect 40 8 42 10
rect 44 8 46 10
<< labels >>
rlabel alu0 12 29 12 29 6 an
rlabel alu0 38 28 38 28 6 an
rlabel alu0 50 16 50 16 6 an
rlabel alu0 55 52 55 52 6 an
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 40 20 40 6 b
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel alu1 52 32 52 32 6 a1
rlabel alu1 36 56 36 56 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 24 60 24 6 a2
rlabel alu1 68 28 68 28 6 a2
rlabel alu1 60 40 60 40 6 a1
<< end >>
