magic
tech scmos
timestamp 1199203452
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 16 59 18 64
rect 26 59 28 64
rect 36 59 38 64
rect 48 59 50 64
rect 58 59 60 64
rect 16 43 18 46
rect 2 41 18 43
rect 2 39 4 41
rect 6 39 11 41
rect 2 37 11 39
rect 9 26 11 37
rect 26 35 28 38
rect 16 33 22 35
rect 16 31 18 33
rect 20 31 22 33
rect 16 29 22 31
rect 26 33 32 35
rect 26 31 28 33
rect 30 31 32 33
rect 26 29 32 31
rect 19 26 21 29
rect 26 26 28 29
rect 36 26 38 38
rect 48 35 50 38
rect 58 35 60 38
rect 46 33 53 35
rect 46 31 49 33
rect 51 31 53 33
rect 46 29 53 31
rect 57 33 63 35
rect 57 31 59 33
rect 61 31 63 33
rect 72 33 78 35
rect 72 31 74 33
rect 76 31 78 33
rect 57 29 63 31
rect 67 29 78 31
rect 46 26 48 29
rect 67 26 69 29
rect 9 8 11 13
rect 19 8 21 13
rect 26 8 28 13
rect 36 4 38 13
rect 46 8 48 13
rect 67 4 69 15
rect 36 2 69 4
<< ndif >>
rect 2 24 9 26
rect 2 22 4 24
rect 6 22 9 24
rect 2 17 9 22
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 11 17 19 26
rect 11 15 14 17
rect 16 15 19 17
rect 11 13 19 15
rect 21 13 26 26
rect 28 24 36 26
rect 28 22 31 24
rect 33 22 36 24
rect 28 13 36 22
rect 38 24 46 26
rect 38 22 41 24
rect 43 22 46 24
rect 38 13 46 22
rect 48 19 53 26
rect 48 17 55 19
rect 48 15 51 17
rect 53 15 55 17
rect 48 13 55 15
rect 59 17 67 26
rect 59 15 61 17
rect 63 15 67 17
rect 69 24 76 26
rect 69 22 72 24
rect 74 22 76 24
rect 69 20 76 22
rect 69 15 74 20
rect 59 13 65 15
<< pdif >>
rect 7 67 14 69
rect 7 65 10 67
rect 12 65 14 67
rect 7 59 14 65
rect 40 67 46 69
rect 40 65 42 67
rect 44 65 46 67
rect 40 59 46 65
rect 7 46 16 59
rect 18 57 26 59
rect 18 55 21 57
rect 23 55 26 57
rect 18 50 26 55
rect 18 48 21 50
rect 23 48 26 50
rect 18 46 26 48
rect 21 38 26 46
rect 28 49 36 59
rect 28 47 31 49
rect 33 47 36 49
rect 28 42 36 47
rect 28 40 31 42
rect 33 40 36 42
rect 28 38 36 40
rect 38 38 48 59
rect 50 42 58 59
rect 50 40 53 42
rect 55 40 58 42
rect 50 38 58 40
rect 60 57 67 59
rect 60 55 63 57
rect 65 55 67 57
rect 60 53 67 55
rect 60 38 65 53
<< alu1 >>
rect -2 67 82 72
rect -2 65 10 67
rect 12 65 42 67
rect 44 65 73 67
rect 75 65 82 67
rect -2 64 82 65
rect 2 54 15 59
rect 19 57 67 58
rect 19 55 21 57
rect 23 55 63 57
rect 65 55 67 57
rect 19 54 67 55
rect 2 41 6 54
rect 19 50 24 54
rect 10 48 21 50
rect 23 48 24 50
rect 10 46 24 48
rect 2 39 4 41
rect 2 29 6 39
rect 10 26 14 46
rect 10 24 35 26
rect 10 22 31 24
rect 33 22 35 24
rect 29 21 35 22
rect 48 33 54 35
rect 66 37 78 43
rect 48 31 49 33
rect 51 31 54 33
rect 48 29 54 31
rect 49 26 54 29
rect 49 22 63 26
rect 73 33 78 37
rect 73 31 74 33
rect 76 31 78 33
rect 73 29 78 31
rect -2 7 82 8
rect -2 5 73 7
rect 75 5 82 7
rect -2 0 82 5
<< ptie >>
rect 71 7 77 9
rect 71 5 73 7
rect 75 5 77 7
rect 71 3 77 5
<< ntie >>
rect 71 67 77 69
rect 71 65 73 67
rect 75 65 77 67
rect 71 40 77 65
<< nmos >>
rect 9 13 11 26
rect 19 13 21 26
rect 26 13 28 26
rect 36 13 38 26
rect 46 13 48 26
rect 67 15 69 26
<< pmos >>
rect 16 46 18 59
rect 26 38 28 59
rect 36 38 38 59
rect 48 38 50 59
rect 58 38 60 59
<< polyct0 >>
rect 18 31 20 33
rect 28 31 30 33
rect 59 31 61 33
<< polyct1 >>
rect 4 39 6 41
rect 49 31 51 33
rect 74 31 76 33
<< ndifct0 >>
rect 4 22 6 24
rect 4 15 6 17
rect 14 15 16 17
rect 41 22 43 24
rect 51 15 53 17
rect 61 15 63 17
rect 72 22 74 24
<< ndifct1 >>
rect 31 22 33 24
<< ntiect1 >>
rect 73 65 75 67
<< ptiect1 >>
rect 73 5 75 7
<< pdifct0 >>
rect 31 47 33 49
rect 31 40 33 42
rect 53 40 55 42
<< pdifct1 >>
rect 10 65 12 67
rect 42 65 44 67
rect 21 55 23 57
rect 21 48 23 50
rect 63 55 65 57
<< alu0 >>
rect 44 50 63 51
rect 29 49 63 50
rect 29 47 31 49
rect 33 47 63 49
rect 29 46 48 47
rect 6 37 7 43
rect 29 42 34 46
rect 52 42 56 44
rect 18 40 31 42
rect 33 40 34 42
rect 18 38 34 40
rect 39 40 53 42
rect 55 40 56 42
rect 39 38 56 40
rect 18 35 22 38
rect 17 33 22 35
rect 39 34 43 38
rect 17 31 18 33
rect 20 31 22 33
rect 17 29 22 31
rect 26 33 43 34
rect 26 31 28 33
rect 30 31 43 33
rect 26 30 43 31
rect 3 24 7 26
rect 3 22 4 24
rect 6 22 7 24
rect 3 17 7 22
rect 39 25 43 30
rect 59 34 63 47
rect 57 33 70 34
rect 57 31 59 33
rect 61 31 70 33
rect 57 30 70 31
rect 39 24 45 25
rect 39 22 41 24
rect 43 22 45 24
rect 66 25 70 30
rect 66 24 76 25
rect 66 22 72 24
rect 74 22 76 24
rect 39 21 45 22
rect 66 21 76 22
rect 3 15 4 17
rect 6 15 7 17
rect 3 8 7 15
rect 12 17 55 18
rect 12 15 14 17
rect 16 15 51 17
rect 53 15 55 17
rect 12 14 55 15
rect 59 17 65 18
rect 59 15 61 17
rect 63 15 65 17
rect 59 8 65 15
<< labels >>
rlabel alu0 20 35 20 35 6 a2n
rlabel alu0 31 44 31 44 6 a2n
rlabel alu0 34 32 34 32 6 a1n
rlabel alu0 41 31 41 31 6 a1n
rlabel alu0 47 40 47 40 6 a1n
rlabel alu0 63 32 63 32 6 a2n
rlabel alu0 71 23 71 23 6 a2n
rlabel alu1 12 36 12 36 6 z
rlabel alu1 4 44 4 44 6 b
rlabel alu1 12 56 12 56 6 b
rlabel alu1 20 24 20 24 6 z
rlabel alu1 28 24 28 24 6 z
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 52 28 52 28 6 a1
rlabel alu1 52 56 52 56 6 z
rlabel alu1 44 56 44 56 6 z
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 60 24 60 24 6 a1
rlabel alu1 76 36 76 36 6 a2
rlabel alu1 68 40 68 40 6 a2
rlabel alu1 60 56 60 56 6 z
<< end >>
