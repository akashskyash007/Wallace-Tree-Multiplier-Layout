magic
tech scmos
timestamp 1199202802
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 37 66 39 70
rect 49 66 51 70
rect 15 59 17 63
rect 25 59 27 63
rect 15 42 17 45
rect 25 42 27 45
rect 15 40 27 42
rect 17 38 19 40
rect 21 38 23 40
rect 17 36 23 38
rect 7 33 13 35
rect 7 31 9 33
rect 11 31 13 33
rect 7 29 14 31
rect 12 26 14 29
rect 19 26 21 36
rect 37 35 39 38
rect 33 33 39 35
rect 33 31 35 33
rect 37 31 39 33
rect 49 35 51 38
rect 49 33 55 35
rect 49 31 51 33
rect 53 31 55 33
rect 26 29 39 31
rect 26 26 28 29
rect 36 26 38 29
rect 43 26 45 31
rect 49 29 55 31
rect 50 26 52 29
rect 12 7 14 12
rect 19 4 21 12
rect 26 8 28 12
rect 36 8 38 12
rect 43 4 45 12
rect 50 7 52 12
rect 19 2 45 4
<< ndif >>
rect 2 23 12 26
rect 2 21 4 23
rect 6 21 12 23
rect 2 16 12 21
rect 2 14 4 16
rect 6 14 12 16
rect 2 12 12 14
rect 14 12 19 26
rect 21 12 26 26
rect 28 24 36 26
rect 28 22 31 24
rect 33 22 36 24
rect 28 12 36 22
rect 38 12 43 26
rect 45 12 50 26
rect 52 23 60 26
rect 52 21 55 23
rect 57 21 60 23
rect 52 16 60 21
rect 52 14 55 16
rect 57 14 60 16
rect 52 12 60 14
<< pdif >>
rect 29 64 37 66
rect 29 62 31 64
rect 33 62 37 64
rect 29 59 37 62
rect 6 57 15 59
rect 6 55 9 57
rect 11 55 15 57
rect 6 45 15 55
rect 17 57 25 59
rect 17 55 20 57
rect 22 55 25 57
rect 17 49 25 55
rect 17 47 20 49
rect 22 47 25 49
rect 17 45 25 47
rect 27 57 37 59
rect 27 55 31 57
rect 33 55 37 57
rect 27 45 37 55
rect 29 38 37 45
rect 39 57 49 66
rect 39 55 43 57
rect 45 55 49 57
rect 39 49 49 55
rect 39 47 43 49
rect 45 47 49 49
rect 39 38 49 47
rect 51 64 59 66
rect 51 62 54 64
rect 56 62 59 64
rect 51 57 59 62
rect 51 55 54 57
rect 56 55 59 57
rect 51 38 59 55
<< alu1 >>
rect -2 67 66 72
rect -2 65 5 67
rect 7 65 66 67
rect -2 64 66 65
rect 18 57 23 59
rect 18 55 20 57
rect 22 55 23 57
rect 9 42 14 51
rect 18 50 23 55
rect 41 57 47 58
rect 41 55 43 57
rect 45 55 47 57
rect 41 50 47 55
rect 18 49 47 50
rect 18 47 20 49
rect 22 47 43 49
rect 45 47 47 49
rect 18 46 47 47
rect 9 40 22 42
rect 9 38 19 40
rect 21 38 22 40
rect 7 33 14 34
rect 7 31 9 33
rect 11 31 14 33
rect 7 30 14 31
rect 10 18 14 30
rect 18 29 22 38
rect 26 22 30 46
rect 34 38 47 42
rect 34 33 38 38
rect 34 31 35 33
rect 37 31 38 33
rect 34 29 38 31
rect 42 33 55 34
rect 42 31 51 33
rect 53 31 55 33
rect 42 30 55 31
rect 42 18 46 30
rect 10 14 46 18
rect -2 0 66 8
<< ntie >>
rect 3 67 9 69
rect 3 65 5 67
rect 7 65 9 67
rect 3 63 9 65
<< nmos >>
rect 12 12 14 26
rect 19 12 21 26
rect 26 12 28 26
rect 36 12 38 26
rect 43 12 45 26
rect 50 12 52 26
<< pmos >>
rect 15 45 17 59
rect 25 45 27 59
rect 37 38 39 66
rect 49 38 51 66
<< polyct1 >>
rect 19 38 21 40
rect 9 31 11 33
rect 35 31 37 33
rect 51 31 53 33
<< ndifct0 >>
rect 4 21 6 23
rect 4 14 6 16
rect 31 22 33 24
rect 55 21 57 23
rect 55 14 57 16
<< ntiect1 >>
rect 5 65 7 67
<< pdifct0 >>
rect 31 62 33 64
rect 9 55 11 57
rect 31 55 33 57
rect 54 62 56 64
rect 54 55 56 57
<< pdifct1 >>
rect 20 55 22 57
rect 20 47 22 49
rect 43 55 45 57
rect 43 47 45 49
<< alu0 >>
rect 7 57 13 64
rect 29 62 31 64
rect 33 62 35 64
rect 7 55 9 57
rect 11 55 13 57
rect 7 54 13 55
rect 29 57 35 62
rect 52 62 54 64
rect 56 62 58 64
rect 29 55 31 57
rect 33 55 35 57
rect 29 54 35 55
rect 52 57 58 62
rect 52 55 54 57
rect 56 55 58 57
rect 52 54 58 55
rect 3 23 7 25
rect 3 21 4 23
rect 6 21 7 23
rect 3 16 7 21
rect 3 14 4 16
rect 6 14 7 16
rect 30 24 35 25
rect 30 22 31 24
rect 33 22 35 24
rect 26 21 35 22
rect 54 23 58 25
rect 54 21 55 23
rect 57 21 58 23
rect 54 16 58 21
rect 54 14 55 16
rect 57 14 58 16
rect 3 8 7 14
rect 54 8 58 14
<< labels >>
rlabel alu1 12 24 12 24 6 a
rlabel alu1 12 44 12 44 6 b
rlabel alu1 20 16 20 16 6 a
rlabel alu1 28 16 28 16 6 a
rlabel alu1 20 32 20 32 6 b
rlabel alu1 28 40 28 40 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 36 16 36 16 6 a
rlabel polyct1 36 32 36 32 6 c
rlabel alu1 44 24 44 24 6 a
rlabel alu1 44 40 44 40 6 c
rlabel alu1 36 48 36 48 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 32 68 32 68 6 vdd
rlabel polyct1 52 32 52 32 6 a
<< end >>
