magic
tech scmos
timestamp 1199470138
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -5 48 65 105
<< pwell >>
rect -5 -5 65 48
<< poly >>
rect 23 94 25 98
rect 31 94 33 98
rect 39 94 41 98
rect 47 94 49 98
rect 23 52 25 55
rect 19 50 25 52
rect 19 48 21 50
rect 23 48 25 50
rect 11 46 25 48
rect 11 23 13 46
rect 31 43 33 55
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 23 37 35 39
rect 23 23 25 37
rect 39 33 41 55
rect 47 52 49 55
rect 47 50 53 52
rect 47 48 49 50
rect 51 48 53 50
rect 47 46 53 48
rect 35 31 43 33
rect 35 29 39 31
rect 41 29 43 31
rect 35 27 43 29
rect 35 23 37 27
rect 47 23 49 46
rect 11 12 13 17
rect 23 12 25 17
rect 35 12 37 17
rect 47 12 49 17
<< ndif >>
rect 3 17 11 23
rect 13 21 23 23
rect 13 19 17 21
rect 19 19 23 21
rect 13 17 23 19
rect 25 17 35 23
rect 37 21 47 23
rect 37 19 41 21
rect 43 19 47 21
rect 37 17 47 19
rect 49 21 57 23
rect 49 19 53 21
rect 55 19 57 21
rect 49 17 57 19
rect 3 11 9 17
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 27 11 33 17
rect 27 9 29 11
rect 31 9 33 11
rect 27 7 33 9
<< pdif >>
rect 18 73 23 94
rect 15 71 23 73
rect 15 69 17 71
rect 19 69 23 71
rect 15 61 23 69
rect 15 59 17 61
rect 19 59 23 61
rect 15 57 23 59
rect 18 55 23 57
rect 25 55 31 94
rect 33 55 39 94
rect 41 55 47 94
rect 49 91 57 94
rect 49 89 53 91
rect 55 89 57 91
rect 49 81 57 89
rect 49 79 53 81
rect 55 79 57 81
rect 49 55 57 79
<< alu1 >>
rect -2 95 62 100
rect -2 93 5 95
rect 7 93 62 95
rect -2 91 62 93
rect -2 89 53 91
rect 55 89 62 91
rect -2 88 62 89
rect 52 81 56 88
rect 52 79 53 81
rect 55 79 56 81
rect 52 77 56 79
rect 16 71 22 73
rect 16 69 17 71
rect 19 69 22 71
rect 16 63 22 69
rect 37 68 53 72
rect 8 61 22 63
rect 8 59 17 61
rect 19 59 22 61
rect 8 57 22 59
rect 8 22 12 57
rect 28 53 32 63
rect 18 50 32 53
rect 18 48 21 50
rect 23 48 32 50
rect 18 47 32 48
rect 18 37 22 47
rect 38 43 42 53
rect 47 50 53 68
rect 47 48 49 50
rect 51 48 53 50
rect 47 47 53 48
rect 28 41 42 43
rect 28 39 31 41
rect 33 39 42 41
rect 28 37 42 39
rect 28 27 32 37
rect 48 32 52 43
rect 37 31 52 32
rect 37 29 39 31
rect 41 29 52 31
rect 37 27 52 29
rect 8 21 45 22
rect 8 19 17 21
rect 19 19 41 21
rect 43 19 45 21
rect 8 17 45 19
rect 52 21 56 23
rect 52 19 53 21
rect 55 19 56 21
rect 52 12 56 19
rect -2 11 62 12
rect -2 9 5 11
rect 7 9 29 11
rect 31 9 62 11
rect -2 7 62 9
rect -2 5 41 7
rect 43 5 51 7
rect 53 5 62 7
rect -2 0 62 5
<< ptie >>
rect 39 7 55 9
rect 39 5 41 7
rect 43 5 51 7
rect 53 5 55 7
rect 39 3 55 5
<< ntie >>
rect 3 95 9 97
rect 3 93 5 95
rect 7 93 9 95
rect 3 91 9 93
<< nmos >>
rect 11 17 13 23
rect 23 17 25 23
rect 35 17 37 23
rect 47 17 49 23
<< pmos >>
rect 23 55 25 94
rect 31 55 33 94
rect 39 55 41 94
rect 47 55 49 94
<< polyct1 >>
rect 21 48 23 50
rect 31 39 33 41
rect 49 48 51 50
rect 39 29 41 31
<< ndifct1 >>
rect 17 19 19 21
rect 41 19 43 21
rect 53 19 55 21
rect 5 9 7 11
rect 29 9 31 11
<< ntiect1 >>
rect 5 93 7 95
<< ptiect1 >>
rect 41 5 43 7
rect 51 5 53 7
<< pdifct1 >>
rect 17 69 19 71
rect 17 59 19 61
rect 53 89 55 91
rect 53 79 55 81
<< labels >>
rlabel alu1 10 40 10 40 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 20 45 20 45 6 d
rlabel alu1 20 65 20 65 6 z
rlabel alu1 30 20 30 20 6 z
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 40 20 40 20 6 z
rlabel alu1 30 35 30 35 6 c
rlabel alu1 40 45 40 45 6 c
rlabel polyct1 40 30 40 30 6 b
rlabel alu1 30 55 30 55 6 d
rlabel alu1 40 70 40 70 6 a
rlabel alu1 30 94 30 94 6 vdd
rlabel alu1 50 35 50 35 6 b
rlabel alu1 50 60 50 60 6 a
<< end >>
