magic
tech scmos
timestamp 1199203695
<< ab >>
rect 0 0 168 80
<< nwell >>
rect -5 36 173 88
<< pwell >>
rect -5 -8 173 36
<< poly >>
rect 11 70 13 74
rect 19 70 21 74
rect 27 70 29 74
rect 37 70 39 74
rect 44 70 46 74
rect 54 70 56 74
rect 75 70 77 74
rect 104 70 106 74
rect 114 70 116 74
rect 121 70 123 74
rect 131 70 133 74
rect 139 70 141 74
rect 147 70 149 74
rect 86 46 92 48
rect 86 44 88 46
rect 90 44 92 46
rect 86 42 92 44
rect 159 47 165 49
rect 159 45 161 47
rect 163 45 165 47
rect 159 43 165 45
rect 11 39 13 42
rect 19 39 21 42
rect 27 39 29 42
rect 37 39 39 42
rect 44 39 46 42
rect 54 39 56 42
rect 75 39 77 42
rect 86 39 88 42
rect 2 37 13 39
rect 2 35 4 37
rect 6 35 13 37
rect 2 33 13 35
rect 17 37 23 39
rect 17 35 19 37
rect 21 35 23 37
rect 17 33 23 35
rect 27 37 40 39
rect 27 35 36 37
rect 38 35 40 37
rect 44 36 48 39
rect 54 36 58 39
rect 27 33 40 35
rect 11 30 13 33
rect 19 30 21 33
rect 27 30 29 33
rect 37 30 39 33
rect 46 32 48 36
rect 46 30 52 32
rect 46 28 48 30
rect 50 28 52 30
rect 46 26 52 28
rect 46 23 48 26
rect 56 23 58 36
rect 62 37 77 39
rect 62 35 64 37
rect 66 35 77 37
rect 62 33 77 35
rect 83 37 88 39
rect 104 38 106 42
rect 68 30 70 33
rect 11 11 13 16
rect 19 11 21 16
rect 27 11 29 16
rect 37 11 39 16
rect 83 22 85 37
rect 92 36 106 38
rect 92 34 94 36
rect 96 34 106 36
rect 92 32 106 34
rect 104 29 106 32
rect 114 29 116 42
rect 121 39 123 42
rect 131 39 133 42
rect 139 39 141 42
rect 147 39 149 42
rect 159 39 161 43
rect 121 37 133 39
rect 121 35 123 37
rect 125 35 133 37
rect 121 33 133 35
rect 137 37 143 39
rect 137 35 139 37
rect 141 35 143 37
rect 137 33 143 35
rect 147 37 161 39
rect 121 29 123 33
rect 131 29 133 33
rect 139 29 141 33
rect 147 29 149 37
rect 79 20 85 22
rect 79 18 81 20
rect 83 18 85 20
rect 79 16 85 18
rect 160 21 166 23
rect 160 19 162 21
rect 164 19 166 21
rect 160 17 166 19
rect 68 12 70 16
rect 104 12 106 16
rect 46 6 48 11
rect 56 8 58 11
rect 114 8 116 16
rect 121 12 123 16
rect 131 12 133 16
rect 139 12 141 16
rect 147 12 149 16
rect 160 8 162 17
rect 56 6 162 8
<< ndif >>
rect 3 16 11 30
rect 13 16 19 30
rect 21 16 27 30
rect 29 28 37 30
rect 29 26 32 28
rect 34 26 37 28
rect 29 16 37 26
rect 39 23 44 30
rect 60 23 68 30
rect 39 16 46 23
rect 3 11 9 16
rect 41 11 46 16
rect 48 20 56 23
rect 48 18 51 20
rect 53 18 56 20
rect 48 11 56 18
rect 58 22 68 23
rect 58 20 62 22
rect 64 20 68 22
rect 58 16 68 20
rect 70 22 75 30
rect 70 20 77 22
rect 70 18 73 20
rect 75 18 77 20
rect 70 16 77 18
rect 97 20 104 29
rect 97 18 99 20
rect 101 18 104 20
rect 97 16 104 18
rect 106 27 114 29
rect 106 25 109 27
rect 111 25 114 27
rect 106 20 114 25
rect 106 18 109 20
rect 111 18 114 20
rect 106 16 114 18
rect 116 16 121 29
rect 123 21 131 29
rect 123 19 126 21
rect 128 19 131 21
rect 123 16 131 19
rect 133 16 139 29
rect 141 16 147 29
rect 149 27 158 29
rect 149 25 154 27
rect 156 25 158 27
rect 149 20 158 25
rect 149 18 154 20
rect 156 18 158 20
rect 149 16 158 18
rect 58 15 66 16
rect 58 13 62 15
rect 64 13 66 15
rect 58 11 66 13
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
<< pdif >>
rect 3 68 11 70
rect 3 66 6 68
rect 8 66 11 68
rect 3 42 11 66
rect 13 42 19 70
rect 21 42 27 70
rect 29 53 37 70
rect 29 51 32 53
rect 34 51 37 53
rect 29 42 37 51
rect 39 42 44 70
rect 46 61 54 70
rect 46 59 49 61
rect 51 59 54 61
rect 46 42 54 59
rect 56 68 75 70
rect 56 66 60 68
rect 62 66 70 68
rect 72 66 75 68
rect 56 42 75 66
rect 77 48 82 70
rect 97 68 104 70
rect 97 66 99 68
rect 101 66 104 68
rect 77 46 84 48
rect 77 44 80 46
rect 82 44 84 46
rect 77 42 84 44
rect 97 42 104 66
rect 106 46 114 70
rect 106 44 109 46
rect 111 44 114 46
rect 106 42 114 44
rect 116 42 121 70
rect 123 53 131 70
rect 123 51 126 53
rect 128 51 131 53
rect 123 42 131 51
rect 133 42 139 70
rect 141 42 147 70
rect 149 63 155 70
rect 149 61 157 63
rect 149 59 152 61
rect 154 59 157 61
rect 149 42 157 59
<< alu1 >>
rect -2 81 170 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 170 81
rect -2 68 170 79
rect 10 53 141 54
rect 10 51 32 53
rect 34 51 126 53
rect 128 51 141 53
rect 10 50 141 51
rect 10 29 14 50
rect 25 42 73 46
rect 25 39 30 42
rect 18 37 30 39
rect 137 46 141 50
rect 137 42 150 46
rect 18 35 19 37
rect 21 35 30 37
rect 18 33 30 35
rect 34 37 68 38
rect 34 35 36 37
rect 38 35 64 37
rect 66 35 68 37
rect 34 34 68 35
rect 73 36 97 38
rect 73 34 94 36
rect 96 34 97 36
rect 93 32 97 34
rect 10 28 36 29
rect 10 26 32 28
rect 34 26 36 28
rect 10 25 36 26
rect 146 22 150 42
rect 154 33 166 39
rect 124 21 150 22
rect 124 19 126 21
rect 128 19 150 21
rect 124 18 150 19
rect 161 21 166 33
rect 161 19 162 21
rect 164 19 166 21
rect 161 17 166 19
rect -2 11 170 12
rect -2 9 5 11
rect 7 9 170 11
rect -2 1 170 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 170 1
rect -2 -2 170 -1
<< ptie >>
rect 0 1 168 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 115 1
rect 117 -1 123 1
rect 125 -1 131 1
rect 133 -1 139 1
rect 141 -1 147 1
rect 149 -1 155 1
rect 157 -1 163 1
rect 165 -1 168 1
rect 0 -3 168 -1
<< ntie >>
rect 0 81 168 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 115 81
rect 117 79 123 81
rect 125 79 131 81
rect 133 79 139 81
rect 141 79 147 81
rect 149 79 155 81
rect 157 79 163 81
rect 165 79 168 81
rect 0 77 168 79
<< nmos >>
rect 11 16 13 30
rect 19 16 21 30
rect 27 16 29 30
rect 37 16 39 30
rect 46 11 48 23
rect 56 11 58 23
rect 68 16 70 30
rect 104 16 106 29
rect 114 16 116 29
rect 121 16 123 29
rect 131 16 133 29
rect 139 16 141 29
rect 147 16 149 29
<< pmos >>
rect 11 42 13 70
rect 19 42 21 70
rect 27 42 29 70
rect 37 42 39 70
rect 44 42 46 70
rect 54 42 56 70
rect 75 42 77 70
rect 104 42 106 70
rect 114 42 116 70
rect 121 42 123 70
rect 131 42 133 70
rect 139 42 141 70
rect 147 42 149 70
<< polyct0 >>
rect 88 44 90 46
rect 161 45 163 47
rect 4 35 6 37
rect 48 28 50 30
rect 123 35 125 37
rect 139 35 141 37
rect 81 18 83 20
<< polyct1 >>
rect 19 35 21 37
rect 36 35 38 37
rect 64 35 66 37
rect 94 34 96 36
rect 162 19 164 21
<< ndifct0 >>
rect 51 18 53 20
rect 62 20 64 22
rect 73 18 75 20
rect 99 18 101 20
rect 109 25 111 27
rect 109 18 111 20
rect 154 25 156 27
rect 154 18 156 20
rect 62 13 64 15
<< ndifct1 >>
rect 32 26 34 28
rect 126 19 128 21
rect 5 9 7 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
rect 115 79 117 81
rect 123 79 125 81
rect 131 79 133 81
rect 139 79 141 81
rect 147 79 149 81
rect 155 79 157 81
rect 163 79 165 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
rect 115 -1 117 1
rect 123 -1 125 1
rect 131 -1 133 1
rect 139 -1 141 1
rect 147 -1 149 1
rect 155 -1 157 1
rect 163 -1 165 1
<< pdifct0 >>
rect 6 66 8 68
rect 49 59 51 61
rect 60 66 62 68
rect 70 66 72 68
rect 99 66 101 68
rect 80 44 82 46
rect 109 44 111 46
rect 152 59 154 61
<< pdifct1 >>
rect 32 51 34 53
rect 126 51 128 53
<< alu0 >>
rect 4 66 6 68
rect 8 66 10 68
rect 4 65 10 66
rect 58 66 60 68
rect 62 66 70 68
rect 72 66 74 68
rect 58 65 74 66
rect 97 66 99 68
rect 101 66 103 68
rect 97 65 103 66
rect 3 61 148 62
rect 3 59 49 61
rect 51 59 148 61
rect 3 58 148 59
rect 3 37 7 58
rect 144 54 148 58
rect 151 61 155 68
rect 151 59 152 61
rect 154 59 155 61
rect 151 57 155 59
rect 3 35 4 37
rect 6 35 7 37
rect 3 21 7 35
rect 144 50 164 54
rect 78 46 104 47
rect 73 42 75 46
rect 78 44 80 46
rect 82 44 88 46
rect 90 44 104 46
rect 78 43 104 44
rect 71 38 75 42
rect 100 38 104 43
rect 107 46 113 47
rect 160 47 164 50
rect 107 44 109 46
rect 111 44 134 46
rect 107 42 134 44
rect 160 45 161 47
rect 163 45 164 47
rect 160 43 164 45
rect 130 38 134 42
rect 71 34 73 38
rect 100 37 127 38
rect 100 35 123 37
rect 125 35 127 37
rect 100 34 127 35
rect 130 37 143 38
rect 130 35 139 37
rect 141 35 143 37
rect 130 34 143 35
rect 46 30 52 31
rect 130 30 134 34
rect 46 28 48 30
rect 50 29 89 30
rect 107 29 134 30
rect 50 28 134 29
rect 46 27 134 28
rect 46 26 109 27
rect 85 25 109 26
rect 111 26 134 27
rect 111 25 113 26
rect 60 22 66 23
rect 3 20 55 21
rect 3 18 51 20
rect 53 18 55 20
rect 3 17 55 18
rect 60 20 62 22
rect 64 20 66 22
rect 60 15 66 20
rect 71 20 85 21
rect 71 18 73 20
rect 75 18 81 20
rect 83 18 85 20
rect 71 17 85 18
rect 97 20 103 21
rect 97 18 99 20
rect 101 18 103 20
rect 60 13 62 15
rect 64 13 66 15
rect 60 12 66 13
rect 88 12 92 16
rect 97 12 103 18
rect 107 20 113 25
rect 107 18 109 20
rect 111 18 113 20
rect 153 27 157 29
rect 153 25 154 27
rect 156 25 157 27
rect 153 20 157 25
rect 153 18 154 20
rect 156 18 157 20
rect 107 17 113 18
rect 153 12 157 18
<< labels >>
rlabel alu0 5 39 5 39 6 an
rlabel alu0 29 19 29 19 6 an
rlabel alu0 67 28 67 28 6 bn
rlabel alu0 78 19 78 19 6 cn
rlabel alu0 110 23 110 23 6 bn
rlabel alu0 113 36 113 36 6 cn
rlabel alu0 91 45 91 45 6 cn
rlabel alu0 120 44 120 44 6 bn
rlabel alu0 136 36 136 36 6 bn
rlabel alu0 162 48 162 48 6 an
rlabel alu0 75 60 75 60 6 an
rlabel polyct1 20 36 20 36 6 b
rlabel alu1 28 40 28 40 6 b
rlabel alu1 12 36 12 36 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 44 36 44 6 b
rlabel alu1 44 36 44 36 6 c
rlabel alu1 44 44 44 44 6 b
rlabel alu1 52 36 52 36 6 c
rlabel alu1 52 44 52 44 6 b
rlabel alu1 60 36 60 36 6 c
rlabel alu1 60 44 60 44 6 b
rlabel alu1 36 52 36 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 60 52 60 52 6 z
rlabel alu1 84 6 84 6 6 vss
rlabel alu1 68 44 68 44 6 b
rlabel alu1 76 36 76 36 6 b
rlabel alu1 84 36 84 36 6 b
rlabel alu1 92 36 92 36 6 b
rlabel alu1 76 52 76 52 6 z
rlabel alu1 84 52 84 52 6 z
rlabel alu1 92 52 92 52 6 z
rlabel alu1 68 52 68 52 6 z
rlabel alu1 84 74 84 74 6 vdd
rlabel alu1 132 20 132 20 6 z
rlabel alu1 108 52 108 52 6 z
rlabel alu1 116 52 116 52 6 z
rlabel alu1 124 52 124 52 6 z
rlabel alu1 132 52 132 52 6 z
rlabel alu1 100 52 100 52 6 z
rlabel alu1 164 28 164 28 6 a
rlabel alu1 140 20 140 20 6 z
rlabel alu1 148 32 148 32 6 z
rlabel alu1 140 44 140 44 6 z
rlabel alu1 156 36 156 36 6 a
<< end >>
