magic
tech scmos
timestamp 1199202645
<< ab >>
rect 0 0 48 80
<< nwell >>
rect -5 36 53 88
<< pwell >>
rect -5 -8 53 36
<< poly >>
rect 9 66 11 71
rect 19 66 21 71
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 32 39
rect 19 35 27 37
rect 29 35 32 37
rect 40 37 46 39
rect 40 35 42 37
rect 44 35 46 37
rect 19 33 32 35
rect 13 30 15 33
rect 20 30 22 33
rect 30 30 32 33
rect 37 33 46 35
rect 37 30 39 33
rect 13 6 15 10
rect 20 6 22 10
rect 30 6 32 10
rect 37 6 39 10
<< ndif >>
rect 5 14 13 30
rect 5 12 8 14
rect 10 12 13 14
rect 5 10 13 12
rect 15 10 20 30
rect 22 21 30 30
rect 22 19 25 21
rect 27 19 30 21
rect 22 10 30 19
rect 32 10 37 30
rect 39 21 46 30
rect 39 19 42 21
rect 44 19 46 21
rect 39 14 46 19
rect 39 12 42 14
rect 44 12 46 14
rect 39 10 46 12
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 56 9 62
rect 2 54 4 56
rect 6 54 9 56
rect 2 42 9 54
rect 11 53 19 66
rect 11 51 14 53
rect 16 51 19 53
rect 11 46 19 51
rect 11 44 14 46
rect 16 44 19 46
rect 11 42 19 44
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 56 29 62
rect 21 54 24 56
rect 26 54 29 56
rect 21 42 29 54
<< alu1 >>
rect -2 81 50 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 50 81
rect -2 68 50 79
rect 12 53 18 54
rect 12 51 14 53
rect 16 51 18 53
rect 12 47 18 51
rect 2 46 18 47
rect 2 44 14 46
rect 16 44 18 46
rect 2 43 18 44
rect 2 22 6 43
rect 25 42 39 46
rect 10 37 19 39
rect 10 35 11 37
rect 13 35 19 37
rect 10 33 19 35
rect 25 37 31 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 40 37 46 38
rect 40 35 42 37
rect 44 35 46 37
rect 15 30 19 33
rect 40 30 46 35
rect 15 26 46 30
rect 2 21 31 22
rect 2 19 25 21
rect 27 19 31 21
rect 2 18 31 19
rect -2 1 50 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 50 1
rect -2 -2 50 -1
<< ptie >>
rect 0 1 48 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 48 1
rect 0 -3 48 -1
<< ntie >>
rect 0 81 48 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 48 81
rect 0 77 48 79
<< nmos >>
rect 13 10 15 30
rect 20 10 22 30
rect 30 10 32 30
rect 37 10 39 30
<< pmos >>
rect 9 42 11 66
rect 19 42 21 66
<< polyct1 >>
rect 11 35 13 37
rect 27 35 29 37
rect 42 35 44 37
<< ndifct0 >>
rect 8 12 10 14
rect 42 19 44 21
rect 42 12 44 14
<< ndifct1 >>
rect 25 19 27 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
<< pdifct0 >>
rect 4 62 6 64
rect 4 54 6 56
rect 24 62 26 64
rect 24 54 26 56
<< pdifct1 >>
rect 14 51 16 53
rect 14 44 16 46
<< alu0 >>
rect 3 64 7 68
rect 3 62 4 64
rect 6 62 7 64
rect 3 56 7 62
rect 3 54 4 56
rect 6 54 7 56
rect 23 64 27 68
rect 23 62 24 64
rect 26 62 27 64
rect 23 56 27 62
rect 23 54 24 56
rect 26 54 27 56
rect 3 52 7 54
rect 23 52 27 54
rect 40 21 46 22
rect 40 19 42 21
rect 44 19 46 21
rect 6 14 12 15
rect 6 12 8 14
rect 10 12 12 14
rect 40 14 46 19
rect 40 12 42 14
rect 44 12 46 14
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 12 20 12 20 6 z
rlabel polyct1 12 36 12 36 6 a
rlabel alu1 20 28 20 28 6 a
rlabel alu1 24 6 24 6 6 vss
rlabel alu1 28 20 28 20 6 z
rlabel alu1 28 28 28 28 6 a
rlabel alu1 28 40 28 40 6 b
rlabel alu1 24 74 24 74 6 vdd
rlabel alu1 36 28 36 28 6 a
rlabel alu1 36 44 36 44 6 b
<< end >>
