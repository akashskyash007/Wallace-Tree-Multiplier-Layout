magic
tech scmos
timestamp 1199543664
<< ab >>
rect 0 0 110 100
<< nwell >>
rect -2 48 112 104
<< pwell >>
rect -2 -4 112 48
<< poly >>
rect 35 95 37 98
rect 47 95 49 98
rect 57 95 59 98
rect 81 95 83 98
rect 93 95 95 98
rect 11 84 13 87
rect 23 84 25 87
rect 11 43 13 55
rect 23 53 25 55
rect 35 53 37 55
rect 21 51 25 53
rect 33 51 37 53
rect 21 43 23 51
rect 33 43 35 51
rect 7 41 13 43
rect 7 39 9 41
rect 11 39 13 41
rect 7 37 13 39
rect 17 41 23 43
rect 17 39 19 41
rect 21 39 23 41
rect 17 37 23 39
rect 27 41 35 43
rect 27 39 29 41
rect 31 39 35 41
rect 47 43 49 55
rect 57 43 59 55
rect 81 53 83 55
rect 93 53 95 55
rect 75 51 95 53
rect 75 49 77 51
rect 79 49 95 51
rect 75 47 95 49
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 27 37 35 39
rect 11 35 13 37
rect 21 35 23 37
rect 33 35 35 37
rect 45 37 53 39
rect 57 41 63 43
rect 57 39 59 41
rect 61 39 63 41
rect 57 37 63 39
rect 45 35 47 37
rect 57 35 59 37
rect 81 35 83 47
rect 93 35 95 47
rect 33 20 35 23
rect 45 20 47 23
rect 11 14 13 17
rect 21 14 23 17
rect 57 20 59 23
rect 81 12 83 15
rect 93 12 95 15
<< ndif >>
rect 3 17 11 35
rect 13 17 21 35
rect 23 23 33 35
rect 35 23 45 35
rect 47 23 57 35
rect 59 23 67 35
rect 23 21 31 23
rect 23 19 27 21
rect 29 19 31 21
rect 37 21 43 23
rect 23 17 31 19
rect 37 19 39 21
rect 41 19 43 21
rect 37 17 43 19
rect 3 11 9 17
rect 49 11 55 23
rect 61 21 67 23
rect 61 19 63 21
rect 65 19 67 21
rect 61 17 67 19
rect 73 31 81 35
rect 73 29 75 31
rect 77 29 81 31
rect 73 21 81 29
rect 73 19 75 21
rect 77 19 81 21
rect 73 15 81 19
rect 83 31 93 35
rect 83 29 87 31
rect 89 29 93 31
rect 83 21 93 29
rect 83 19 87 21
rect 89 19 93 21
rect 83 15 93 19
rect 95 31 103 35
rect 95 29 99 31
rect 101 29 103 31
rect 95 21 103 29
rect 95 19 99 21
rect 101 19 103 21
rect 95 15 103 19
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 49 9 51 11
rect 53 9 55 11
rect 49 7 55 9
<< pdif >>
rect 15 91 21 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 84 21 89
rect 28 84 35 95
rect 3 81 11 84
rect 3 79 5 81
rect 7 79 11 81
rect 3 55 11 79
rect 13 55 23 84
rect 25 81 35 84
rect 25 79 29 81
rect 31 79 35 81
rect 25 55 35 79
rect 37 71 47 95
rect 37 69 41 71
rect 43 69 47 71
rect 37 55 47 69
rect 49 55 57 95
rect 59 81 67 95
rect 59 79 63 81
rect 65 79 67 81
rect 59 55 67 79
rect 73 91 81 95
rect 73 89 75 91
rect 77 89 81 91
rect 73 81 81 89
rect 73 79 75 81
rect 77 79 81 81
rect 73 55 81 79
rect 83 81 93 95
rect 83 79 87 81
rect 89 79 93 81
rect 83 71 93 79
rect 83 69 87 71
rect 89 69 93 71
rect 83 61 93 69
rect 83 59 87 61
rect 89 59 93 61
rect 83 55 93 59
rect 95 91 103 95
rect 95 89 99 91
rect 101 89 103 91
rect 95 81 103 89
rect 95 79 99 81
rect 101 79 103 81
rect 95 71 103 79
rect 95 69 99 71
rect 101 69 103 71
rect 95 61 103 69
rect 95 59 99 61
rect 101 59 103 61
rect 95 55 103 59
<< alu1 >>
rect -2 91 112 100
rect -2 89 17 91
rect 19 89 75 91
rect 77 89 99 91
rect 101 89 112 91
rect -2 88 112 89
rect 4 81 8 82
rect 28 81 32 82
rect 62 81 66 82
rect 4 79 5 81
rect 7 79 29 81
rect 31 79 63 81
rect 65 79 66 81
rect 4 78 8 79
rect 28 78 32 79
rect 62 78 66 79
rect 74 81 78 88
rect 74 79 75 81
rect 77 79 78 81
rect 74 78 78 79
rect 86 81 92 82
rect 86 79 87 81
rect 89 79 92 81
rect 86 78 92 79
rect 88 72 92 78
rect 8 41 12 72
rect 8 39 9 41
rect 11 39 12 41
rect 8 18 12 39
rect 18 41 22 72
rect 18 39 19 41
rect 21 39 22 41
rect 18 28 22 39
rect 28 41 32 72
rect 40 71 44 72
rect 86 71 92 72
rect 28 39 29 41
rect 31 39 32 41
rect 28 38 32 39
rect 39 69 41 71
rect 43 69 79 71
rect 39 68 44 69
rect 39 31 41 68
rect 29 29 41 31
rect 48 41 52 62
rect 48 39 49 41
rect 51 39 52 41
rect 29 22 31 29
rect 48 28 52 39
rect 58 41 62 62
rect 77 52 79 69
rect 86 69 87 71
rect 89 69 92 71
rect 86 68 92 69
rect 88 62 92 68
rect 86 61 92 62
rect 86 59 87 61
rect 89 59 92 61
rect 86 58 92 59
rect 98 81 102 88
rect 98 79 99 81
rect 101 79 102 81
rect 98 71 102 79
rect 98 69 99 71
rect 101 69 102 71
rect 98 61 102 69
rect 98 59 99 61
rect 101 59 102 61
rect 98 58 102 59
rect 76 51 80 52
rect 76 49 77 51
rect 79 49 80 51
rect 76 48 80 49
rect 58 39 59 41
rect 61 39 62 41
rect 58 28 62 39
rect 88 32 92 58
rect 74 31 78 32
rect 74 29 75 31
rect 77 29 78 31
rect 26 21 31 22
rect 26 19 27 21
rect 29 19 31 21
rect 38 21 42 22
rect 62 21 66 22
rect 38 19 39 21
rect 41 19 63 21
rect 65 19 66 21
rect 26 18 30 19
rect 38 18 42 19
rect 62 18 66 19
rect 74 21 78 29
rect 86 31 92 32
rect 86 29 87 31
rect 89 29 92 31
rect 86 28 92 29
rect 88 22 92 28
rect 74 19 75 21
rect 77 19 78 21
rect 74 12 78 19
rect 86 21 92 22
rect 86 19 87 21
rect 89 19 92 21
rect 86 18 92 19
rect 98 31 102 32
rect 98 29 99 31
rect 101 29 102 31
rect 98 21 102 29
rect 98 19 99 21
rect 101 19 102 21
rect 98 12 102 19
rect -2 11 112 12
rect -2 9 5 11
rect 7 9 51 11
rect 53 9 112 11
rect -2 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 112 9
rect -2 5 63 7
rect 65 5 75 7
rect 77 5 87 7
rect 89 5 99 7
rect 101 5 112 7
rect -2 0 112 5
<< ptie >>
rect 21 9 43 11
rect 21 7 23 9
rect 25 7 31 9
rect 33 7 39 9
rect 41 7 43 9
rect 61 7 103 9
rect 21 5 43 7
rect 61 5 63 7
rect 65 5 75 7
rect 77 5 87 7
rect 89 5 99 7
rect 101 5 103 7
rect 61 3 103 5
<< nmos >>
rect 11 17 13 35
rect 21 17 23 35
rect 33 23 35 35
rect 45 23 47 35
rect 57 23 59 35
rect 81 15 83 35
rect 93 15 95 35
<< pmos >>
rect 11 55 13 84
rect 23 55 25 84
rect 35 55 37 95
rect 47 55 49 95
rect 57 55 59 95
rect 81 55 83 95
rect 93 55 95 95
<< polyct1 >>
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 77 49 79 51
rect 49 39 51 41
rect 59 39 61 41
<< ndifct1 >>
rect 27 19 29 21
rect 39 19 41 21
rect 63 19 65 21
rect 75 29 77 31
rect 75 19 77 21
rect 87 29 89 31
rect 87 19 89 21
rect 99 29 101 31
rect 99 19 101 21
rect 5 9 7 11
rect 51 9 53 11
<< ptiect1 >>
rect 23 7 25 9
rect 31 7 33 9
rect 39 7 41 9
rect 63 5 65 7
rect 75 5 77 7
rect 87 5 89 7
rect 99 5 101 7
<< pdifct1 >>
rect 17 89 19 91
rect 5 79 7 81
rect 29 79 31 81
rect 41 69 43 71
rect 63 79 65 81
rect 75 89 77 91
rect 75 79 77 81
rect 87 79 89 81
rect 87 69 89 71
rect 87 59 89 61
rect 99 89 101 91
rect 99 79 101 81
rect 99 69 101 71
rect 99 59 101 61
<< labels >>
rlabel alu1 10 45 10 45 6 i0
rlabel alu1 20 50 20 50 6 i1
rlabel alu1 30 55 30 55 6 i4
rlabel alu1 55 6 55 6 6 vss
rlabel alu1 50 45 50 45 6 i2
rlabel alu1 60 45 60 45 6 i3
rlabel alu1 55 94 55 94 6 vdd
rlabel alu1 90 50 90 50 6 q
<< end >>
