magic
tech scmos
timestamp 1199179204
<< ab >>
rect -715 0 17435 3960
<< alu1 >>
rect -660 3620 -440 3850
rect -660 3420 -650 3620
rect -450 3420 -440 3620
rect -660 2740 -440 3420
rect -660 2540 -650 2740
rect -450 2540 -440 2740
rect -660 1860 -440 2540
rect -660 1660 -650 1860
rect -450 1660 -440 1860
rect -660 980 -440 1660
rect -660 780 -650 980
rect -450 780 -440 980
rect -660 440 -440 780
rect 17160 440 17380 3850
rect -660 220 17380 440
rect -660 110 -440 220
rect 17160 110 17380 220
<< alu2 >>
rect -715 3620 17435 3630
rect -715 3420 -650 3620
rect -450 3420 17435 3620
rect -715 3410 17435 3420
rect -715 2740 17435 2750
rect -715 2540 -650 2740
rect -450 2540 17435 2740
rect -715 2530 17435 2540
rect -715 1860 17435 1870
rect -715 1660 -650 1860
rect -450 1660 17435 1860
rect -715 1650 17435 1660
rect -715 980 17435 990
rect -715 780 -650 980
rect -450 780 120 980
rect 320 780 1000 980
rect 1200 780 1880 980
rect 2080 780 2760 980
rect 2960 780 3640 980
rect 3840 780 4520 980
rect 4720 780 5400 980
rect 5600 780 6280 980
rect 6480 780 7160 980
rect 7360 780 8040 980
rect 8240 780 8920 980
rect 9120 780 9800 980
rect 10000 780 10680 980
rect 10880 780 11560 980
rect 11760 780 12440 980
rect 12640 780 13320 980
rect 13520 780 14200 980
rect 14400 780 15080 980
rect 15280 780 15960 980
rect 16160 780 16840 980
rect 17040 780 17435 980
rect -715 770 17435 780
<< alu3 >>
rect 110 3180 330 3850
rect 110 2980 120 3180
rect 320 2980 330 3180
rect 110 2300 330 2980
rect 110 2100 120 2300
rect 320 2100 330 2300
rect 110 1420 330 2100
rect 110 1220 120 1420
rect 320 1220 330 1420
rect 110 980 330 1220
rect 110 780 120 980
rect 320 780 330 980
rect 110 540 330 780
rect 110 340 120 540
rect 320 340 330 540
rect 110 110 330 340
rect 990 980 1210 3850
rect 990 780 1000 980
rect 1200 780 1210 980
rect 990 110 1210 780
rect 1870 980 2090 3850
rect 1870 780 1880 980
rect 2080 780 2090 980
rect 1870 110 2090 780
rect 2750 980 2970 3850
rect 2750 780 2760 980
rect 2960 780 2970 980
rect 2750 110 2970 780
rect 3630 980 3850 3850
rect 3630 780 3640 980
rect 3840 780 3850 980
rect 3630 110 3850 780
rect 4510 980 4730 3850
rect 4510 780 4520 980
rect 4720 780 4730 980
rect 4510 110 4730 780
rect 5390 980 5610 3850
rect 5390 780 5400 980
rect 5600 780 5610 980
rect 5390 110 5610 780
rect 6270 980 6490 3850
rect 6270 780 6280 980
rect 6480 780 6490 980
rect 6270 110 6490 780
rect 7150 980 7370 3850
rect 7150 780 7160 980
rect 7360 780 7370 980
rect 7150 110 7370 780
rect 8030 980 8250 3850
rect 8030 780 8040 980
rect 8240 780 8250 980
rect 8030 110 8250 780
rect 8910 980 9130 3850
rect 8910 780 8920 980
rect 9120 780 9130 980
rect 8910 110 9130 780
rect 9790 980 10010 3850
rect 9790 780 9800 980
rect 10000 780 10010 980
rect 9790 110 10010 780
rect 10670 980 10890 3850
rect 10670 780 10680 980
rect 10880 780 10890 980
rect 10670 110 10890 780
rect 11550 980 11770 3850
rect 11550 780 11560 980
rect 11760 780 11770 980
rect 11550 110 11770 780
rect 12430 980 12650 3850
rect 12430 780 12440 980
rect 12640 780 12650 980
rect 12430 110 12650 780
rect 13310 980 13530 3850
rect 13310 780 13320 980
rect 13520 780 13530 980
rect 13310 110 13530 780
rect 14190 980 14410 3850
rect 14190 780 14200 980
rect 14400 780 14410 980
rect 14190 110 14410 780
rect 15070 980 15290 3850
rect 15070 780 15080 980
rect 15280 780 15290 980
rect 15070 110 15290 780
rect 15950 980 16170 3850
rect 15950 780 15960 980
rect 16160 780 16170 980
rect 15950 110 16170 780
rect 16830 980 17050 3850
rect 16830 780 16840 980
rect 17040 780 17050 980
rect 16830 110 17050 780
<< alu4 >>
rect -715 3180 17435 3190
rect -715 2980 120 3180
rect 320 2980 17435 3180
rect -715 2970 17435 2980
rect -715 2300 17435 2310
rect -715 2100 120 2300
rect 320 2100 17435 2300
rect -715 2090 17435 2100
rect -715 1420 17435 1430
rect -715 1220 120 1420
rect 320 1220 17435 1420
rect -715 1210 17435 1220
rect -715 540 17435 550
rect -715 340 -320 540
rect -120 340 120 540
rect 320 340 560 540
rect 760 340 1440 540
rect 1640 340 2320 540
rect 2520 340 3200 540
rect 3400 340 4080 540
rect 4280 340 4960 540
rect 5160 340 5840 540
rect 6040 340 6720 540
rect 6920 340 7600 540
rect 7800 340 8480 540
rect 8680 340 9360 540
rect 9560 340 10240 540
rect 10440 340 11120 540
rect 11320 340 12000 540
rect 12200 340 12880 540
rect 13080 340 13760 540
rect 13960 340 14640 540
rect 14840 340 15520 540
rect 15720 340 16400 540
rect 16600 340 17435 540
rect -715 330 17435 340
<< alu5 >>
rect -330 540 -110 3850
rect -330 340 -320 540
rect -120 340 -110 540
rect -330 110 -110 340
rect 550 540 770 3850
rect 550 340 560 540
rect 760 340 770 540
rect 550 110 770 340
rect 1430 540 1650 3850
rect 1430 340 1440 540
rect 1640 340 1650 540
rect 1430 110 1650 340
rect 2310 540 2530 3850
rect 2310 340 2320 540
rect 2520 340 2530 540
rect 2310 110 2530 340
rect 3190 540 3410 3850
rect 3190 340 3200 540
rect 3400 340 3410 540
rect 3190 110 3410 340
rect 4070 540 4290 3850
rect 4070 340 4080 540
rect 4280 340 4290 540
rect 4070 110 4290 340
rect 4950 540 5170 3850
rect 4950 340 4960 540
rect 5160 340 5170 540
rect 4950 110 5170 340
rect 5830 540 6050 3850
rect 5830 340 5840 540
rect 6040 340 6050 540
rect 5830 110 6050 340
rect 6710 540 6930 3850
rect 6710 340 6720 540
rect 6920 340 6930 540
rect 6710 110 6930 340
rect 7590 540 7810 3850
rect 7590 340 7600 540
rect 7800 340 7810 540
rect 7590 110 7810 340
rect 8470 540 8690 3850
rect 8470 340 8480 540
rect 8680 340 8690 540
rect 8470 110 8690 340
rect 9350 540 9570 3850
rect 9350 340 9360 540
rect 9560 340 9570 540
rect 9350 110 9570 340
rect 10230 540 10450 3850
rect 10230 340 10240 540
rect 10440 340 10450 540
rect 10230 110 10450 340
rect 11110 540 11330 3850
rect 11110 340 11120 540
rect 11320 340 11330 540
rect 11110 110 11330 340
rect 11990 540 12210 3850
rect 11990 340 12000 540
rect 12200 340 12210 540
rect 11990 110 12210 340
rect 12870 540 13090 3850
rect 12870 340 12880 540
rect 13080 340 13090 540
rect 12870 110 13090 340
rect 13750 540 13970 3850
rect 13750 340 13760 540
rect 13960 340 13970 540
rect 13750 110 13970 340
rect 14630 540 14850 3850
rect 14630 340 14640 540
rect 14840 340 14850 540
rect 14630 110 14850 340
rect 15510 540 15730 3850
rect 15510 340 15520 540
rect 15720 340 15730 540
rect 15510 110 15730 340
rect 16390 540 16610 3850
rect 16390 340 16400 540
rect 16600 340 16610 540
rect 16390 110 16610 340
<< via1 >>
rect -650 3420 -450 3620
rect -650 2540 -450 2740
rect -650 1660 -450 1860
rect -650 780 -450 980
<< via2 >>
rect 120 780 320 980
rect 1000 780 1200 980
rect 1880 780 2080 980
rect 2760 780 2960 980
rect 3640 780 3840 980
rect 4520 780 4720 980
rect 5400 780 5600 980
rect 6280 780 6480 980
rect 7160 780 7360 980
rect 8040 780 8240 980
rect 8920 780 9120 980
rect 9800 780 10000 980
rect 10680 780 10880 980
rect 11560 780 11760 980
rect 12440 780 12640 980
rect 13320 780 13520 980
rect 14200 780 14400 980
rect 15080 780 15280 980
rect 15960 780 16160 980
rect 16840 780 17040 980
<< via3 >>
rect 120 2980 320 3180
rect 120 2100 320 2300
rect 120 1220 320 1420
rect 120 340 320 540
<< via4 >>
rect -320 340 -120 540
rect 560 340 760 540
rect 1440 340 1640 540
rect 2320 340 2520 540
rect 3200 340 3400 540
rect 4080 340 4280 540
rect 4960 340 5160 540
rect 5840 340 6040 540
rect 6720 340 6920 540
rect 7600 340 7800 540
rect 8480 340 8680 540
rect 9360 340 9560 540
rect 10240 340 10440 540
rect 11120 340 11320 540
rect 12000 340 12200 540
rect 12880 340 13080 540
rect 13760 340 13960 540
rect 14640 340 14840 540
rect 15520 340 15720 540
rect 16400 340 16600 540
<< end >>
