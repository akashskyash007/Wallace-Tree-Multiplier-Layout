magic
tech scmos
timestamp 1199202453
<< ab >>
rect 0 0 56 80
<< nwell >>
rect -5 36 61 88
<< pwell >>
rect -5 -8 61 36
<< poly >>
rect 10 70 12 74
rect 18 70 20 74
rect 28 70 30 74
rect 36 70 38 74
rect 48 62 54 64
rect 48 60 50 62
rect 52 60 54 62
rect 45 58 54 60
rect 45 55 47 58
rect 10 42 12 45
rect 18 42 20 45
rect 28 42 30 45
rect 36 42 38 45
rect 45 43 47 46
rect 9 39 12 42
rect 16 40 22 42
rect 9 31 11 39
rect 16 38 18 40
rect 20 38 22 40
rect 16 36 22 38
rect 26 40 32 42
rect 36 40 40 42
rect 45 41 50 43
rect 26 38 28 40
rect 30 38 32 40
rect 26 36 32 38
rect 38 37 40 40
rect 26 32 28 36
rect 38 35 44 37
rect 38 33 40 35
rect 42 33 44 35
rect 38 32 44 33
rect 2 29 11 31
rect 2 27 4 29
rect 6 27 11 29
rect 2 25 11 27
rect 9 22 11 25
rect 16 30 28 32
rect 35 31 44 32
rect 35 30 41 31
rect 16 22 18 30
rect 35 27 37 30
rect 48 27 50 41
rect 26 22 28 26
rect 45 25 50 27
rect 45 22 47 25
rect 35 12 37 16
rect 9 6 11 10
rect 16 6 18 10
rect 26 8 28 11
rect 45 8 47 16
rect 26 6 47 8
<< ndif >>
rect 30 22 35 27
rect 2 14 9 22
rect 2 12 4 14
rect 6 12 9 14
rect 2 10 9 12
rect 11 10 16 22
rect 18 20 26 22
rect 18 18 21 20
rect 23 18 26 20
rect 18 11 26 18
rect 28 16 35 22
rect 37 22 42 27
rect 37 20 45 22
rect 37 18 40 20
rect 42 18 45 20
rect 37 16 45 18
rect 47 20 54 22
rect 47 18 50 20
rect 52 18 54 20
rect 47 16 54 18
rect 28 11 33 16
rect 18 10 23 11
<< pdif >>
rect 2 68 10 70
rect 2 66 4 68
rect 6 66 10 68
rect 2 61 10 66
rect 2 59 4 61
rect 6 59 10 61
rect 2 45 10 59
rect 12 45 18 70
rect 20 61 28 70
rect 20 59 23 61
rect 25 59 28 61
rect 20 45 28 59
rect 30 45 36 70
rect 38 68 45 70
rect 38 66 41 68
rect 43 66 45 68
rect 38 63 45 66
rect 38 55 43 63
rect 38 46 45 55
rect 47 53 54 55
rect 47 51 50 53
rect 52 51 54 53
rect 47 49 54 51
rect 47 46 52 49
rect 38 45 43 46
<< alu1 >>
rect -2 81 58 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 58 81
rect -2 68 58 79
rect 10 61 27 63
rect 48 62 54 63
rect 10 59 23 61
rect 25 59 27 61
rect 10 58 27 59
rect 32 60 50 62
rect 52 60 54 62
rect 32 58 54 60
rect 10 32 14 58
rect 32 54 36 58
rect 18 50 36 54
rect 18 40 22 50
rect 20 38 22 40
rect 18 36 22 38
rect 50 38 54 47
rect 2 29 6 31
rect 2 27 4 29
rect 2 22 6 27
rect 10 28 23 32
rect 2 18 15 22
rect 19 21 23 28
rect 38 35 54 38
rect 38 33 40 35
rect 42 33 54 35
rect 38 32 54 33
rect 19 20 25 21
rect 19 18 21 20
rect 23 18 25 20
rect 19 17 25 18
rect -2 1 58 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 58 1
rect -2 -2 58 -1
<< ptie >>
rect 0 1 56 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 56 1
rect 0 -3 56 -1
<< ntie >>
rect 0 81 56 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 56 81
rect 0 77 56 79
<< nmos >>
rect 9 10 11 22
rect 16 10 18 22
rect 26 11 28 22
rect 35 16 37 27
rect 45 16 47 22
<< pmos >>
rect 10 45 12 70
rect 18 45 20 70
rect 28 45 30 70
rect 36 45 38 70
rect 45 46 47 55
<< polyct0 >>
rect 28 38 30 40
<< polyct1 >>
rect 50 60 52 62
rect 18 38 20 40
rect 40 33 42 35
rect 4 27 6 29
<< ndifct0 >>
rect 4 12 6 14
rect 40 18 42 20
rect 50 18 52 20
<< ndifct1 >>
rect 21 18 23 20
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
<< pdifct0 >>
rect 4 66 6 68
rect 4 59 6 61
rect 41 66 43 68
rect 50 51 52 53
<< pdifct1 >>
rect 23 59 25 61
<< alu0 >>
rect 3 66 4 68
rect 6 66 7 68
rect 3 61 7 66
rect 39 66 41 68
rect 43 66 45 68
rect 39 65 45 66
rect 3 59 4 61
rect 6 59 7 61
rect 3 57 7 59
rect 42 53 54 54
rect 42 51 50 53
rect 52 51 54 53
rect 42 50 54 51
rect 17 36 18 42
rect 42 46 46 50
rect 30 42 46 46
rect 30 41 34 42
rect 26 40 34 41
rect 26 38 28 40
rect 30 38 34 40
rect 26 37 34 38
rect 6 22 7 31
rect 30 28 34 37
rect 30 24 54 28
rect 38 20 44 21
rect 38 18 40 20
rect 42 18 44 20
rect 2 14 8 15
rect 2 12 4 14
rect 6 12 8 14
rect 38 12 44 18
rect 48 20 54 24
rect 48 18 50 20
rect 52 18 54 20
rect 48 17 54 18
<< labels >>
rlabel alu0 32 35 32 35 6 sn
rlabel alu0 51 22 51 22 6 sn
rlabel alu0 48 52 48 52 6 sn
rlabel alu1 4 28 4 28 6 a0
rlabel alu1 12 20 12 20 6 a0
rlabel alu1 20 44 20 44 6 s
rlabel alu1 12 48 12 48 6 z
rlabel alu1 20 60 20 60 6 z
rlabel alu1 28 6 28 6 6 vss
rlabel alu1 28 52 28 52 6 s
rlabel alu1 36 60 36 60 6 s
rlabel alu1 28 74 28 74 6 vdd
rlabel alu1 44 36 44 36 6 a1
rlabel alu1 52 40 52 40 6 a1
rlabel alu1 44 60 44 60 6 s
<< end >>
