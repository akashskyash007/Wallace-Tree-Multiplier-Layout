magic
tech scmos
timestamp 1199203152
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 13 66 15 70
rect 21 66 23 70
rect 31 66 33 70
rect 39 66 41 70
rect 13 36 15 39
rect 21 36 23 39
rect 9 34 15 36
rect 9 32 11 34
rect 13 32 15 34
rect 9 30 15 32
rect 19 34 25 36
rect 31 35 33 39
rect 39 36 41 39
rect 19 32 21 34
rect 23 32 25 34
rect 19 30 25 32
rect 29 33 35 35
rect 29 31 31 33
rect 33 31 35 33
rect 9 26 11 30
rect 19 26 21 30
rect 29 29 35 31
rect 39 34 48 36
rect 39 32 44 34
rect 46 32 48 34
rect 39 30 48 32
rect 29 23 31 29
rect 41 23 43 30
rect 9 7 11 12
rect 19 7 21 12
rect 29 7 31 12
rect 41 7 43 12
<< ndif >>
rect 4 18 9 26
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 12 19 22
rect 21 23 26 26
rect 21 16 29 23
rect 21 14 24 16
rect 26 14 29 16
rect 21 12 29 14
rect 31 12 41 23
rect 43 18 48 23
rect 43 16 50 18
rect 43 14 46 16
rect 48 14 50 16
rect 43 12 50 14
rect 33 7 39 12
rect 33 5 35 7
rect 37 5 39 7
rect 33 3 39 5
<< pdif >>
rect 5 64 13 66
rect 5 62 8 64
rect 10 62 13 64
rect 5 39 13 62
rect 15 39 21 66
rect 23 57 31 66
rect 23 55 26 57
rect 28 55 31 57
rect 23 39 31 55
rect 33 39 39 66
rect 41 64 48 66
rect 41 62 44 64
rect 46 62 48 64
rect 41 57 48 62
rect 41 55 44 57
rect 46 55 48 57
rect 41 39 48 55
<< alu1 >>
rect -2 64 58 72
rect 2 57 30 58
rect 2 55 26 57
rect 28 55 30 57
rect 2 54 30 55
rect 2 25 6 54
rect 34 50 38 59
rect 10 46 23 50
rect 34 46 47 50
rect 10 34 14 46
rect 10 32 11 34
rect 13 32 14 34
rect 10 29 14 32
rect 18 38 39 42
rect 18 34 24 38
rect 43 34 47 46
rect 18 32 21 34
rect 23 32 24 34
rect 18 29 24 32
rect 29 33 39 34
rect 29 31 31 33
rect 33 31 39 33
rect 29 30 39 31
rect 43 32 44 34
rect 46 32 47 34
rect 43 30 47 32
rect 33 26 39 30
rect 2 24 18 25
rect 2 22 14 24
rect 16 22 18 24
rect 33 22 47 26
rect 2 21 18 22
rect -2 7 58 8
rect -2 5 35 7
rect 37 5 58 7
rect -2 0 58 5
<< nmos >>
rect 9 12 11 26
rect 19 12 21 26
rect 29 12 31 23
rect 41 12 43 23
<< pmos >>
rect 13 39 15 66
rect 21 39 23 66
rect 31 39 33 66
rect 39 39 41 66
<< polyct1 >>
rect 11 32 13 34
rect 21 32 23 34
rect 31 31 33 33
rect 44 32 46 34
<< ndifct0 >>
rect 4 14 6 16
rect 24 14 26 16
rect 46 14 48 16
<< ndifct1 >>
rect 14 22 16 24
rect 35 5 37 7
<< pdifct0 >>
rect 8 62 10 64
rect 44 62 46 64
rect 44 55 46 57
<< pdifct1 >>
rect 26 55 28 57
<< alu0 >>
rect 6 62 8 64
rect 10 62 12 64
rect 6 61 12 62
rect 42 62 44 64
rect 46 62 48 64
rect 42 57 48 62
rect 42 55 44 57
rect 46 55 48 57
rect 42 54 48 55
rect 2 16 50 17
rect 2 14 4 16
rect 6 14 24 16
rect 26 14 46 16
rect 48 14 50 16
rect 2 13 50 14
<< labels >>
rlabel alu0 26 15 26 15 6 n3
rlabel alu1 4 36 4 36 6 z
rlabel alu1 20 32 20 32 6 b2
rlabel alu1 12 36 12 36 6 b1
rlabel alu1 20 48 20 48 6 b1
rlabel alu1 20 56 20 56 6 z
rlabel alu1 12 56 12 56 6 z
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 36 28 36 28 6 a2
rlabel alu1 36 40 36 40 6 b2
rlabel alu1 28 40 28 40 6 b2
rlabel alu1 36 56 36 56 6 a1
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 24 44 24 6 a2
rlabel alu1 44 48 44 48 6 a1
<< end >>
