magic
tech scmos
timestamp 1199203520
<< ab >>
rect 0 0 184 72
<< nwell >>
rect -5 32 189 77
<< pwell >>
rect -5 -5 189 32
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 29 68 53 70
rect 29 65 31 68
rect 39 65 41 68
rect 51 51 53 68
rect 63 66 65 70
rect 73 66 75 70
rect 83 66 85 70
rect 93 66 95 70
rect 116 66 118 70
rect 123 66 125 70
rect 133 66 135 70
rect 151 66 153 70
rect 161 66 163 70
rect 48 49 54 51
rect 48 47 50 49
rect 52 47 54 49
rect 48 45 54 47
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 63 37 65 40
rect 73 37 75 40
rect 9 33 22 35
rect 29 33 41 35
rect 61 35 75 37
rect 83 35 85 38
rect 93 35 95 38
rect 116 35 118 38
rect 61 33 67 35
rect 16 31 18 33
rect 20 31 22 33
rect 16 29 22 31
rect 9 24 11 29
rect 16 27 28 29
rect 16 24 18 27
rect 26 24 28 27
rect 33 24 35 33
rect 61 31 63 33
rect 65 31 67 33
rect 80 33 108 35
rect 80 31 82 33
rect 45 26 47 31
rect 55 29 67 31
rect 55 26 57 29
rect 65 26 67 29
rect 75 29 82 31
rect 102 31 104 33
rect 106 31 108 33
rect 102 29 108 31
rect 112 33 118 35
rect 112 31 114 33
rect 116 31 118 33
rect 123 35 125 38
rect 133 35 135 38
rect 151 35 153 38
rect 161 35 163 38
rect 123 32 126 35
rect 133 33 153 35
rect 157 33 163 35
rect 112 29 118 31
rect 75 26 77 29
rect 86 26 92 28
rect 114 26 116 29
rect 124 26 126 32
rect 137 31 139 33
rect 141 31 148 33
rect 137 29 148 31
rect 157 31 159 33
rect 161 31 163 33
rect 157 29 163 31
rect 146 26 148 29
rect 86 24 88 26
rect 90 24 92 26
rect 86 23 92 24
rect 85 21 97 23
rect 85 18 87 21
rect 95 18 97 21
rect 9 4 11 12
rect 16 8 18 12
rect 26 8 28 12
rect 33 4 35 12
rect 9 2 35 4
rect 45 4 47 12
rect 55 8 57 12
rect 65 8 67 12
rect 75 4 77 12
rect 133 16 139 18
rect 133 14 135 16
rect 137 14 139 16
rect 158 23 160 29
rect 133 12 139 14
rect 114 7 116 12
rect 124 9 126 12
rect 133 9 135 12
rect 146 10 148 15
rect 124 7 135 9
rect 45 2 77 4
rect 85 2 87 6
rect 95 2 97 6
rect 158 7 160 12
<< ndif >>
rect 37 24 45 26
rect 4 18 9 24
rect 2 16 9 18
rect 2 14 4 16
rect 6 14 9 16
rect 2 12 9 14
rect 11 12 16 24
rect 18 22 26 24
rect 18 20 21 22
rect 23 20 26 22
rect 18 12 26 20
rect 28 12 33 24
rect 35 12 45 24
rect 47 24 55 26
rect 47 22 50 24
rect 52 22 55 24
rect 47 12 55 22
rect 57 16 65 26
rect 57 14 60 16
rect 62 14 65 16
rect 57 12 65 14
rect 67 24 75 26
rect 67 22 70 24
rect 72 22 75 24
rect 67 17 75 22
rect 67 15 70 17
rect 72 15 75 17
rect 67 12 75 15
rect 77 18 82 26
rect 109 19 114 26
rect 77 16 85 18
rect 77 14 80 16
rect 82 14 85 16
rect 77 12 85 14
rect 37 7 43 12
rect 37 5 39 7
rect 41 5 43 7
rect 37 3 43 5
rect 80 6 85 12
rect 87 16 95 18
rect 87 14 90 16
rect 92 14 95 16
rect 87 6 95 14
rect 97 9 103 18
rect 107 17 114 19
rect 107 15 109 17
rect 111 15 114 17
rect 107 13 114 15
rect 109 12 114 13
rect 116 24 124 26
rect 116 22 119 24
rect 121 22 124 24
rect 116 12 124 22
rect 126 24 133 26
rect 126 22 129 24
rect 131 22 133 24
rect 126 20 133 22
rect 139 24 146 26
rect 139 22 141 24
rect 143 22 146 24
rect 139 20 146 22
rect 126 12 131 20
rect 141 15 146 20
rect 148 23 156 26
rect 148 15 158 23
rect 97 7 105 9
rect 150 12 158 15
rect 160 18 165 23
rect 160 16 167 18
rect 160 14 163 16
rect 165 14 167 16
rect 160 12 167 14
rect 97 6 101 7
rect 99 5 101 6
rect 103 5 105 7
rect 99 3 105 5
rect 150 7 156 12
rect 150 5 152 7
rect 154 5 156 7
rect 150 3 156 5
<< pdif >>
rect 4 59 9 65
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 50 9 55
rect 2 48 4 50
rect 6 48 9 50
rect 2 46 9 48
rect 4 38 9 46
rect 11 49 19 65
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 57 29 65
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 42 39 65
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 59 46 65
rect 41 57 48 59
rect 41 55 44 57
rect 46 55 48 57
rect 41 53 48 55
rect 41 38 46 53
rect 56 64 63 66
rect 56 62 58 64
rect 60 62 63 64
rect 56 57 63 62
rect 56 55 58 57
rect 60 55 63 57
rect 56 40 63 55
rect 65 57 73 66
rect 65 55 68 57
rect 70 55 73 57
rect 65 50 73 55
rect 65 48 68 50
rect 70 48 73 50
rect 65 40 73 48
rect 75 64 83 66
rect 75 62 78 64
rect 80 62 83 64
rect 75 40 83 62
rect 78 38 83 40
rect 85 44 93 66
rect 85 42 88 44
rect 90 42 93 44
rect 85 38 93 42
rect 95 64 116 66
rect 95 62 98 64
rect 100 62 106 64
rect 108 62 116 64
rect 95 57 116 62
rect 95 55 106 57
rect 108 55 116 57
rect 95 38 116 55
rect 118 38 123 66
rect 125 58 133 66
rect 125 56 128 58
rect 130 56 133 58
rect 125 38 133 56
rect 135 60 140 66
rect 135 58 142 60
rect 135 56 138 58
rect 140 56 142 58
rect 135 54 142 56
rect 135 38 140 54
rect 146 50 151 66
rect 144 48 151 50
rect 144 46 146 48
rect 148 46 151 48
rect 144 44 151 46
rect 146 38 151 44
rect 153 64 161 66
rect 153 62 156 64
rect 158 62 161 64
rect 153 38 161 62
rect 163 51 168 66
rect 163 49 170 51
rect 163 47 166 49
rect 168 47 170 49
rect 163 42 170 47
rect 163 40 166 42
rect 168 40 170 42
rect 163 38 170 40
<< alu1 >>
rect -2 67 186 72
rect -2 65 174 67
rect 176 65 186 67
rect -2 64 186 65
rect 2 57 48 58
rect 2 55 4 57
rect 6 55 24 57
rect 26 55 44 57
rect 46 55 48 57
rect 2 54 48 55
rect 2 50 6 54
rect 2 48 4 50
rect 2 26 6 48
rect 57 33 87 34
rect 57 31 63 33
rect 65 31 87 33
rect 57 30 87 31
rect 2 22 24 26
rect 20 20 21 22
rect 23 20 24 22
rect 81 28 87 30
rect 81 26 91 28
rect 81 24 88 26
rect 90 24 91 26
rect 81 22 91 24
rect 20 18 24 20
rect 20 16 64 18
rect 20 14 60 16
rect 62 14 64 16
rect 58 13 64 14
rect 129 38 142 42
rect 138 33 142 38
rect 154 35 158 51
rect 138 31 139 33
rect 141 31 142 33
rect 138 29 142 31
rect 146 33 162 35
rect 146 31 159 33
rect 161 31 162 33
rect 146 29 162 31
rect 154 21 158 29
rect -2 7 186 8
rect -2 5 39 7
rect 41 5 101 7
rect 103 5 139 7
rect 141 5 152 7
rect 154 5 173 7
rect 175 5 186 7
rect -2 0 186 5
<< ptie >>
rect 137 7 143 9
rect 137 5 139 7
rect 141 5 143 7
rect 137 3 143 5
rect 171 7 177 26
rect 171 5 173 7
rect 175 5 177 7
rect 171 3 177 5
<< ntie >>
rect 172 67 178 69
rect 172 65 174 67
rect 176 65 178 67
rect 172 55 178 65
<< nmos >>
rect 9 12 11 24
rect 16 12 18 24
rect 26 12 28 24
rect 33 12 35 24
rect 45 12 47 26
rect 55 12 57 26
rect 65 12 67 26
rect 75 12 77 26
rect 85 6 87 18
rect 95 6 97 18
rect 114 12 116 26
rect 124 12 126 26
rect 146 15 148 26
rect 158 12 160 23
<< pmos >>
rect 9 38 11 65
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 65
rect 63 40 65 66
rect 73 40 75 66
rect 83 38 85 66
rect 93 38 95 66
rect 116 38 118 66
rect 123 38 125 66
rect 133 38 135 66
rect 151 38 153 66
rect 161 38 163 66
<< polyct0 >>
rect 50 47 52 49
rect 18 31 20 33
rect 104 31 106 33
rect 114 31 116 33
rect 135 14 137 16
<< polyct1 >>
rect 63 31 65 33
rect 139 31 141 33
rect 159 31 161 33
rect 88 24 90 26
<< ndifct0 >>
rect 4 14 6 16
rect 50 22 52 24
rect 70 22 72 24
rect 70 15 72 17
rect 80 14 82 16
rect 90 14 92 16
rect 109 15 111 17
rect 119 22 121 24
rect 129 22 131 24
rect 141 22 143 24
rect 163 14 165 16
<< ndifct1 >>
rect 21 20 23 22
rect 60 14 62 16
rect 39 5 41 7
rect 101 5 103 7
rect 152 5 154 7
<< ntiect1 >>
rect 174 65 176 67
<< ptiect1 >>
rect 139 5 141 7
rect 173 5 175 7
<< pdifct0 >>
rect 14 47 16 49
rect 14 40 16 42
rect 34 40 36 42
rect 58 62 60 64
rect 58 55 60 57
rect 68 55 70 57
rect 68 48 70 50
rect 78 62 80 64
rect 88 42 90 44
rect 98 62 100 64
rect 106 62 108 64
rect 106 55 108 57
rect 128 56 130 58
rect 138 56 140 58
rect 146 46 148 48
rect 156 62 158 64
rect 166 47 168 49
rect 166 40 168 42
<< pdifct1 >>
rect 4 55 6 57
rect 4 48 6 50
rect 24 55 26 57
rect 44 55 46 57
<< alu0 >>
rect 56 62 58 64
rect 60 62 62 64
rect 56 57 62 62
rect 77 62 78 64
rect 80 62 81 64
rect 77 60 81 62
rect 97 62 98 64
rect 100 62 101 64
rect 97 60 101 62
rect 105 62 106 64
rect 108 62 109 64
rect 56 55 58 57
rect 60 55 62 57
rect 56 54 62 55
rect 67 57 71 59
rect 67 55 68 57
rect 70 55 71 57
rect 67 54 71 55
rect 105 57 109 62
rect 154 62 156 64
rect 158 62 160 64
rect 154 61 160 62
rect 105 55 106 57
rect 108 55 109 57
rect 6 46 7 54
rect 67 50 99 54
rect 105 53 109 55
rect 113 58 132 59
rect 113 56 128 58
rect 130 56 132 58
rect 113 55 132 56
rect 136 58 142 59
rect 136 56 138 58
rect 140 56 169 58
rect 12 49 68 50
rect 12 47 14 49
rect 16 47 50 49
rect 52 48 68 49
rect 70 48 71 50
rect 52 47 71 48
rect 12 46 71 47
rect 12 42 17 46
rect 87 44 91 46
rect 12 40 14 42
rect 16 40 17 42
rect 12 38 17 40
rect 32 42 38 43
rect 87 42 88 44
rect 90 42 91 44
rect 32 40 34 42
rect 36 40 38 42
rect 32 34 38 40
rect 48 38 91 42
rect 48 34 52 38
rect 16 33 52 34
rect 16 31 18 33
rect 20 31 52 33
rect 16 30 52 31
rect 48 25 52 30
rect 48 24 74 25
rect 48 22 50 24
rect 52 22 70 24
rect 72 22 74 24
rect 48 21 74 22
rect 3 16 7 18
rect 3 14 4 16
rect 6 14 7 16
rect 3 8 7 14
rect 69 17 74 21
rect 95 17 99 50
rect 113 49 117 55
rect 136 54 169 56
rect 103 45 117 49
rect 121 48 150 49
rect 121 46 146 48
rect 148 46 150 48
rect 121 45 150 46
rect 103 33 107 45
rect 121 34 125 45
rect 103 31 104 33
rect 106 31 107 33
rect 103 25 107 31
rect 112 33 131 34
rect 112 31 114 33
rect 116 31 131 33
rect 112 30 131 31
rect 127 25 131 30
rect 165 49 169 54
rect 165 47 166 49
rect 168 47 169 49
rect 165 42 169 47
rect 165 40 166 42
rect 168 40 169 42
rect 103 24 123 25
rect 103 22 119 24
rect 121 22 123 24
rect 103 21 123 22
rect 127 24 145 25
rect 127 22 129 24
rect 131 22 141 24
rect 143 22 145 24
rect 127 21 145 22
rect 69 15 70 17
rect 72 15 74 17
rect 69 13 74 15
rect 78 16 84 17
rect 78 14 80 16
rect 82 14 84 16
rect 78 8 84 14
rect 88 16 99 17
rect 88 14 90 16
rect 92 14 99 16
rect 88 13 99 14
rect 107 17 113 18
rect 165 17 169 40
rect 107 15 109 17
rect 111 16 169 17
rect 111 15 135 16
rect 107 14 135 15
rect 137 14 163 16
rect 165 14 169 16
rect 107 13 169 14
<< labels >>
rlabel alu0 35 36 35 36 6 zn
rlabel alu0 14 44 14 44 6 cn
rlabel alu0 71 19 71 19 6 zn
rlabel alu0 61 23 61 23 6 zn
rlabel alu0 41 48 41 48 6 cn
rlabel alu0 93 15 93 15 6 cn
rlabel alu0 113 23 113 23 6 iz
rlabel alu0 123 39 123 39 6 bn
rlabel alu0 105 35 105 35 6 iz
rlabel alu0 89 42 89 42 6 zn
rlabel alu0 122 57 122 57 6 iz
rlabel alu0 83 52 83 52 6 cn
rlabel alu0 138 15 138 15 6 an
rlabel alu0 136 23 136 23 6 bn
rlabel alu0 135 47 135 47 6 bn
rlabel alu0 139 56 139 56 6 an
rlabel alu0 167 35 167 35 6 an
rlabel alu1 28 16 28 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 20 24 20 24 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 20 56 20 56 6 z
rlabel alu1 12 56 12 56 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 60 16 60 16 6 z
rlabel alu1 52 16 52 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 76 32 76 32 6 c
rlabel alu1 84 28 84 28 6 c
rlabel alu1 60 32 60 32 6 c
rlabel alu1 68 32 68 32 6 c
rlabel alu1 44 56 44 56 6 z
rlabel alu1 92 4 92 4 6 vss
rlabel alu1 132 40 132 40 6 b
rlabel alu1 92 68 92 68 6 vdd
rlabel polyct1 140 32 140 32 6 b
rlabel alu1 148 32 148 32 6 a
rlabel alu1 156 24 156 24 6 a
rlabel alu1 156 36 156 36 6 a
<< end >>
