magic
tech scmos
timestamp 1199203398
<< ab >>
rect 0 0 24 80
<< nwell >>
rect -5 36 29 88
<< pwell >>
rect -5 -8 29 36
<< poly >>
rect 12 61 14 65
rect 12 40 14 43
rect 4 38 14 40
rect 4 36 6 38
rect 8 36 14 38
rect 4 34 14 36
rect 12 30 14 34
rect 12 6 14 10
<< ndif >>
rect 3 28 12 30
rect 3 26 5 28
rect 7 26 12 28
rect 3 21 12 26
rect 3 19 5 21
rect 7 19 12 21
rect 3 10 12 19
rect 14 21 22 30
rect 14 19 18 21
rect 20 19 22 21
rect 14 14 22 19
rect 14 12 18 14
rect 20 12 22 14
rect 14 10 22 12
<< pdif >>
rect 3 71 10 73
rect 3 69 6 71
rect 8 69 10 71
rect 3 63 10 69
rect 3 61 6 63
rect 8 61 10 63
rect 3 55 12 61
rect 3 53 6 55
rect 8 53 12 55
rect 3 47 12 53
rect 3 45 6 47
rect 8 45 12 47
rect 3 43 12 45
rect 14 55 22 61
rect 14 53 18 55
rect 20 53 22 55
rect 14 47 22 53
rect 14 45 18 47
rect 20 45 22 47
rect 14 43 22 45
<< alu1 >>
rect -2 81 26 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 26 81
rect -2 71 26 79
rect -2 69 6 71
rect 8 69 26 71
rect -2 68 26 69
rect 17 55 22 63
rect 17 53 18 55
rect 20 53 22 55
rect 17 47 22 53
rect 17 45 18 47
rect 20 45 22 47
rect 17 31 22 45
rect 2 28 22 31
rect 2 26 5 28
rect 7 26 22 28
rect 2 25 22 26
rect 2 21 8 25
rect 2 19 5 21
rect 7 19 8 21
rect 2 17 8 19
rect -2 1 26 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 26 1
rect -2 -2 26 -1
<< ptie >>
rect 0 1 24 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 24 1
rect 0 -3 24 -1
<< ntie >>
rect 0 81 24 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 24 81
rect 0 77 24 79
<< nmos >>
rect 12 10 14 30
<< pmos >>
rect 12 43 14 61
<< polyct0 >>
rect 6 36 8 38
<< ndifct0 >>
rect 18 19 20 21
rect 18 12 20 14
<< ndifct1 >>
rect 5 26 7 28
rect 5 19 7 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
<< pdifct0 >>
rect 6 61 8 63
rect 6 53 8 55
rect 6 45 8 47
<< pdifct1 >>
rect 6 69 8 71
rect 18 53 20 55
rect 18 45 20 47
<< alu0 >>
rect 4 63 10 68
rect 4 61 6 63
rect 8 61 10 63
rect 4 55 10 61
rect 4 53 6 55
rect 8 53 10 55
rect 4 47 10 53
rect 4 45 6 47
rect 8 45 10 47
rect 4 38 10 45
rect 4 36 6 38
rect 8 36 10 38
rect 4 35 10 36
rect 16 21 22 22
rect 16 19 18 21
rect 20 19 22 21
rect 16 14 22 19
rect 16 12 18 14
rect 20 12 22 14
<< labels >>
rlabel alu1 4 24 4 24 6 z
rlabel alu1 12 6 12 6 6 vss
rlabel alu1 12 28 12 28 6 z
rlabel alu1 12 74 12 74 6 vdd
rlabel alu1 20 44 20 44 6 z
<< end >>
