magic
tech scmos
timestamp 1199203426
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 47 66 49 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 36 31 39
rect 58 52 60 57
rect 68 52 70 57
rect 29 35 39 36
rect 47 35 49 38
rect 58 35 60 38
rect 68 35 70 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 29 34 42 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 36 33 42 34
rect 36 31 38 33
rect 40 31 42 33
rect 13 26 15 29
rect 20 26 22 29
rect 30 26 32 30
rect 36 29 42 31
rect 40 26 42 29
rect 47 33 54 35
rect 58 33 78 35
rect 47 31 50 33
rect 52 31 54 33
rect 47 29 54 31
rect 47 26 49 29
rect 63 26 65 33
rect 72 31 74 33
rect 76 31 78 33
rect 72 29 78 31
rect 13 8 15 13
rect 20 8 22 13
rect 40 8 42 12
rect 47 8 49 12
rect 30 4 32 7
rect 63 4 65 13
rect 30 2 65 4
<< ndif >>
rect 4 13 13 26
rect 15 13 20 26
rect 22 17 30 26
rect 22 15 25 17
rect 27 15 30 17
rect 22 13 30 15
rect 4 7 11 13
rect 25 7 30 13
rect 32 22 40 26
rect 32 20 35 22
rect 37 20 40 22
rect 32 12 40 20
rect 42 12 47 26
rect 49 17 63 26
rect 49 15 58 17
rect 60 15 63 17
rect 49 13 63 15
rect 65 24 72 26
rect 65 22 68 24
rect 70 22 72 24
rect 65 20 72 22
rect 65 13 70 20
rect 49 12 61 13
rect 32 7 37 12
rect 4 5 7 7
rect 9 5 11 7
rect 4 3 11 5
<< pdif >>
rect 4 59 9 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 53 9 55
rect 4 38 9 53
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 38 19 47
rect 21 49 29 66
rect 21 47 24 49
rect 26 47 29 49
rect 21 39 29 47
rect 31 64 38 66
rect 31 62 34 64
rect 36 62 38 64
rect 31 55 38 62
rect 31 39 36 55
rect 42 51 47 66
rect 40 49 47 51
rect 40 47 42 49
rect 44 47 47 49
rect 40 45 47 47
rect 21 38 26 39
rect 42 38 47 45
rect 49 64 56 66
rect 49 62 52 64
rect 54 62 56 64
rect 72 67 78 69
rect 72 65 74 67
rect 76 65 78 67
rect 49 52 56 62
rect 72 52 78 65
rect 49 38 58 52
rect 60 49 68 52
rect 60 47 63 49
rect 65 47 68 49
rect 60 42 68 47
rect 60 40 63 42
rect 65 40 68 42
rect 60 38 68 40
rect 70 38 78 52
<< alu1 >>
rect -2 67 82 72
rect -2 65 63 67
rect 65 65 74 67
rect 76 65 82 67
rect -2 64 82 65
rect 64 54 78 59
rect 2 49 17 51
rect 2 47 14 49
rect 16 47 17 49
rect 2 45 17 47
rect 2 18 6 45
rect 34 33 46 35
rect 34 31 38 33
rect 40 31 46 33
rect 34 29 46 31
rect 50 33 54 35
rect 52 31 54 33
rect 2 17 31 18
rect 2 15 25 17
rect 27 15 31 17
rect 2 14 31 15
rect 42 13 46 29
rect 50 26 54 31
rect 74 35 78 54
rect 73 33 78 35
rect 73 31 74 33
rect 76 31 78 33
rect 73 29 78 31
rect 50 22 63 26
rect 50 13 54 22
rect -2 7 82 8
rect -2 5 7 7
rect 9 5 73 7
rect 75 5 82 7
rect -2 0 82 5
<< ptie >>
rect 71 7 77 9
rect 71 5 73 7
rect 75 5 77 7
rect 71 3 77 5
<< ntie >>
rect 60 67 68 69
rect 60 65 63 67
rect 65 65 68 67
rect 60 63 68 65
<< nmos >>
rect 13 13 15 26
rect 20 13 22 26
rect 30 7 32 26
rect 40 12 42 26
rect 47 12 49 26
rect 63 13 65 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 39 31 66
rect 47 38 49 66
rect 58 38 60 52
rect 68 38 70 52
<< polyct0 >>
rect 11 31 13 33
rect 21 31 23 33
<< polyct1 >>
rect 38 31 40 33
rect 50 31 52 33
rect 74 31 76 33
<< ndifct0 >>
rect 35 20 37 22
rect 58 15 60 17
rect 68 22 70 24
<< ndifct1 >>
rect 25 15 27 17
rect 7 5 9 7
<< ntiect1 >>
rect 63 65 65 67
<< ptiect1 >>
rect 73 5 75 7
<< pdifct0 >>
rect 4 55 6 57
rect 24 47 26 49
rect 34 62 36 64
rect 42 47 44 49
rect 52 62 54 64
rect 63 47 65 49
rect 63 40 65 42
<< pdifct1 >>
rect 14 47 16 49
rect 74 65 76 67
<< alu0 >>
rect 32 62 34 64
rect 36 62 38 64
rect 32 61 38 62
rect 50 62 52 64
rect 54 62 56 64
rect 50 61 56 62
rect 2 57 54 58
rect 2 55 4 57
rect 6 55 54 57
rect 2 54 54 55
rect 20 49 46 50
rect 20 47 24 49
rect 26 47 42 49
rect 44 47 46 49
rect 20 46 46 47
rect 20 42 24 46
rect 50 43 54 54
rect 61 49 67 50
rect 61 47 63 49
rect 65 47 67 49
rect 61 43 67 47
rect 10 38 24 42
rect 27 42 70 43
rect 27 40 63 42
rect 65 40 70 42
rect 27 39 70 40
rect 10 33 14 38
rect 27 34 31 39
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 19 33 31 34
rect 19 31 21 33
rect 23 31 31 33
rect 19 30 31 31
rect 49 29 50 35
rect 10 22 38 26
rect 34 20 35 22
rect 37 20 38 22
rect 34 18 38 20
rect 66 26 70 39
rect 66 24 71 26
rect 66 22 68 24
rect 70 22 71 24
rect 66 20 71 22
rect 57 17 61 19
rect 57 15 58 17
rect 60 15 61 17
rect 57 8 61 15
<< labels >>
rlabel polyct0 12 32 12 32 6 an
rlabel alu0 25 32 25 32 6 bn
rlabel alu0 24 24 24 24 6 an
rlabel alu0 33 48 33 48 6 an
rlabel alu0 28 56 28 56 6 bn
rlabel alu0 68 31 68 31 6 bn
rlabel alu0 48 41 48 41 6 bn
rlabel alu0 64 44 64 44 6 bn
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 36 32 36 32 6 a2
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 44 24 44 24 6 a2
rlabel alu1 52 24 52 24 6 a1
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 60 24 60 24 6 a1
rlabel alu1 76 44 76 44 6 b
rlabel alu1 68 56 68 56 6 b
<< end >>
