magic
tech scmos
timestamp 1199202616
<< ab >>
rect 0 0 72 72
<< nwell >>
rect -5 32 77 77
<< pwell >>
rect -5 -5 77 32
<< poly >>
rect 9 62 11 67
rect 19 65 21 70
rect 29 65 31 70
rect 39 62 41 67
rect 49 62 51 67
rect 59 56 61 61
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 49 35 51 38
rect 59 35 61 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 33 35
rect 19 31 27 33
rect 29 31 33 33
rect 19 29 33 31
rect 12 26 14 29
rect 19 26 21 29
rect 31 26 33 29
rect 38 33 51 35
rect 38 31 43 33
rect 45 31 51 33
rect 38 29 51 31
rect 55 33 63 35
rect 55 31 59 33
rect 61 31 63 33
rect 55 29 63 31
rect 38 26 40 29
rect 48 26 50 29
rect 55 26 57 29
rect 12 2 14 6
rect 19 2 21 6
rect 31 2 33 6
rect 38 2 40 6
rect 48 2 50 6
rect 55 2 57 6
<< ndif >>
rect 5 24 12 26
rect 5 22 7 24
rect 9 22 12 24
rect 5 17 12 22
rect 5 15 7 17
rect 9 15 12 17
rect 5 13 12 15
rect 7 6 12 13
rect 14 6 19 26
rect 21 10 31 26
rect 21 8 25 10
rect 27 8 31 10
rect 21 6 31 8
rect 33 6 38 26
rect 40 17 48 26
rect 40 15 43 17
rect 45 15 48 17
rect 40 6 48 15
rect 50 6 55 26
rect 57 10 65 26
rect 57 8 60 10
rect 62 8 65 10
rect 57 6 65 8
<< pdif >>
rect 14 62 19 65
rect 2 60 9 62
rect 2 58 4 60
rect 6 58 9 60
rect 2 52 9 58
rect 2 50 4 52
rect 6 50 9 52
rect 2 38 9 50
rect 11 49 19 62
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 63 29 65
rect 21 61 24 63
rect 26 61 29 63
rect 21 56 29 61
rect 21 54 24 56
rect 26 54 29 56
rect 21 38 29 54
rect 31 62 36 65
rect 31 57 39 62
rect 31 55 34 57
rect 36 55 39 57
rect 31 49 39 55
rect 31 47 34 49
rect 36 47 39 49
rect 31 38 39 47
rect 41 60 49 62
rect 41 58 44 60
rect 46 58 49 60
rect 41 38 49 58
rect 51 56 56 62
rect 51 49 59 56
rect 51 47 54 49
rect 56 47 59 49
rect 51 38 59 47
rect 61 54 68 56
rect 61 52 64 54
rect 66 52 68 54
rect 61 38 68 52
<< alu1 >>
rect -2 67 74 72
rect -2 65 63 67
rect 65 65 74 67
rect -2 64 74 65
rect 33 57 38 59
rect 33 55 34 57
rect 36 55 38 57
rect 33 50 38 55
rect 12 49 58 50
rect 12 47 14 49
rect 16 47 34 49
rect 36 47 54 49
rect 56 47 58 49
rect 12 46 58 47
rect 12 43 18 46
rect 2 42 18 43
rect 2 40 14 42
rect 16 40 18 42
rect 2 39 18 40
rect 2 25 6 39
rect 25 38 63 42
rect 10 33 21 35
rect 10 31 11 33
rect 13 31 21 33
rect 10 29 21 31
rect 25 33 31 38
rect 25 31 27 33
rect 29 31 31 33
rect 25 30 31 31
rect 41 33 47 34
rect 41 31 43 33
rect 45 31 47 33
rect 17 26 21 29
rect 41 26 47 31
rect 57 33 63 38
rect 57 31 59 33
rect 61 31 63 33
rect 57 30 63 31
rect 2 24 11 25
rect 2 22 7 24
rect 9 22 11 24
rect 17 22 47 26
rect 2 21 11 22
rect 5 18 11 21
rect 5 17 47 18
rect 5 15 7 17
rect 9 15 43 17
rect 45 15 47 17
rect 5 14 47 15
rect -2 0 74 8
<< ntie >>
rect 61 67 67 69
rect 61 65 63 67
rect 65 65 67 67
rect 61 63 67 65
<< nmos >>
rect 12 6 14 26
rect 19 6 21 26
rect 31 6 33 26
rect 38 6 40 26
rect 48 6 50 26
rect 55 6 57 26
<< pmos >>
rect 9 38 11 62
rect 19 38 21 65
rect 29 38 31 65
rect 39 38 41 62
rect 49 38 51 62
rect 59 38 61 56
<< polyct1 >>
rect 11 31 13 33
rect 27 31 29 33
rect 43 31 45 33
rect 59 31 61 33
<< ndifct0 >>
rect 25 8 27 10
rect 60 8 62 10
<< ndifct1 >>
rect 7 22 9 24
rect 7 15 9 17
rect 43 15 45 17
<< ntiect1 >>
rect 63 65 65 67
<< pdifct0 >>
rect 4 58 6 60
rect 4 50 6 52
rect 24 61 26 63
rect 24 54 26 56
rect 44 58 46 60
rect 64 52 66 54
<< pdifct1 >>
rect 14 47 16 49
rect 14 40 16 42
rect 34 55 36 57
rect 34 47 36 49
rect 54 47 56 49
<< alu0 >>
rect 3 60 7 64
rect 3 58 4 60
rect 6 58 7 60
rect 3 52 7 58
rect 22 63 28 64
rect 22 61 24 63
rect 26 61 28 63
rect 22 56 28 61
rect 43 60 47 64
rect 22 54 24 56
rect 26 54 28 56
rect 22 53 28 54
rect 43 58 44 60
rect 46 58 47 60
rect 43 56 47 58
rect 3 50 4 52
rect 6 50 7 52
rect 63 54 67 64
rect 63 52 64 54
rect 66 52 67 54
rect 63 50 67 52
rect 3 48 7 50
rect 23 10 29 11
rect 23 8 25 10
rect 27 8 29 10
rect 58 10 64 11
rect 58 8 60 10
rect 62 8 64 10
<< labels >>
rlabel alu1 12 16 12 16 6 z
rlabel polyct1 12 32 12 32 6 b
rlabel alu1 4 32 4 32 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 24 20 24 6 b
rlabel alu1 28 24 28 24 6 b
rlabel alu1 28 36 28 36 6 a
rlabel alu1 20 48 20 48 6 z
rlabel alu1 28 48 28 48 6 z
rlabel alu1 36 4 36 4 6 vss
rlabel ndifct1 44 16 44 16 6 z
rlabel alu1 36 16 36 16 6 z
rlabel alu1 36 24 36 24 6 b
rlabel alu1 44 28 44 28 6 b
rlabel alu1 44 40 44 40 6 a
rlabel alu1 52 40 52 40 6 a
rlabel alu1 36 40 36 40 6 a
rlabel alu1 36 52 36 52 6 z
rlabel alu1 52 48 52 48 6 z
rlabel alu1 44 48 44 48 6 z
rlabel alu1 36 68 36 68 6 vdd
rlabel alu1 60 36 60 36 6 a
<< end >>
