magic
tech scmos
timestamp 1199202361
<< ab >>
rect 0 0 64 72
<< nwell >>
rect -5 32 69 77
<< pwell >>
rect -5 -5 69 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 54 51 59
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 39 35 41 38
rect 9 33 41 35
rect 22 31 37 33
rect 39 31 41 33
rect 22 29 41 31
rect 49 35 51 38
rect 49 33 55 35
rect 49 31 51 33
rect 53 31 55 33
rect 49 29 55 31
rect 22 26 24 29
rect 32 26 34 29
rect 22 5 24 10
rect 32 5 34 10
<< ndif >>
rect 14 22 22 26
rect 14 20 17 22
rect 19 20 22 22
rect 14 14 22 20
rect 14 12 17 14
rect 19 12 22 14
rect 14 10 22 12
rect 24 24 32 26
rect 24 22 27 24
rect 29 22 32 24
rect 24 17 32 22
rect 24 15 27 17
rect 29 15 32 17
rect 24 10 32 15
rect 34 22 42 26
rect 34 20 37 22
rect 39 20 42 22
rect 34 14 42 20
rect 34 12 37 14
rect 39 12 42 14
rect 34 10 42 12
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 42 19 47
rect 11 40 14 42
rect 16 40 19 42
rect 11 38 19 40
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 57 29 62
rect 21 55 24 57
rect 26 55 29 57
rect 21 38 29 55
rect 31 49 39 66
rect 31 47 34 49
rect 36 47 39 49
rect 31 42 39 47
rect 31 40 34 42
rect 36 40 39 42
rect 31 38 39 40
rect 41 54 47 66
rect 41 52 49 54
rect 41 50 44 52
rect 46 50 49 52
rect 41 38 49 50
rect 51 51 56 54
rect 51 49 58 51
rect 51 47 54 49
rect 56 47 58 49
rect 51 42 58 47
rect 51 40 54 42
rect 56 40 58 42
rect 51 38 58 40
<< alu1 >>
rect -2 67 66 72
rect -2 65 55 67
rect 57 65 66 67
rect -2 64 66 65
rect 33 49 38 51
rect 33 47 34 49
rect 36 47 38 49
rect 53 49 62 51
rect 33 42 38 47
rect 53 47 54 49
rect 56 47 62 49
rect 53 45 62 47
rect 53 42 57 45
rect 9 40 14 42
rect 16 40 34 42
rect 36 40 54 42
rect 56 40 57 42
rect 9 38 57 40
rect 26 24 30 38
rect 35 33 55 34
rect 35 31 37 33
rect 39 31 51 33
rect 53 31 55 33
rect 35 30 55 31
rect 26 22 27 24
rect 29 22 30 24
rect 26 17 30 22
rect 26 15 27 17
rect 29 15 30 17
rect 26 13 30 15
rect 49 22 55 30
rect -2 7 66 8
rect -2 5 5 7
rect 7 5 53 7
rect 55 5 66 7
rect -2 0 66 5
<< ptie >>
rect 3 7 9 24
rect 3 5 5 7
rect 7 5 9 7
rect 51 7 57 24
rect 51 5 53 7
rect 55 5 57 7
rect 3 3 9 5
rect 51 3 57 5
<< ntie >>
rect 51 67 61 69
rect 51 65 55 67
rect 57 65 61 67
rect 51 61 61 65
<< nmos >>
rect 22 10 24 26
rect 32 10 34 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 38 41 66
rect 49 38 51 54
<< polyct1 >>
rect 37 31 39 33
rect 51 31 53 33
<< ndifct0 >>
rect 17 20 19 22
rect 17 12 19 14
rect 37 20 39 22
rect 37 12 39 14
<< ndifct1 >>
rect 27 22 29 24
rect 27 15 29 17
<< ntiect1 >>
rect 55 65 57 67
<< ptiect1 >>
rect 5 5 7 7
rect 53 5 55 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 47 16 49
rect 24 62 26 64
rect 24 55 26 57
rect 44 50 46 52
<< pdifct1 >>
rect 14 40 16 42
rect 34 47 36 49
rect 34 40 36 42
rect 54 47 56 49
rect 54 40 56 42
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 22 62 24 64
rect 26 62 28 64
rect 22 57 28 62
rect 22 55 24 57
rect 26 55 28 57
rect 22 54 28 55
rect 43 52 47 64
rect 13 49 17 51
rect 13 47 14 49
rect 16 47 17 49
rect 13 42 17 47
rect 43 50 44 52
rect 46 50 47 52
rect 43 48 47 50
rect 16 22 20 24
rect 16 20 17 22
rect 19 20 20 22
rect 16 14 20 20
rect 16 12 17 14
rect 19 12 20 14
rect 36 22 40 24
rect 36 20 37 22
rect 39 20 40 22
rect 36 14 40 20
rect 16 8 20 12
rect 36 12 37 14
rect 39 12 40 14
rect 36 8 40 12
<< labels >>
rlabel alu1 12 40 12 40 6 z
rlabel alu1 28 28 28 28 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 32 4 32 4 6 vss
rlabel alu1 44 32 44 32 6 a
rlabel alu1 44 40 44 40 6 z
rlabel alu1 36 44 36 44 6 z
rlabel alu1 32 68 32 68 6 vdd
rlabel alu1 52 28 52 28 6 a
rlabel alu1 52 40 52 40 6 z
rlabel alu1 60 48 60 48 6 z
<< end >>
