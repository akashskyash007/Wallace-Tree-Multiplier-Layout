magic
tech scmos
timestamp 1199543382
<< ab >>
rect 0 0 80 100
<< nwell >>
rect -5 48 85 105
<< pwell >>
rect -5 -5 85 48
<< poly >>
rect 19 94 21 98
rect 27 94 29 98
rect 35 94 37 98
rect 43 94 45 98
rect 55 94 57 98
rect 67 94 69 98
rect 19 53 21 56
rect 17 51 23 53
rect 17 49 19 51
rect 21 49 23 51
rect 11 47 23 49
rect 11 25 13 47
rect 27 43 29 56
rect 35 53 37 56
rect 43 53 45 56
rect 55 53 57 56
rect 67 53 69 56
rect 35 51 39 53
rect 43 51 49 53
rect 55 51 69 53
rect 37 43 39 51
rect 47 43 49 51
rect 57 49 59 51
rect 61 49 63 51
rect 57 47 63 49
rect 27 41 33 43
rect 27 39 29 41
rect 31 39 33 41
rect 23 37 33 39
rect 37 41 43 43
rect 37 39 39 41
rect 41 39 43 41
rect 37 37 43 39
rect 47 41 53 43
rect 47 39 49 41
rect 51 39 53 41
rect 47 37 53 39
rect 23 25 25 37
rect 37 29 39 37
rect 47 29 49 37
rect 57 31 63 33
rect 57 29 59 31
rect 61 29 63 31
rect 33 27 39 29
rect 45 27 49 29
rect 55 27 69 29
rect 33 24 35 27
rect 45 24 47 27
rect 55 24 57 27
rect 67 24 69 27
rect 11 11 13 15
rect 23 11 25 15
rect 33 11 35 15
rect 45 11 47 15
rect 55 2 57 6
rect 67 2 69 6
<< ndif >>
rect 3 15 11 25
rect 13 21 23 25
rect 13 19 17 21
rect 19 19 23 21
rect 13 15 23 19
rect 25 24 30 25
rect 25 15 33 24
rect 35 21 45 24
rect 35 19 39 21
rect 41 19 45 21
rect 35 15 45 19
rect 47 15 55 24
rect 3 11 9 15
rect 3 9 5 11
rect 7 9 9 11
rect 3 7 9 9
rect 27 9 31 15
rect 49 9 55 15
rect 27 7 33 9
rect 27 5 29 7
rect 31 5 33 7
rect 27 3 33 5
rect 47 7 55 9
rect 47 5 49 7
rect 51 6 55 7
rect 57 21 67 24
rect 57 19 61 21
rect 63 19 67 21
rect 57 6 67 19
rect 69 11 77 24
rect 69 9 73 11
rect 75 9 77 11
rect 69 6 77 9
rect 51 5 53 6
rect 47 3 53 5
<< pdif >>
rect 11 85 19 94
rect 7 81 19 85
rect 7 79 9 81
rect 11 79 19 81
rect 7 71 19 79
rect 7 69 9 71
rect 11 69 19 71
rect 7 61 19 69
rect 7 59 9 61
rect 11 59 19 61
rect 7 56 19 59
rect 21 56 27 94
rect 29 56 35 94
rect 37 56 43 94
rect 45 91 55 94
rect 45 89 49 91
rect 51 89 55 91
rect 45 56 55 89
rect 57 81 67 94
rect 57 79 61 81
rect 63 79 67 81
rect 57 71 67 79
rect 57 69 61 71
rect 63 69 67 71
rect 57 61 67 69
rect 57 59 61 61
rect 63 59 67 61
rect 57 56 67 59
rect 69 91 77 94
rect 69 89 73 91
rect 75 89 77 91
rect 69 81 77 89
rect 69 79 73 81
rect 75 79 77 81
rect 69 71 77 79
rect 69 69 73 71
rect 75 69 77 71
rect 69 56 77 69
rect 7 55 13 56
<< alu1 >>
rect -2 91 82 100
rect -2 89 49 91
rect 51 89 73 91
rect 75 89 82 91
rect -2 88 82 89
rect 8 81 12 83
rect 8 79 9 81
rect 11 79 12 81
rect 8 71 12 79
rect 8 69 9 71
rect 11 69 12 71
rect 8 61 12 69
rect 8 59 9 61
rect 11 59 12 61
rect 8 22 12 59
rect 18 51 22 83
rect 18 49 19 51
rect 21 49 22 51
rect 18 27 22 49
rect 28 41 32 83
rect 28 39 29 41
rect 31 39 32 41
rect 28 27 32 39
rect 38 41 42 83
rect 38 39 39 41
rect 41 39 42 41
rect 38 27 42 39
rect 48 41 52 83
rect 58 82 62 83
rect 58 81 65 82
rect 58 79 61 81
rect 63 79 65 81
rect 58 78 65 79
rect 72 81 76 88
rect 72 79 73 81
rect 75 79 76 81
rect 58 72 62 78
rect 58 71 65 72
rect 58 69 61 71
rect 63 69 65 71
rect 58 68 65 69
rect 72 71 76 79
rect 72 69 73 71
rect 75 69 76 71
rect 58 62 62 68
rect 72 67 76 69
rect 68 62 72 63
rect 58 61 72 62
rect 58 59 61 61
rect 63 59 72 61
rect 58 58 72 59
rect 58 57 62 58
rect 48 39 49 41
rect 51 39 52 41
rect 48 37 52 39
rect 58 51 62 53
rect 58 49 59 51
rect 61 49 62 51
rect 58 32 62 49
rect 48 31 62 32
rect 48 29 59 31
rect 61 29 62 31
rect 48 28 62 29
rect 48 22 52 28
rect 58 27 62 28
rect 68 22 72 58
rect 8 21 52 22
rect 8 19 17 21
rect 19 19 39 21
rect 41 19 52 21
rect 8 18 52 19
rect 59 21 72 22
rect 59 19 61 21
rect 63 19 72 21
rect 59 18 72 19
rect 68 17 72 18
rect -2 11 82 12
rect -2 9 5 11
rect 7 9 73 11
rect 75 9 82 11
rect -2 7 82 9
rect -2 5 29 7
rect 31 5 49 7
rect 51 5 82 7
rect -2 0 82 5
<< nmos >>
rect 11 15 13 25
rect 23 15 25 25
rect 33 15 35 24
rect 45 15 47 24
rect 55 6 57 24
rect 67 6 69 24
<< pmos >>
rect 19 56 21 94
rect 27 56 29 94
rect 35 56 37 94
rect 43 56 45 94
rect 55 56 57 94
rect 67 56 69 94
<< polyct1 >>
rect 19 49 21 51
rect 59 49 61 51
rect 29 39 31 41
rect 39 39 41 41
rect 49 39 51 41
rect 59 29 61 31
<< ndifct1 >>
rect 17 19 19 21
rect 39 19 41 21
rect 5 9 7 11
rect 29 5 31 7
rect 49 5 51 7
rect 61 19 63 21
rect 73 9 75 11
<< pdifct1 >>
rect 9 79 11 81
rect 9 69 11 71
rect 9 59 11 61
rect 49 89 51 91
rect 61 79 63 81
rect 61 69 63 71
rect 61 59 63 61
rect 73 89 75 91
rect 73 79 75 81
rect 73 69 75 71
<< labels >>
rlabel alu1 20 55 20 55 6 i1
rlabel alu1 30 55 30 55 6 i0
rlabel alu1 40 6 40 6 6 vss
rlabel alu1 40 55 40 55 6 i2
rlabel alu1 50 60 50 60 6 i3
rlabel alu1 40 94 40 94 6 vdd
rlabel alu1 70 40 70 40 6 q
rlabel alu1 60 70 60 70 6 q
<< end >>
