magic
tech scmos
timestamp 1199203037
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 12 66 14 70
rect 19 66 21 70
rect 26 66 28 70
rect 12 35 14 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 29 21 38
rect 26 35 28 38
rect 26 33 38 35
rect 29 31 34 33
rect 36 31 38 33
rect 29 29 38 31
rect 9 25 11 29
rect 19 27 25 29
rect 19 25 21 27
rect 23 25 25 27
rect 19 23 25 25
rect 19 20 21 23
rect 29 20 31 29
rect 9 11 11 15
rect 19 5 21 10
rect 29 5 31 10
<< ndif >>
rect 4 21 9 25
rect 2 19 9 21
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 20 17 25
rect 11 15 19 20
rect 13 10 19 15
rect 21 17 29 20
rect 21 15 24 17
rect 26 15 29 17
rect 21 10 29 15
rect 31 14 38 20
rect 31 12 34 14
rect 36 12 38 14
rect 31 10 38 12
rect 13 9 17 10
rect 11 7 17 9
rect 11 5 13 7
rect 15 5 17 7
rect 11 3 17 5
<< pdif >>
rect 7 59 12 66
rect 5 57 12 59
rect 5 55 7 57
rect 9 55 12 57
rect 5 50 12 55
rect 5 48 7 50
rect 9 48 12 50
rect 5 46 12 48
rect 7 38 12 46
rect 14 38 19 66
rect 21 38 26 66
rect 28 64 38 66
rect 28 62 34 64
rect 36 62 38 64
rect 28 57 38 62
rect 28 55 34 57
rect 36 55 38 57
rect 28 38 38 55
<< alu1 >>
rect -2 64 42 72
rect 5 57 11 58
rect 5 55 7 57
rect 9 55 11 57
rect 5 51 11 55
rect 2 50 11 51
rect 2 48 7 50
rect 9 48 11 50
rect 2 47 11 48
rect 2 21 6 47
rect 18 43 22 51
rect 34 43 38 51
rect 10 39 22 43
rect 10 33 14 39
rect 26 37 38 43
rect 10 31 11 33
rect 13 31 14 33
rect 10 29 14 31
rect 18 30 22 35
rect 18 27 24 30
rect 18 26 21 27
rect 20 25 21 26
rect 23 26 24 27
rect 23 25 31 26
rect 20 22 31 25
rect 2 19 7 21
rect 2 17 4 19
rect 6 18 7 19
rect 6 17 28 18
rect 2 15 24 17
rect 26 15 28 17
rect 2 14 28 15
rect -2 7 42 8
rect -2 5 13 7
rect 15 5 42 7
rect -2 0 42 5
<< nmos >>
rect 9 15 11 25
rect 19 10 21 20
rect 29 10 31 20
<< pmos >>
rect 12 38 14 66
rect 19 38 21 66
rect 26 38 28 66
<< polyct0 >>
rect 34 31 36 33
<< polyct1 >>
rect 11 31 13 33
rect 21 25 23 27
<< ndifct0 >>
rect 34 12 36 14
<< ndifct1 >>
rect 4 17 6 19
rect 24 15 26 17
rect 13 5 15 7
<< pdifct0 >>
rect 34 62 36 64
rect 34 55 36 57
<< pdifct1 >>
rect 7 55 9 57
rect 7 48 9 50
<< alu0 >>
rect 32 62 34 64
rect 36 62 38 64
rect 32 57 38 62
rect 32 55 34 57
rect 36 55 38 57
rect 32 54 38 55
rect 33 33 37 37
rect 33 31 34 33
rect 36 31 37 33
rect 33 29 37 31
rect 33 14 37 16
rect 33 12 34 14
rect 36 12 37 14
rect 33 8 37 12
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 12 36 12 36 6 c
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 20 16 20 16 6 z
rlabel alu1 20 32 20 32 6 b
rlabel alu1 28 24 28 24 6 b
rlabel alu1 28 40 28 40 6 a
rlabel alu1 20 48 20 48 6 c
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 20 68 20 68 6 vdd
rlabel alu1 36 44 36 44 6 a
<< end >>
