magic
tech scmos
timestamp 1199202397
<< ab >>
rect 0 0 40 72
<< nwell >>
rect -5 32 45 77
<< pwell >>
rect -5 -5 45 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 9 33 31 35
rect 9 31 17 33
rect 19 31 21 33
rect 9 29 21 31
rect 9 26 11 29
rect 19 26 21 29
rect 9 5 11 10
rect 19 5 21 10
<< ndif >>
rect 2 14 9 26
rect 2 12 4 14
rect 6 12 9 14
rect 2 10 9 12
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 17 19 22
rect 11 15 14 17
rect 16 15 19 17
rect 11 10 19 15
rect 21 17 28 26
rect 21 15 24 17
rect 26 15 28 17
rect 21 13 28 15
rect 21 10 27 13
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 64 19 66
rect 11 62 14 64
rect 16 62 19 64
rect 11 57 19 62
rect 11 55 14 57
rect 16 55 19 57
rect 11 38 19 55
rect 21 49 29 66
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 64 38 66
rect 31 62 34 64
rect 36 62 38 64
rect 31 57 38 62
rect 31 55 34 57
rect 36 55 38 57
rect 31 38 38 55
<< alu1 >>
rect -2 64 42 72
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 2 40 4 42
rect 6 40 24 42
rect 26 40 31 42
rect 2 38 31 40
rect 2 26 6 38
rect 15 33 31 34
rect 15 31 17 33
rect 19 31 31 33
rect 15 30 31 31
rect 2 24 17 26
rect 2 22 14 24
rect 16 22 17 24
rect 25 22 31 30
rect 2 21 17 22
rect 13 17 17 21
rect 13 15 14 17
rect 16 15 17 17
rect 13 13 17 15
rect -2 7 42 8
rect -2 5 33 7
rect 35 5 42 7
rect -2 0 42 5
<< ptie >>
rect 31 7 37 9
rect 31 5 33 7
rect 35 5 37 7
rect 31 3 37 5
<< nmos >>
rect 9 10 11 26
rect 19 10 21 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
<< polyct1 >>
rect 17 31 19 33
<< ndifct0 >>
rect 4 12 6 14
rect 24 15 26 17
<< ndifct1 >>
rect 14 22 16 24
rect 14 15 16 17
<< ptiect1 >>
rect 33 5 35 7
<< pdifct0 >>
rect 14 62 16 64
rect 14 55 16 57
rect 24 47 26 49
rect 34 62 36 64
rect 34 55 36 57
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 24 40 26 42
<< alu0 >>
rect 13 62 14 64
rect 16 62 17 64
rect 13 57 17 62
rect 13 55 14 57
rect 16 55 17 57
rect 13 53 17 55
rect 32 62 34 64
rect 36 62 38 64
rect 32 57 38 62
rect 32 55 34 57
rect 36 55 38 57
rect 32 54 38 55
rect 23 49 27 51
rect 23 47 24 49
rect 26 47 27 49
rect 23 42 27 47
rect 3 14 7 16
rect 3 12 4 14
rect 6 12 7 14
rect 22 17 28 18
rect 22 15 24 17
rect 26 15 28 17
rect 3 8 7 12
rect 22 8 28 15
<< labels >>
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 24 12 24 6 z
rlabel alu1 12 40 12 40 6 z
rlabel alu1 20 4 20 4 6 vss
rlabel alu1 20 32 20 32 6 a
rlabel alu1 28 28 28 28 6 a
rlabel alu1 28 40 28 40 6 z
rlabel alu1 20 40 20 40 6 z
rlabel alu1 20 68 20 68 6 vdd
<< end >>
