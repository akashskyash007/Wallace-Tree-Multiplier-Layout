magic
tech scmos
timestamp 1199201767
<< ab >>
rect 0 0 96 72
<< nwell >>
rect -5 32 101 77
<< pwell >>
rect -5 -5 101 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 59 66 61 70
rect 78 57 84 59
rect 78 55 80 57
rect 82 55 84 57
rect 78 53 84 55
rect 71 41 77 43
rect 9 35 11 38
rect 19 35 21 38
rect 9 33 24 35
rect 9 31 20 33
rect 22 31 24 33
rect 29 31 31 40
rect 39 37 41 40
rect 49 37 51 40
rect 38 35 44 37
rect 38 33 40 35
rect 42 33 44 35
rect 38 31 44 33
rect 48 35 55 37
rect 48 33 51 35
rect 53 33 55 35
rect 48 31 55 33
rect 59 35 61 40
rect 71 39 73 41
rect 75 39 77 41
rect 71 37 77 39
rect 59 33 66 35
rect 59 31 62 33
rect 64 31 66 33
rect 9 29 24 31
rect 28 29 34 31
rect 9 26 11 29
rect 19 26 21 29
rect 28 27 30 29
rect 32 27 34 29
rect 9 11 11 15
rect 28 25 35 27
rect 33 22 35 25
rect 40 22 42 31
rect 48 27 50 31
rect 59 27 66 31
rect 47 25 50 27
rect 54 25 66 27
rect 47 22 49 25
rect 54 22 56 25
rect 64 22 66 25
rect 71 22 73 37
rect 82 33 84 53
rect 78 31 84 33
rect 78 22 80 31
rect 88 29 94 31
rect 88 27 90 29
rect 92 27 94 29
rect 85 25 94 27
rect 85 22 87 25
rect 19 5 21 9
rect 33 2 35 6
rect 40 2 42 6
rect 47 2 49 6
rect 54 2 56 6
rect 64 2 66 6
rect 71 2 73 6
rect 78 2 80 6
rect 85 2 87 6
<< ndif >>
rect 2 19 9 26
rect 2 17 4 19
rect 6 17 9 19
rect 2 15 9 17
rect 11 24 19 26
rect 11 22 14 24
rect 16 22 19 24
rect 11 15 19 22
rect 14 9 19 15
rect 21 22 26 26
rect 21 10 33 22
rect 21 9 26 10
rect 23 8 26 9
rect 28 8 33 10
rect 23 6 33 8
rect 35 6 40 22
rect 42 6 47 22
rect 49 6 54 22
rect 56 17 64 22
rect 56 15 59 17
rect 61 15 64 17
rect 56 6 64 15
rect 66 6 71 22
rect 73 6 78 22
rect 80 6 85 22
rect 87 17 94 22
rect 87 15 90 17
rect 92 15 94 17
rect 87 10 94 15
rect 87 8 90 10
rect 92 8 94 10
rect 87 6 94 8
<< pdif >>
rect 2 64 9 66
rect 2 62 4 64
rect 6 62 9 64
rect 2 57 9 62
rect 2 55 4 57
rect 6 55 9 57
rect 2 38 9 55
rect 11 57 19 66
rect 11 55 14 57
rect 16 55 19 57
rect 11 50 19 55
rect 11 48 14 50
rect 16 48 19 50
rect 11 38 19 48
rect 21 64 29 66
rect 21 62 24 64
rect 26 62 29 64
rect 21 56 29 62
rect 21 54 24 56
rect 26 54 29 56
rect 21 40 29 54
rect 31 53 39 66
rect 31 51 34 53
rect 36 51 39 53
rect 31 45 39 51
rect 31 43 34 45
rect 36 43 39 45
rect 31 40 39 43
rect 41 64 49 66
rect 41 62 44 64
rect 46 62 49 64
rect 41 40 49 62
rect 51 57 59 66
rect 51 55 54 57
rect 56 55 59 57
rect 51 40 59 55
rect 61 64 69 66
rect 61 62 64 64
rect 66 62 69 64
rect 61 40 69 62
rect 21 38 27 40
<< alu1 >>
rect -2 67 98 72
rect -2 65 79 67
rect 81 65 89 67
rect 91 65 98 67
rect -2 64 98 65
rect 65 57 87 58
rect 65 55 80 57
rect 82 55 87 57
rect 65 54 87 55
rect 10 43 14 51
rect 65 50 69 54
rect 2 37 14 43
rect 10 26 14 37
rect 42 46 69 50
rect 73 46 87 50
rect 42 36 46 46
rect 73 42 77 46
rect 38 35 46 36
rect 38 33 40 35
rect 42 33 46 35
rect 38 32 46 33
rect 50 41 77 42
rect 50 39 73 41
rect 75 39 77 41
rect 50 38 77 39
rect 81 38 87 42
rect 50 35 54 38
rect 50 33 51 35
rect 53 33 54 35
rect 81 34 86 38
rect 50 31 54 33
rect 60 33 86 34
rect 60 31 62 33
rect 64 31 86 33
rect 10 24 17 26
rect 10 22 14 24
rect 16 22 17 24
rect 10 20 17 22
rect 29 29 33 31
rect 60 30 86 31
rect 29 27 30 29
rect 32 27 33 29
rect 29 26 33 27
rect 90 29 94 31
rect 92 27 94 29
rect 90 26 94 27
rect 29 22 94 26
rect 74 21 94 22
rect 74 13 78 21
rect -2 7 98 8
rect -2 5 5 7
rect 7 5 98 7
rect -2 0 98 5
<< ptie >>
rect 3 7 9 9
rect 3 5 5 7
rect 7 5 9 7
rect 3 3 9 5
<< ntie >>
rect 77 67 93 69
rect 77 65 79 67
rect 81 65 89 67
rect 91 65 93 67
rect 77 63 93 65
<< nmos >>
rect 9 15 11 26
rect 19 9 21 26
rect 33 6 35 22
rect 40 6 42 22
rect 47 6 49 22
rect 54 6 56 22
rect 64 6 66 22
rect 71 6 73 22
rect 78 6 80 22
rect 85 6 87 22
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 40 31 66
rect 39 40 41 66
rect 49 40 51 66
rect 59 40 61 66
<< polyct0 >>
rect 20 31 22 33
<< polyct1 >>
rect 80 55 82 57
rect 40 33 42 35
rect 51 33 53 35
rect 73 39 75 41
rect 62 31 64 33
rect 30 27 32 29
rect 90 27 92 29
<< ndifct0 >>
rect 4 17 6 19
rect 26 8 28 10
rect 59 15 61 17
rect 90 15 92 17
rect 90 8 92 10
<< ndifct1 >>
rect 14 22 16 24
<< ntiect1 >>
rect 79 65 81 67
rect 89 65 91 67
<< ptiect1 >>
rect 5 5 7 7
<< pdifct0 >>
rect 4 62 6 64
rect 4 55 6 57
rect 14 55 16 57
rect 14 48 16 50
rect 24 62 26 64
rect 24 54 26 56
rect 34 51 36 53
rect 34 43 36 45
rect 44 62 46 64
rect 54 55 56 57
rect 64 62 66 64
<< alu0 >>
rect 2 62 4 64
rect 6 62 8 64
rect 2 57 8 62
rect 23 62 24 64
rect 26 62 27 64
rect 2 55 4 57
rect 6 55 8 57
rect 2 54 8 55
rect 13 57 17 59
rect 13 55 14 57
rect 16 55 17 57
rect 13 51 17 55
rect 23 56 27 62
rect 42 62 44 64
rect 46 62 48 64
rect 42 61 48 62
rect 62 62 64 64
rect 66 62 68 64
rect 62 61 68 62
rect 23 54 24 56
rect 26 54 27 56
rect 23 52 27 54
rect 33 57 58 58
rect 33 55 54 57
rect 56 55 58 57
rect 33 54 58 55
rect 33 53 37 54
rect 14 50 17 51
rect 16 48 17 50
rect 14 46 17 48
rect 33 51 34 53
rect 36 51 37 53
rect 33 45 37 51
rect 21 43 34 45
rect 36 43 37 45
rect 21 41 37 43
rect 21 34 25 41
rect 18 33 25 34
rect 18 31 20 33
rect 22 31 25 33
rect 18 30 25 31
rect 3 19 7 21
rect 3 17 4 19
rect 6 17 7 19
rect 3 8 7 17
rect 21 18 25 30
rect 89 26 90 31
rect 21 17 63 18
rect 21 15 59 17
rect 61 15 63 17
rect 21 14 63 15
rect 88 17 94 18
rect 88 15 90 17
rect 92 15 94 17
rect 24 10 30 11
rect 24 8 26 10
rect 28 8 30 10
rect 88 10 94 15
rect 88 8 90 10
rect 92 8 94 10
<< labels >>
rlabel alu0 23 29 23 29 6 zn
rlabel alu0 35 49 35 49 6 zn
rlabel alu0 42 16 42 16 6 zn
rlabel alu0 45 56 45 56 6 zn
rlabel alu1 12 36 12 36 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 48 4 48 4 6 vss
rlabel alu1 36 24 36 24 6 a
rlabel alu1 52 24 52 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 44 40 44 40 6 b
rlabel alu1 52 48 52 48 6 b
rlabel alu1 48 68 48 68 6 vdd
rlabel alu1 60 24 60 24 6 a
rlabel alu1 68 24 68 24 6 a
rlabel alu1 76 20 76 20 6 a
rlabel alu1 76 32 76 32 6 d
rlabel alu1 68 32 68 32 6 d
rlabel alu1 60 40 60 40 6 c
rlabel alu1 68 40 68 40 6 c
rlabel alu1 60 48 60 48 6 b
rlabel alu1 76 48 76 48 6 c
rlabel alu1 76 56 76 56 6 b
rlabel alu1 68 56 68 56 6 b
rlabel alu1 92 24 92 24 6 a
rlabel alu1 84 24 84 24 6 a
rlabel alu1 84 40 84 40 6 d
rlabel alu1 84 48 84 48 6 c
rlabel alu1 84 56 84 56 6 b
<< end >>
