magic
tech scmos
timestamp 1199469243
<< ab >>
rect 0 0 50 100
<< nwell >>
rect -5 48 55 105
<< pwell >>
rect -5 -5 55 48
<< poly >>
rect 13 94 15 98
rect 25 94 27 98
rect 37 94 39 98
rect 13 43 15 56
rect 25 43 27 56
rect 37 53 39 56
rect 32 51 39 53
rect 32 49 34 51
rect 36 49 39 51
rect 32 47 39 49
rect 13 41 27 43
rect 13 39 23 41
rect 25 39 27 41
rect 13 37 27 39
rect 13 34 15 37
rect 25 34 27 37
rect 37 34 39 47
rect 13 11 15 15
rect 25 10 27 15
rect 37 10 39 15
<< ndif >>
rect 4 21 13 34
rect 4 19 7 21
rect 9 19 13 21
rect 4 15 13 19
rect 15 31 25 34
rect 15 29 19 31
rect 21 29 25 31
rect 15 21 25 29
rect 15 19 19 21
rect 21 19 25 21
rect 15 15 25 19
rect 27 31 37 34
rect 27 29 31 31
rect 33 29 37 31
rect 27 21 37 29
rect 27 19 31 21
rect 33 19 37 21
rect 27 15 37 19
rect 39 32 47 34
rect 39 30 43 32
rect 45 30 47 32
rect 39 24 47 30
rect 39 22 43 24
rect 45 22 47 24
rect 39 20 47 22
rect 39 15 44 20
<< pdif >>
rect 4 91 13 94
rect 4 89 7 91
rect 9 89 13 91
rect 4 81 13 89
rect 4 79 7 81
rect 9 79 13 81
rect 4 71 13 79
rect 4 69 7 71
rect 9 69 13 71
rect 4 56 13 69
rect 15 71 25 94
rect 15 69 19 71
rect 21 69 25 71
rect 15 61 25 69
rect 15 59 19 61
rect 21 59 25 61
rect 15 56 25 59
rect 27 91 37 94
rect 27 89 31 91
rect 33 89 37 91
rect 27 81 37 89
rect 27 79 31 81
rect 33 79 37 81
rect 27 56 37 79
rect 39 70 44 94
rect 39 68 47 70
rect 39 66 43 68
rect 45 66 47 68
rect 39 60 47 66
rect 39 58 43 60
rect 45 58 47 60
rect 39 56 47 58
<< alu1 >>
rect -2 91 52 100
rect -2 89 7 91
rect 9 89 31 91
rect 33 89 52 91
rect -2 88 52 89
rect 6 81 10 88
rect 6 79 7 81
rect 9 79 10 81
rect 6 71 10 79
rect 30 81 34 88
rect 30 79 31 81
rect 33 79 34 81
rect 30 77 34 79
rect 6 69 7 71
rect 9 69 10 71
rect 6 67 10 69
rect 18 71 22 73
rect 18 69 19 71
rect 21 69 22 71
rect 18 63 22 69
rect 8 61 22 63
rect 8 59 19 61
rect 21 59 22 61
rect 8 57 22 59
rect 8 33 12 57
rect 28 52 32 73
rect 42 68 46 70
rect 42 66 43 68
rect 45 66 46 68
rect 42 60 46 66
rect 42 58 43 60
rect 45 58 46 60
rect 17 51 38 52
rect 17 49 34 51
rect 36 49 38 51
rect 17 48 38 49
rect 42 42 46 58
rect 21 41 46 42
rect 21 39 23 41
rect 25 39 46 41
rect 21 38 46 39
rect 8 31 22 33
rect 8 29 19 31
rect 21 29 22 31
rect 8 27 22 29
rect 6 21 10 23
rect 6 19 7 21
rect 9 19 10 21
rect 6 12 10 19
rect 18 21 22 27
rect 18 19 19 21
rect 21 19 22 21
rect 18 17 22 19
rect 30 31 34 33
rect 30 29 31 31
rect 33 29 34 31
rect 30 21 34 29
rect 30 19 31 21
rect 33 19 34 21
rect 42 32 46 38
rect 42 30 43 32
rect 45 30 46 32
rect 42 24 46 30
rect 42 22 43 24
rect 45 22 46 24
rect 42 20 46 22
rect 30 12 34 19
rect -2 7 52 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 52 7
rect -2 0 52 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< nmos >>
rect 13 15 15 34
rect 25 15 27 34
rect 37 15 39 34
<< pmos >>
rect 13 56 15 94
rect 25 56 27 94
rect 37 56 39 94
<< polyct1 >>
rect 34 49 36 51
rect 23 39 25 41
<< ndifct1 >>
rect 7 19 9 21
rect 19 29 21 31
rect 19 19 21 21
rect 31 29 33 31
rect 31 19 33 21
rect 43 30 45 32
rect 43 22 45 24
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 7 89 9 91
rect 7 79 9 81
rect 7 69 9 71
rect 19 69 21 71
rect 19 59 21 61
rect 31 89 33 91
rect 31 79 33 81
rect 43 66 45 68
rect 43 58 45 60
<< labels >>
rlabel polyct1 24 40 24 40 6 an
rlabel ndifct1 44 23 44 23 6 an
rlabel ndifct1 44 31 44 31 6 an
rlabel pdifct1 44 59 44 59 6 an
rlabel pdifct1 44 67 44 67 6 an
rlabel alu1 20 25 20 25 6 z
rlabel alu1 10 45 10 45 6 z
rlabel alu1 20 50 20 50 6 a
rlabel alu1 20 65 20 65 6 z
rlabel alu1 25 6 25 6 6 vss
rlabel alu1 30 60 30 60 6 a
rlabel alu1 25 94 25 94 6 vdd
<< end >>
