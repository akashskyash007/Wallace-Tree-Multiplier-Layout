magic
tech scmos
timestamp 1199542175
<< ab >>
rect 0 0 130 100
<< nwell >>
rect -2 48 132 104
<< pwell >>
rect -2 -4 132 48
<< poly >>
rect 27 95 29 98
rect 39 95 41 98
rect 51 95 53 98
rect 59 95 61 98
rect 71 95 73 98
rect 83 95 85 98
rect 91 95 93 98
rect 115 95 117 98
rect 15 69 17 72
rect 15 53 17 55
rect 7 51 17 53
rect 7 49 9 51
rect 11 49 17 51
rect 7 47 17 49
rect 15 37 17 47
rect 27 53 29 75
rect 39 73 41 75
rect 33 71 41 73
rect 33 69 35 71
rect 37 69 41 71
rect 33 67 41 69
rect 27 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 15 26 17 29
rect 27 23 29 47
rect 39 41 41 67
rect 51 63 53 75
rect 47 61 53 63
rect 47 59 49 61
rect 51 59 53 61
rect 47 57 53 59
rect 47 51 53 53
rect 59 51 61 75
rect 71 73 73 75
rect 83 73 85 75
rect 47 49 49 51
rect 51 49 61 51
rect 47 47 53 49
rect 39 39 53 41
rect 33 31 41 33
rect 33 29 35 31
rect 37 29 41 31
rect 33 27 41 29
rect 39 23 41 27
rect 51 23 53 39
rect 59 23 61 49
rect 69 71 73 73
rect 79 71 85 73
rect 69 33 71 71
rect 79 53 81 71
rect 91 63 93 75
rect 103 69 105 72
rect 85 61 93 63
rect 85 59 87 61
rect 89 59 93 61
rect 85 57 93 59
rect 75 51 81 53
rect 103 51 105 55
rect 75 49 77 51
rect 79 49 105 51
rect 75 47 81 49
rect 79 39 81 47
rect 65 31 71 33
rect 65 29 67 31
rect 69 29 71 31
rect 65 27 71 29
rect 75 37 81 39
rect 85 41 93 43
rect 85 39 87 41
rect 89 39 93 41
rect 85 37 93 39
rect 75 23 77 37
rect 81 31 87 33
rect 81 29 83 31
rect 85 29 87 31
rect 81 27 87 29
rect 71 21 77 23
rect 71 19 73 21
rect 83 19 85 27
rect 91 19 93 37
rect 103 35 105 49
rect 115 43 117 55
rect 111 41 117 43
rect 111 39 113 41
rect 115 39 117 41
rect 111 37 117 39
rect 115 35 117 37
rect 103 26 105 29
rect 27 8 29 11
rect 39 8 41 11
rect 51 8 53 11
rect 59 8 61 11
rect 115 12 117 15
rect 71 4 73 7
rect 83 4 85 7
rect 91 4 93 7
<< ndif >>
rect 7 29 15 37
rect 17 33 25 37
rect 17 31 21 33
rect 23 31 25 33
rect 17 29 25 31
rect 7 21 13 29
rect 43 31 49 33
rect 43 29 45 31
rect 47 29 49 31
rect 43 23 49 29
rect 7 19 9 21
rect 11 19 13 21
rect 7 17 13 19
rect 19 21 27 23
rect 19 19 21 21
rect 23 19 27 21
rect 19 11 27 19
rect 29 11 39 23
rect 41 11 51 23
rect 53 11 59 23
rect 61 21 69 23
rect 61 19 65 21
rect 67 19 69 21
rect 95 33 103 35
rect 95 31 97 33
rect 99 31 103 33
rect 95 29 103 31
rect 105 29 115 35
rect 95 21 101 23
rect 95 19 97 21
rect 99 19 101 21
rect 61 11 71 19
rect 63 7 71 11
rect 73 11 83 19
rect 73 9 77 11
rect 79 9 83 11
rect 73 7 83 9
rect 85 7 91 19
rect 93 7 101 19
rect 107 15 115 29
rect 117 31 125 35
rect 117 29 121 31
rect 123 29 125 31
rect 117 21 125 29
rect 117 19 121 21
rect 123 19 125 21
rect 117 15 125 19
rect 107 11 113 15
rect 107 9 109 11
rect 111 9 113 11
rect 107 7 113 9
<< pdif >>
rect 7 81 13 83
rect 7 79 9 81
rect 11 79 13 81
rect 7 69 13 79
rect 19 81 27 95
rect 19 79 21 81
rect 23 79 27 81
rect 19 75 27 79
rect 29 75 39 95
rect 41 75 51 95
rect 53 75 59 95
rect 61 81 71 95
rect 61 79 65 81
rect 67 79 71 81
rect 61 75 71 79
rect 73 91 83 95
rect 73 89 77 91
rect 79 89 83 91
rect 73 75 83 89
rect 85 75 91 95
rect 93 81 101 95
rect 93 79 97 81
rect 99 79 101 81
rect 93 75 101 79
rect 107 93 115 95
rect 107 91 109 93
rect 111 91 115 93
rect 7 55 15 69
rect 17 61 25 69
rect 17 59 21 61
rect 23 59 25 61
rect 17 55 25 59
rect 43 71 49 75
rect 43 69 45 71
rect 47 69 49 71
rect 43 67 49 69
rect 107 69 115 91
rect 95 61 103 69
rect 95 59 97 61
rect 99 59 103 61
rect 95 55 103 59
rect 105 55 115 69
rect 117 81 125 95
rect 117 79 121 81
rect 123 79 125 81
rect 117 71 125 79
rect 117 69 121 71
rect 123 69 125 71
rect 117 61 125 69
rect 117 59 121 61
rect 123 59 125 61
rect 117 55 125 59
<< alu1 >>
rect -2 93 132 100
rect -2 91 109 93
rect 111 91 132 93
rect -2 89 77 91
rect 79 89 132 91
rect -2 88 132 89
rect 8 81 12 88
rect 8 79 9 81
rect 11 79 12 81
rect 8 78 12 79
rect 20 81 68 82
rect 20 79 21 81
rect 23 79 65 81
rect 67 79 68 81
rect 20 78 68 79
rect 96 81 100 82
rect 96 79 97 81
rect 99 79 100 81
rect 96 72 100 79
rect 118 81 124 82
rect 118 79 121 81
rect 123 79 124 81
rect 118 78 124 79
rect 118 72 122 78
rect 8 71 12 72
rect 34 71 38 72
rect 8 69 35 71
rect 37 69 38 71
rect 8 51 12 69
rect 34 68 38 69
rect 44 71 111 72
rect 118 71 124 72
rect 44 69 45 71
rect 47 69 112 71
rect 44 68 112 69
rect 20 61 52 62
rect 8 49 9 51
rect 11 49 12 51
rect 8 28 12 49
rect 18 59 21 61
rect 23 59 49 61
rect 51 59 52 61
rect 18 58 52 59
rect 18 34 22 58
rect 28 51 32 52
rect 28 49 29 51
rect 31 49 32 51
rect 28 41 32 49
rect 39 51 52 52
rect 39 49 49 51
rect 51 49 52 51
rect 39 48 52 49
rect 58 42 62 68
rect 55 41 62 42
rect 54 39 62 41
rect 68 52 72 62
rect 78 61 90 62
rect 78 59 87 61
rect 89 59 90 61
rect 78 58 90 59
rect 96 61 100 62
rect 96 59 97 61
rect 99 59 102 61
rect 96 58 102 59
rect 86 52 90 58
rect 68 51 80 52
rect 68 49 77 51
rect 79 49 80 51
rect 68 48 80 49
rect 86 48 92 52
rect 54 38 61 39
rect 68 38 72 48
rect 86 42 90 48
rect 78 41 90 42
rect 78 39 87 41
rect 89 39 90 41
rect 78 38 90 39
rect 18 33 24 34
rect 18 31 21 33
rect 23 32 24 33
rect 54 32 58 38
rect 98 34 102 58
rect 96 33 102 34
rect 96 32 97 33
rect 23 31 38 32
rect 20 30 35 31
rect 21 29 35 30
rect 37 29 38 31
rect 21 28 38 29
rect 44 31 58 32
rect 44 29 45 31
rect 47 29 58 31
rect 66 31 97 32
rect 99 31 102 33
rect 66 29 67 31
rect 69 29 83 31
rect 85 29 102 31
rect 108 42 112 68
rect 118 69 121 71
rect 123 69 124 71
rect 118 68 124 69
rect 118 62 122 68
rect 118 61 124 62
rect 118 59 121 61
rect 123 59 124 61
rect 118 58 124 59
rect 118 52 122 58
rect 118 48 126 52
rect 108 41 116 42
rect 108 39 113 41
rect 115 39 116 41
rect 108 38 116 39
rect 44 28 57 29
rect 66 28 101 29
rect 108 22 112 38
rect 122 32 126 48
rect 8 21 12 22
rect 8 19 9 21
rect 11 19 12 21
rect 8 12 12 19
rect 20 21 68 22
rect 20 19 21 21
rect 23 19 65 21
rect 67 19 68 21
rect 20 18 68 19
rect 96 21 112 22
rect 96 19 97 21
rect 99 19 112 21
rect 118 31 126 32
rect 118 29 121 31
rect 123 29 126 31
rect 118 28 126 29
rect 118 22 122 28
rect 118 21 124 22
rect 118 19 121 21
rect 123 19 124 21
rect 96 18 111 19
rect 118 18 124 19
rect -2 11 132 12
rect -2 9 77 11
rect 79 9 109 11
rect 111 9 132 11
rect -2 0 132 9
<< nmos >>
rect 15 29 17 37
rect 27 11 29 23
rect 39 11 41 23
rect 51 11 53 23
rect 59 11 61 23
rect 103 29 105 35
rect 71 7 73 19
rect 83 7 85 19
rect 91 7 93 19
rect 115 15 117 35
<< pmos >>
rect 27 75 29 95
rect 39 75 41 95
rect 51 75 53 95
rect 59 75 61 95
rect 71 75 73 95
rect 83 75 85 95
rect 91 75 93 95
rect 15 55 17 69
rect 103 55 105 69
rect 115 55 117 95
<< polyct1 >>
rect 9 49 11 51
rect 35 69 37 71
rect 29 49 31 51
rect 49 59 51 61
rect 49 49 51 51
rect 35 29 37 31
rect 87 59 89 61
rect 77 49 79 51
rect 67 29 69 31
rect 87 39 89 41
rect 83 29 85 31
rect 113 39 115 41
<< ndifct1 >>
rect 21 31 23 33
rect 45 29 47 31
rect 9 19 11 21
rect 21 19 23 21
rect 65 19 67 21
rect 97 31 99 33
rect 97 19 99 21
rect 77 9 79 11
rect 121 29 123 31
rect 121 19 123 21
rect 109 9 111 11
<< pdifct1 >>
rect 9 79 11 81
rect 21 79 23 81
rect 65 79 67 81
rect 77 89 79 91
rect 97 79 99 81
rect 109 91 111 93
rect 21 59 23 61
rect 45 69 47 71
rect 97 59 99 61
rect 121 79 123 81
rect 121 69 123 71
rect 121 59 123 61
<< labels >>
rlabel polyct1 10 50 10 50 6 cmd1
rlabel polyct1 30 50 30 50 6 i2
rlabel alu1 65 6 65 6 6 vss
rlabel polyct1 50 50 50 50 6 i1
rlabel alu1 70 50 70 50 6 cmd0
rlabel alu1 65 94 65 94 6 vdd
rlabel alu1 80 40 80 40 6 i0
rlabel alu1 90 50 90 50 6 i0
rlabel alu1 80 60 80 60 6 i0
rlabel alu1 120 25 120 25 6 q
rlabel alu1 120 65 120 65 6 q
<< end >>
