magic
tech scmos
timestamp 1199203647
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 22 70 24 74
rect 32 70 34 74
rect 42 70 44 74
rect 52 70 54 74
rect 2 61 8 63
rect 2 59 4 61
rect 6 59 8 61
rect 2 57 11 59
rect 9 54 11 57
rect 61 54 63 58
rect 9 40 11 43
rect 22 40 24 43
rect 9 38 24 40
rect 32 39 34 43
rect 42 39 44 43
rect 52 40 54 43
rect 61 40 63 43
rect 9 30 11 38
rect 19 30 21 38
rect 32 37 38 39
rect 32 35 34 37
rect 36 35 38 37
rect 26 30 28 34
rect 32 33 38 35
rect 42 37 48 39
rect 52 38 63 40
rect 42 35 44 37
rect 46 35 48 37
rect 42 33 48 35
rect 36 30 38 33
rect 43 30 45 33
rect 54 30 56 38
rect 9 19 11 24
rect 54 18 56 24
rect 64 20 70 22
rect 64 18 66 20
rect 68 18 70 20
rect 19 13 21 18
rect 26 10 28 18
rect 36 14 38 18
rect 43 14 45 18
rect 54 16 70 18
rect 54 10 56 16
rect 26 8 56 10
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 24 9 26
rect 11 28 19 30
rect 11 26 14 28
rect 16 26 19 28
rect 11 24 19 26
rect 13 18 19 24
rect 21 18 26 30
rect 28 22 36 30
rect 28 20 31 22
rect 33 20 36 22
rect 28 18 36 20
rect 38 18 43 30
rect 45 24 54 30
rect 56 28 63 30
rect 56 26 59 28
rect 61 26 63 28
rect 56 24 63 26
rect 45 22 52 24
rect 45 20 48 22
rect 50 20 52 22
rect 45 18 52 20
<< pdif >>
rect 13 66 22 70
rect 13 64 17 66
rect 19 64 22 66
rect 13 54 22 64
rect 4 49 9 54
rect 2 47 9 49
rect 2 45 4 47
rect 6 45 9 47
rect 2 43 9 45
rect 11 43 22 54
rect 24 62 32 70
rect 24 60 27 62
rect 29 60 32 62
rect 24 43 32 60
rect 34 47 42 70
rect 34 45 37 47
rect 39 45 42 47
rect 34 43 42 45
rect 44 62 52 70
rect 44 60 47 62
rect 49 60 52 62
rect 44 43 52 60
rect 54 64 61 70
rect 54 62 57 64
rect 59 62 61 64
rect 54 60 61 62
rect 54 54 59 60
rect 54 43 61 54
rect 63 49 68 54
rect 63 47 70 49
rect 63 45 66 47
rect 68 45 70 47
rect 63 43 70 45
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 61 7 63
rect 2 59 4 61
rect 6 59 7 61
rect 2 58 7 59
rect 2 54 14 58
rect 10 49 14 54
rect 35 47 41 48
rect 35 46 37 47
rect 26 45 37 46
rect 39 45 41 47
rect 26 42 41 45
rect 26 23 30 42
rect 26 22 35 23
rect 26 20 31 22
rect 33 20 35 22
rect 26 19 35 20
rect 66 22 70 31
rect 57 20 70 22
rect 57 18 66 20
rect 68 18 70 20
rect 57 17 70 18
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 9 24 11 30
rect 19 18 21 30
rect 26 18 28 30
rect 36 18 38 30
rect 43 18 45 30
rect 54 24 56 30
<< pmos >>
rect 9 43 11 54
rect 22 43 24 70
rect 32 43 34 70
rect 42 43 44 70
rect 52 43 54 70
rect 61 43 63 54
<< polyct0 >>
rect 34 35 36 37
rect 44 35 46 37
<< polyct1 >>
rect 4 59 6 61
rect 66 18 68 20
<< ndifct0 >>
rect 4 26 6 28
rect 14 26 16 28
rect 59 26 61 28
rect 48 20 50 22
<< ndifct1 >>
rect 31 20 33 22
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 17 64 19 66
rect 4 45 6 47
rect 27 60 29 62
rect 47 60 49 62
rect 57 62 59 64
rect 66 45 68 47
<< pdifct1 >>
rect 37 45 39 47
<< alu0 >>
rect 16 66 20 68
rect 16 64 17 66
rect 19 64 20 66
rect 16 62 20 64
rect 56 64 60 68
rect 25 62 51 63
rect 25 60 27 62
rect 29 60 47 62
rect 49 60 51 62
rect 56 62 57 64
rect 59 62 60 64
rect 56 60 60 62
rect 25 59 51 60
rect 18 51 49 55
rect 3 47 7 49
rect 3 45 4 47
rect 6 45 7 47
rect 18 45 22 51
rect 3 41 22 45
rect 3 28 7 41
rect 3 26 4 28
rect 6 26 7 28
rect 3 24 7 26
rect 13 28 17 30
rect 13 26 14 28
rect 16 26 17 28
rect 13 12 17 26
rect 33 37 38 39
rect 45 38 49 51
rect 33 35 34 37
rect 36 35 38 37
rect 33 33 38 35
rect 42 37 49 38
rect 42 35 44 37
rect 46 35 49 37
rect 42 34 49 35
rect 59 47 70 48
rect 59 45 66 47
rect 68 45 70 47
rect 59 44 70 45
rect 34 31 38 33
rect 59 31 63 44
rect 34 28 63 31
rect 34 27 59 28
rect 57 26 59 27
rect 61 26 63 28
rect 57 25 63 26
rect 46 22 52 23
rect 46 20 48 22
rect 50 20 52 22
rect 46 12 52 20
<< labels >>
rlabel alu0 5 36 5 36 6 an
rlabel alu0 36 33 36 33 6 bn
rlabel alu0 47 44 47 44 6 an
rlabel alu0 38 61 38 61 6 n3
rlabel alu0 61 36 61 36 6 bn
rlabel alu0 64 46 64 46 6 bn
rlabel alu1 12 52 12 52 6 a
rlabel alu1 4 60 4 60 6 a
rlabel alu1 28 32 28 32 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 44 36 44 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 20 60 20 6 b
rlabel alu1 68 24 68 24 6 b
<< end >>
