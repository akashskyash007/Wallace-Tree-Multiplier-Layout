magic
tech scmos
timestamp 1199203010
<< ab >>
rect 0 0 64 80
<< nwell >>
rect -5 36 69 88
<< pwell >>
rect -5 -8 69 36
<< poly >>
rect 11 70 13 74
rect 18 70 20 74
rect 25 70 27 74
rect 35 70 37 74
rect 42 70 44 74
rect 49 70 51 74
rect 11 31 13 42
rect 18 39 20 42
rect 25 39 27 42
rect 35 39 37 42
rect 18 36 21 39
rect 25 37 37 39
rect 19 31 21 36
rect 35 31 37 37
rect 9 29 15 31
rect 9 27 11 29
rect 13 27 15 29
rect 9 25 15 27
rect 19 29 25 31
rect 19 27 21 29
rect 23 27 25 29
rect 19 25 25 27
rect 31 29 37 31
rect 31 27 33 29
rect 35 27 37 29
rect 42 33 44 42
rect 49 39 51 42
rect 49 37 58 39
rect 52 35 54 37
rect 56 35 58 37
rect 52 33 58 35
rect 42 31 48 33
rect 42 29 44 31
rect 46 29 48 31
rect 42 27 48 29
rect 31 25 37 27
rect 9 22 11 25
rect 21 22 23 25
rect 31 22 33 25
rect 9 7 11 12
rect 21 7 23 12
rect 31 7 33 12
<< ndif >>
rect 2 20 9 22
rect 2 18 4 20
rect 6 18 9 20
rect 2 16 9 18
rect 4 12 9 16
rect 11 12 21 22
rect 23 20 31 22
rect 23 18 26 20
rect 28 18 31 20
rect 23 12 31 18
rect 33 12 42 22
rect 13 11 19 12
rect 13 9 15 11
rect 17 9 19 11
rect 13 7 19 9
rect 35 11 42 12
rect 35 9 37 11
rect 39 9 42 11
rect 35 7 42 9
<< pdif >>
rect 4 68 11 70
rect 4 66 6 68
rect 8 66 11 68
rect 4 61 11 66
rect 4 59 6 61
rect 8 59 11 61
rect 4 42 11 59
rect 13 42 18 70
rect 20 42 25 70
rect 27 61 35 70
rect 27 59 30 61
rect 32 59 35 61
rect 27 54 35 59
rect 27 52 30 54
rect 32 52 35 54
rect 27 42 35 52
rect 37 42 42 70
rect 44 42 49 70
rect 51 68 58 70
rect 51 66 54 68
rect 56 66 58 68
rect 51 61 58 66
rect 51 59 54 61
rect 56 59 58 61
rect 51 42 58 59
<< alu1 >>
rect -2 81 66 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 66 81
rect -2 68 66 79
rect 2 52 30 54
rect 32 52 39 54
rect 2 50 39 52
rect 2 21 6 50
rect 10 42 55 46
rect 10 29 14 42
rect 51 38 55 42
rect 10 27 11 29
rect 13 27 14 29
rect 10 25 14 27
rect 18 34 47 38
rect 51 37 58 38
rect 51 35 54 37
rect 56 35 58 37
rect 51 34 58 35
rect 18 29 24 34
rect 43 31 47 34
rect 18 27 21 29
rect 23 27 24 29
rect 18 25 24 27
rect 31 29 39 30
rect 31 27 33 29
rect 35 27 39 29
rect 31 26 39 27
rect 43 29 44 31
rect 46 30 47 31
rect 46 29 55 30
rect 43 26 55 29
rect 34 22 39 26
rect 2 20 30 21
rect 2 18 4 20
rect 6 18 26 20
rect 28 18 30 20
rect 2 17 30 18
rect 34 17 47 22
rect -2 11 66 12
rect -2 9 15 11
rect 17 9 37 11
rect 39 9 66 11
rect -2 1 66 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 66 1
rect -2 -2 66 -1
<< ptie >>
rect 0 1 64 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 64 1
rect 0 -3 64 -1
<< ntie >>
rect 0 81 64 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 64 81
rect 0 77 64 79
<< nmos >>
rect 9 12 11 22
rect 21 12 23 22
rect 31 12 33 22
<< pmos >>
rect 11 42 13 70
rect 18 42 20 70
rect 25 42 27 70
rect 35 42 37 70
rect 42 42 44 70
rect 49 42 51 70
<< polyct1 >>
rect 11 27 13 29
rect 21 27 23 29
rect 33 27 35 29
rect 54 35 56 37
rect 44 29 46 31
<< ndifct1 >>
rect 4 18 6 20
rect 26 18 28 20
rect 15 9 17 11
rect 37 9 39 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
<< pdifct0 >>
rect 6 66 8 68
rect 6 59 8 61
rect 30 59 32 61
rect 54 66 56 68
rect 54 59 56 61
<< pdifct1 >>
rect 30 52 32 54
<< alu0 >>
rect 4 66 6 68
rect 8 66 10 68
rect 4 61 10 66
rect 52 66 54 68
rect 56 66 58 68
rect 4 59 6 61
rect 8 59 10 61
rect 4 58 10 59
rect 29 61 33 63
rect 29 59 30 61
rect 32 59 33 61
rect 29 54 33 59
rect 52 61 58 66
rect 52 59 54 61
rect 56 59 58 61
rect 52 58 58 59
<< labels >>
rlabel alu1 12 32 12 32 6 a
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 36 28 36 6 b
rlabel alu1 20 28 20 28 6 b
rlabel alu1 20 44 20 44 6 a
rlabel alu1 28 44 28 44 6 a
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 32 6 32 6 6 vss
rlabel alu1 44 20 44 20 6 c
rlabel alu1 36 24 36 24 6 c
rlabel alu1 36 36 36 36 6 b
rlabel alu1 44 36 44 36 6 b
rlabel alu1 44 44 44 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 36 52 36 52 6 z
rlabel alu1 32 74 32 74 6 vdd
rlabel alu1 52 28 52 28 6 b
rlabel alu1 52 44 52 44 6 a
<< end >>
