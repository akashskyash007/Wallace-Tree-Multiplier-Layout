magic
tech scmos
timestamp 1199544137
<< ab >>
rect 0 0 130 100
<< nwell >>
rect -2 48 132 104
<< pwell >>
rect -2 -4 132 48
<< poly >>
rect 17 95 19 98
rect 29 95 31 98
rect 41 95 43 98
rect 53 95 55 98
rect 65 95 67 98
rect 93 85 95 88
rect 105 85 107 88
rect 117 85 119 88
rect 65 63 67 75
rect 75 65 81 67
rect 75 63 77 65
rect 79 63 81 65
rect 93 63 95 65
rect 65 61 71 63
rect 75 61 95 63
rect 65 59 67 61
rect 69 59 71 61
rect 65 57 71 59
rect 105 57 107 65
rect 117 63 119 65
rect 111 61 119 63
rect 111 59 113 61
rect 115 59 119 61
rect 111 57 119 59
rect 65 55 107 57
rect 17 47 19 55
rect 29 47 31 55
rect 41 47 43 55
rect 53 47 55 55
rect 95 53 97 55
rect 99 53 101 55
rect 95 51 101 53
rect 121 47 127 49
rect 17 45 123 47
rect 125 45 127 47
rect 121 43 127 45
rect 17 37 91 39
rect 17 25 19 37
rect 29 25 31 37
rect 41 25 43 37
rect 53 25 55 37
rect 85 35 87 37
rect 89 35 91 37
rect 85 33 91 35
rect 95 37 119 39
rect 95 35 97 37
rect 99 35 101 37
rect 95 33 101 35
rect 59 31 67 33
rect 59 29 61 31
rect 63 29 67 31
rect 59 27 67 29
rect 75 31 81 33
rect 75 29 77 31
rect 79 29 81 31
rect 105 31 113 33
rect 105 29 109 31
rect 111 29 113 31
rect 75 27 95 29
rect 65 25 67 27
rect 93 25 95 27
rect 105 27 113 29
rect 105 25 107 27
rect 117 25 119 37
rect 65 12 67 15
rect 93 12 95 15
rect 105 12 107 15
rect 117 12 119 15
rect 17 2 19 5
rect 29 2 31 5
rect 41 2 43 5
rect 53 2 55 5
<< ndif >>
rect 9 21 17 25
rect 9 19 11 21
rect 13 19 17 21
rect 9 11 17 19
rect 9 9 11 11
rect 13 9 17 11
rect 9 5 17 9
rect 19 21 29 25
rect 19 19 23 21
rect 25 19 29 21
rect 19 5 29 19
rect 31 21 41 25
rect 31 19 35 21
rect 37 19 41 21
rect 31 11 41 19
rect 31 9 35 11
rect 37 9 41 11
rect 31 5 41 9
rect 43 21 53 25
rect 43 19 47 21
rect 49 19 53 21
rect 43 5 53 19
rect 55 15 65 25
rect 67 21 75 25
rect 67 19 71 21
rect 73 19 75 21
rect 67 15 75 19
rect 85 21 93 25
rect 85 19 87 21
rect 89 19 93 21
rect 85 15 93 19
rect 95 15 105 25
rect 107 21 117 25
rect 107 19 111 21
rect 113 19 117 21
rect 107 15 117 19
rect 119 21 127 25
rect 119 19 123 21
rect 125 19 127 21
rect 119 15 127 19
rect 55 11 63 15
rect 55 9 59 11
rect 61 9 63 11
rect 97 11 103 15
rect 97 9 99 11
rect 101 9 103 11
rect 55 5 63 9
rect 97 7 103 9
<< pdif >>
rect 9 91 17 95
rect 9 89 11 91
rect 13 89 17 91
rect 9 81 17 89
rect 9 79 11 81
rect 13 79 17 81
rect 9 71 17 79
rect 9 69 11 71
rect 13 69 17 71
rect 9 61 17 69
rect 9 59 11 61
rect 13 59 17 61
rect 9 55 17 59
rect 19 81 29 95
rect 19 79 23 81
rect 25 79 29 81
rect 19 71 29 79
rect 19 69 23 71
rect 25 69 29 71
rect 19 61 29 69
rect 19 59 23 61
rect 25 59 29 61
rect 19 55 29 59
rect 31 91 41 95
rect 31 89 35 91
rect 37 89 41 91
rect 31 81 41 89
rect 31 79 35 81
rect 37 79 41 81
rect 31 71 41 79
rect 31 69 35 71
rect 37 69 41 71
rect 31 61 41 69
rect 31 59 35 61
rect 37 59 41 61
rect 31 55 41 59
rect 43 81 53 95
rect 43 79 47 81
rect 49 79 53 81
rect 43 71 53 79
rect 43 69 47 71
rect 49 69 53 71
rect 43 61 53 69
rect 43 59 47 61
rect 49 59 53 61
rect 43 55 53 59
rect 55 91 65 95
rect 55 89 59 91
rect 61 89 65 91
rect 55 75 65 89
rect 67 81 75 95
rect 109 91 115 93
rect 109 89 111 91
rect 113 89 115 91
rect 109 85 115 89
rect 67 79 71 81
rect 73 79 75 81
rect 67 75 75 79
rect 85 81 93 85
rect 85 79 87 81
rect 89 79 93 81
rect 55 55 63 75
rect 85 71 93 79
rect 85 69 87 71
rect 89 69 93 71
rect 85 65 93 69
rect 95 81 105 85
rect 95 79 99 81
rect 101 79 105 81
rect 95 71 105 79
rect 95 69 99 71
rect 101 69 105 71
rect 95 65 105 69
rect 107 65 117 85
rect 119 81 127 85
rect 119 79 123 81
rect 125 79 127 81
rect 119 71 127 79
rect 119 69 123 71
rect 125 69 127 71
rect 119 65 127 69
<< alu1 >>
rect -2 95 132 100
rect -2 93 83 95
rect 85 93 99 95
rect 101 93 132 95
rect -2 91 132 93
rect -2 89 11 91
rect 13 89 35 91
rect 37 89 59 91
rect 61 89 111 91
rect 113 89 132 91
rect -2 88 132 89
rect 10 81 14 88
rect 10 79 11 81
rect 13 79 14 81
rect 10 71 14 79
rect 10 69 11 71
rect 13 69 14 71
rect 10 61 14 69
rect 10 59 11 61
rect 13 59 14 61
rect 10 58 14 59
rect 22 81 26 82
rect 22 79 23 81
rect 25 79 26 81
rect 22 71 26 79
rect 22 69 23 71
rect 25 69 26 71
rect 22 61 26 69
rect 22 59 23 61
rect 25 59 26 61
rect 22 44 26 59
rect 34 81 38 88
rect 34 79 35 81
rect 37 79 38 81
rect 34 71 38 79
rect 46 81 52 82
rect 46 79 47 81
rect 49 79 52 81
rect 46 78 52 79
rect 48 72 52 78
rect 34 69 35 71
rect 37 69 38 71
rect 34 61 38 69
rect 46 71 52 72
rect 46 69 47 71
rect 49 69 52 71
rect 46 68 52 69
rect 48 62 52 68
rect 34 59 35 61
rect 37 59 38 61
rect 34 58 38 59
rect 46 61 52 62
rect 46 59 47 61
rect 49 59 52 61
rect 46 58 52 59
rect 48 44 52 58
rect 22 40 52 44
rect 10 21 14 22
rect 10 19 11 21
rect 13 19 14 21
rect 10 12 14 19
rect 22 21 26 40
rect 48 22 52 40
rect 22 19 23 21
rect 25 19 26 21
rect 22 18 26 19
rect 34 21 38 22
rect 34 19 35 21
rect 37 19 38 21
rect 34 12 38 19
rect 46 21 52 22
rect 46 19 47 21
rect 49 19 52 21
rect 46 18 52 19
rect 58 62 62 82
rect 70 81 79 82
rect 70 79 71 81
rect 73 79 79 81
rect 70 78 79 79
rect 86 81 90 82
rect 86 79 87 81
rect 89 79 90 81
rect 86 78 90 79
rect 98 81 102 82
rect 122 81 126 82
rect 98 79 99 81
rect 101 79 123 81
rect 125 79 126 81
rect 98 78 102 79
rect 122 78 126 79
rect 77 66 79 78
rect 87 72 89 78
rect 99 72 101 78
rect 123 72 125 78
rect 86 71 90 72
rect 86 69 87 71
rect 89 69 90 71
rect 86 68 90 69
rect 98 71 102 72
rect 98 69 99 71
rect 101 69 102 71
rect 98 68 102 69
rect 76 65 80 66
rect 76 63 77 65
rect 79 63 80 65
rect 76 62 80 63
rect 58 61 70 62
rect 58 59 67 61
rect 69 59 70 61
rect 58 58 70 59
rect 58 32 62 58
rect 77 32 79 62
rect 87 38 89 68
rect 108 62 112 72
rect 122 71 126 72
rect 122 69 123 71
rect 125 69 126 71
rect 122 68 126 69
rect 108 61 116 62
rect 108 59 113 61
rect 115 59 116 61
rect 108 58 116 59
rect 96 55 100 56
rect 96 53 97 55
rect 99 53 100 55
rect 96 52 100 53
rect 97 38 99 52
rect 86 37 90 38
rect 86 35 87 37
rect 89 35 90 37
rect 86 34 90 35
rect 96 37 100 38
rect 96 35 97 37
rect 99 35 100 37
rect 96 34 100 35
rect 58 31 64 32
rect 58 29 61 31
rect 63 29 64 31
rect 58 28 64 29
rect 76 31 80 32
rect 76 29 77 31
rect 79 29 80 31
rect 76 28 80 29
rect 58 18 62 28
rect 77 22 79 28
rect 87 22 89 34
rect 108 31 112 58
rect 123 48 125 68
rect 122 47 126 48
rect 122 45 123 47
rect 125 45 126 47
rect 122 44 126 45
rect 108 29 109 31
rect 111 29 112 31
rect 108 28 112 29
rect 123 22 125 44
rect 70 21 79 22
rect 70 19 71 21
rect 73 19 79 21
rect 70 18 79 19
rect 86 21 90 22
rect 110 21 114 22
rect 86 19 87 21
rect 89 19 111 21
rect 113 19 114 21
rect 86 18 90 19
rect 110 18 114 19
rect 122 21 126 22
rect 122 19 123 21
rect 125 19 126 21
rect 122 18 126 19
rect -2 11 132 12
rect -2 9 11 11
rect 13 9 35 11
rect 37 9 59 11
rect 61 9 99 11
rect 101 9 132 11
rect -2 7 132 9
rect -2 5 71 7
rect 73 5 87 7
rect 89 5 111 7
rect 113 5 123 7
rect 125 5 132 7
rect -2 0 132 5
<< ptie >>
rect 69 7 91 9
rect 109 7 127 9
rect 69 5 71 7
rect 73 5 87 7
rect 89 5 91 7
rect 69 3 91 5
rect 109 5 111 7
rect 113 5 123 7
rect 125 5 127 7
rect 109 3 127 5
<< ntie >>
rect 81 95 103 97
rect 81 93 83 95
rect 85 93 99 95
rect 101 93 103 95
rect 81 91 103 93
<< nmos >>
rect 17 5 19 25
rect 29 5 31 25
rect 41 5 43 25
rect 53 5 55 25
rect 65 15 67 25
rect 93 15 95 25
rect 105 15 107 25
rect 117 15 119 25
<< pmos >>
rect 17 55 19 95
rect 29 55 31 95
rect 41 55 43 95
rect 53 55 55 95
rect 65 75 67 95
rect 93 65 95 85
rect 105 65 107 85
rect 117 65 119 85
<< polyct1 >>
rect 77 63 79 65
rect 67 59 69 61
rect 113 59 115 61
rect 97 53 99 55
rect 123 45 125 47
rect 87 35 89 37
rect 97 35 99 37
rect 61 29 63 31
rect 77 29 79 31
rect 109 29 111 31
<< ndifct1 >>
rect 11 19 13 21
rect 11 9 13 11
rect 23 19 25 21
rect 35 19 37 21
rect 35 9 37 11
rect 47 19 49 21
rect 71 19 73 21
rect 87 19 89 21
rect 111 19 113 21
rect 123 19 125 21
rect 59 9 61 11
rect 99 9 101 11
<< ntiect1 >>
rect 83 93 85 95
rect 99 93 101 95
<< ptiect1 >>
rect 71 5 73 7
rect 87 5 89 7
rect 111 5 113 7
rect 123 5 125 7
<< pdifct1 >>
rect 11 89 13 91
rect 11 79 13 81
rect 11 69 13 71
rect 11 59 13 61
rect 23 79 25 81
rect 23 69 25 71
rect 23 59 25 61
rect 35 89 37 91
rect 35 79 37 81
rect 35 69 37 71
rect 35 59 37 61
rect 47 79 49 81
rect 47 69 49 71
rect 47 59 49 61
rect 59 89 61 91
rect 111 89 113 91
rect 71 79 73 81
rect 87 79 89 81
rect 87 69 89 71
rect 99 79 101 81
rect 99 69 101 71
rect 123 79 125 81
rect 123 69 125 71
<< labels >>
rlabel alu1 65 6 65 6 6 vss
rlabel alu1 50 50 50 50 6 q
rlabel alu1 60 50 60 50 6 cmd
rlabel alu1 65 94 65 94 6 vdd
rlabel alu1 110 50 110 50 6 i
<< end >>
