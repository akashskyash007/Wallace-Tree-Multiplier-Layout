magic
tech scmos
timestamp 1199203629
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 29 72 53 74
rect 9 63 11 68
rect 19 63 21 68
rect 29 63 31 72
rect 41 60 43 65
rect 51 63 53 72
rect 51 61 57 63
rect 9 44 11 47
rect 9 42 15 44
rect 9 40 11 42
rect 13 40 15 42
rect 9 38 15 40
rect 19 39 21 47
rect 10 28 12 38
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 34 25 35
rect 17 32 25 34
rect 17 28 19 32
rect 29 30 31 47
rect 51 59 53 61
rect 55 59 57 61
rect 51 57 57 59
rect 57 45 63 47
rect 41 41 43 44
rect 57 43 59 45
rect 61 43 63 45
rect 57 41 63 43
rect 39 39 63 41
rect 39 30 41 39
rect 49 30 51 35
rect 59 30 61 39
rect 10 12 12 17
rect 17 12 19 17
rect 29 14 31 24
rect 39 18 41 22
rect 49 14 51 22
rect 59 19 61 24
rect 29 12 51 14
<< ndif >>
rect 24 28 29 30
rect 5 23 10 28
rect 3 21 10 23
rect 3 19 5 21
rect 7 19 10 21
rect 3 17 10 19
rect 12 17 17 28
rect 19 24 29 28
rect 31 28 39 30
rect 31 26 34 28
rect 36 26 39 28
rect 31 24 39 26
rect 19 17 27 24
rect 21 11 27 17
rect 34 22 39 24
rect 41 27 49 30
rect 41 25 44 27
rect 46 25 49 27
rect 41 22 49 25
rect 51 28 59 30
rect 51 26 54 28
rect 56 26 59 28
rect 51 24 59 26
rect 61 28 68 30
rect 61 26 64 28
rect 66 26 68 28
rect 61 24 68 26
rect 51 22 56 24
rect 21 9 23 11
rect 25 9 27 11
rect 21 7 27 9
<< pdif >>
rect 33 68 39 70
rect 33 66 35 68
rect 37 66 39 68
rect 33 63 39 66
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 57 9 59
rect 4 47 9 57
rect 11 53 19 63
rect 11 51 14 53
rect 16 51 19 53
rect 11 47 19 51
rect 21 51 29 63
rect 21 49 24 51
rect 26 49 29 51
rect 21 47 29 49
rect 31 60 39 63
rect 31 47 41 60
rect 33 44 41 47
rect 43 50 48 60
rect 43 48 50 50
rect 43 46 46 48
rect 48 46 50 48
rect 43 44 50 46
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 49 61 63 62
rect 49 59 53 61
rect 55 59 63 61
rect 49 58 63 59
rect 2 53 18 54
rect 2 51 14 53
rect 16 51 18 53
rect 2 50 18 51
rect 2 22 6 50
rect 57 50 63 58
rect 57 45 70 46
rect 57 43 59 45
rect 61 43 70 45
rect 57 42 70 43
rect 43 27 47 29
rect 43 25 44 27
rect 46 25 47 27
rect 43 22 47 25
rect 66 33 70 42
rect 2 21 47 22
rect 2 19 5 21
rect 7 19 47 21
rect 2 18 47 19
rect -2 11 74 12
rect -2 9 23 11
rect 25 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 10 17 12 28
rect 17 17 19 28
rect 29 24 31 30
rect 39 22 41 30
rect 49 22 51 30
rect 59 24 61 30
<< pmos >>
rect 9 47 11 63
rect 19 47 21 63
rect 29 47 31 63
rect 41 44 43 60
<< polyct0 >>
rect 11 40 13 42
rect 21 35 23 37
<< polyct1 >>
rect 53 59 55 61
rect 59 43 61 45
<< ndifct0 >>
rect 34 26 36 28
rect 54 26 56 28
rect 64 26 66 28
<< ndifct1 >>
rect 5 19 7 21
rect 44 25 46 27
rect 23 9 25 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 35 66 37 68
rect 4 59 6 61
rect 24 49 26 51
rect 46 46 48 48
<< pdifct1 >>
rect 14 51 16 53
<< alu0 >>
rect 33 66 35 68
rect 37 66 39 68
rect 33 65 39 66
rect 2 61 37 62
rect 2 59 4 61
rect 6 59 37 61
rect 2 58 37 59
rect 23 51 27 53
rect 23 49 24 51
rect 26 49 27 51
rect 23 46 27 49
rect 11 44 27 46
rect 10 42 27 44
rect 10 40 11 42
rect 13 40 15 42
rect 10 38 15 40
rect 33 38 37 58
rect 45 48 49 50
rect 45 46 46 48
rect 48 46 49 48
rect 45 38 49 46
rect 11 30 15 38
rect 19 37 57 38
rect 19 35 21 37
rect 23 35 57 37
rect 19 34 57 35
rect 11 28 38 30
rect 11 26 34 28
rect 36 26 38 28
rect 32 25 38 26
rect 53 28 57 34
rect 53 26 54 28
rect 56 26 57 28
rect 53 24 57 26
rect 63 28 67 30
rect 63 26 64 28
rect 66 26 67 28
rect 63 12 67 26
<< labels >>
rlabel alu0 13 36 13 36 6 bn
rlabel alu0 25 47 25 47 6 bn
rlabel alu0 24 28 24 28 6 bn
rlabel alu0 47 42 47 42 6 an
rlabel alu0 19 60 19 60 6 an
rlabel alu0 55 31 55 31 6 an
rlabel alu0 38 36 38 36 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 52 60 52 60 6 b
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 68 36 68 36 6 a
rlabel polyct1 60 44 60 44 6 a
rlabel alu1 60 56 60 56 6 b
<< end >>
