magic
tech scmos
timestamp 1199468916
<< ab >>
rect 0 0 60 100
<< nwell >>
rect -2 48 62 104
<< pwell >>
rect -2 -4 62 48
<< poly >>
rect 11 80 13 85
rect 23 83 25 88
rect 35 83 37 88
rect 47 83 49 88
rect 11 44 13 60
rect 23 53 25 67
rect 35 63 37 67
rect 35 61 43 63
rect 35 60 39 61
rect 37 59 39 60
rect 41 59 43 61
rect 37 57 43 59
rect 23 51 33 53
rect 27 49 29 51
rect 31 49 33 51
rect 27 47 33 49
rect 11 42 23 44
rect 15 40 19 42
rect 21 40 23 42
rect 15 38 23 40
rect 15 33 17 38
rect 29 33 31 47
rect 37 33 39 57
rect 47 42 49 67
rect 47 40 53 42
rect 47 39 49 40
rect 45 38 49 39
rect 51 38 53 40
rect 45 36 53 38
rect 45 33 47 36
rect 15 18 17 23
rect 29 12 31 17
rect 37 12 39 17
rect 45 12 47 17
<< ndif >>
rect 7 31 15 33
rect 7 29 9 31
rect 11 29 15 31
rect 7 27 15 29
rect 10 23 15 27
rect 17 23 29 33
rect 19 21 29 23
rect 19 19 21 21
rect 23 19 29 21
rect 19 17 29 19
rect 31 17 37 33
rect 39 17 45 33
rect 47 23 52 33
rect 47 21 55 23
rect 47 19 51 21
rect 53 19 55 21
rect 47 17 55 19
<< pdif >>
rect 15 91 21 93
rect 39 91 45 93
rect 15 89 17 91
rect 19 89 21 91
rect 15 83 21 89
rect 39 89 41 91
rect 43 89 45 91
rect 39 83 45 89
rect 15 80 23 83
rect 6 74 11 80
rect 3 72 11 74
rect 3 70 5 72
rect 7 70 11 72
rect 3 64 11 70
rect 3 62 5 64
rect 7 62 11 64
rect 3 60 11 62
rect 13 67 23 80
rect 25 81 35 83
rect 25 79 29 81
rect 31 79 35 81
rect 25 67 35 79
rect 37 67 47 83
rect 49 81 57 83
rect 49 79 53 81
rect 55 79 57 81
rect 49 77 57 79
rect 49 67 54 77
rect 13 60 21 67
<< alu1 >>
rect -2 95 62 100
rect -2 93 29 95
rect 31 93 62 95
rect -2 91 62 93
rect -2 89 17 91
rect 19 89 41 91
rect 43 89 62 91
rect -2 88 62 89
rect 18 81 57 82
rect 18 79 29 81
rect 31 79 53 81
rect 55 79 57 81
rect 18 78 57 79
rect 3 72 12 73
rect 3 70 5 72
rect 7 70 12 72
rect 3 69 12 70
rect 8 65 12 69
rect 3 64 12 65
rect 3 62 5 64
rect 7 62 12 64
rect 3 61 12 62
rect 8 33 12 61
rect 18 42 22 78
rect 28 68 53 73
rect 28 51 32 68
rect 28 49 29 51
rect 31 49 32 51
rect 28 47 32 49
rect 38 61 53 63
rect 38 59 39 61
rect 41 59 53 61
rect 38 58 53 59
rect 18 40 19 42
rect 21 40 32 42
rect 18 38 32 40
rect 8 31 22 33
rect 8 29 9 31
rect 11 29 22 31
rect 8 27 22 29
rect 20 21 24 23
rect 20 19 21 21
rect 23 19 24 21
rect 20 12 24 19
rect 28 22 32 38
rect 38 37 42 58
rect 48 40 52 53
rect 48 38 49 40
rect 51 38 52 40
rect 48 32 52 38
rect 37 27 52 32
rect 28 21 55 22
rect 28 19 51 21
rect 53 19 55 21
rect 28 18 55 19
rect -2 7 62 12
rect -2 5 9 7
rect 11 5 19 7
rect 21 5 62 7
rect -2 0 62 5
<< ptie >>
rect 7 7 23 9
rect 7 5 9 7
rect 11 5 19 7
rect 21 5 23 7
rect 7 3 23 5
<< ntie >>
rect 27 95 33 97
rect 27 93 29 95
rect 31 93 33 95
rect 27 91 33 93
<< nmos >>
rect 15 23 17 33
rect 29 17 31 33
rect 37 17 39 33
rect 45 17 47 33
<< pmos >>
rect 11 60 13 80
rect 23 67 25 83
rect 35 67 37 83
rect 47 67 49 83
<< polyct1 >>
rect 39 59 41 61
rect 29 49 31 51
rect 19 40 21 42
rect 49 38 51 40
<< ndifct1 >>
rect 9 29 11 31
rect 21 19 23 21
rect 51 19 53 21
<< ntiect1 >>
rect 29 93 31 95
<< ptiect1 >>
rect 9 5 11 7
rect 19 5 21 7
<< pdifct1 >>
rect 17 89 19 91
rect 41 89 43 91
rect 5 70 7 72
rect 5 62 7 64
rect 29 79 31 81
rect 53 79 55 81
<< labels >>
rlabel alu1 10 50 10 50 6 z
rlabel alu1 20 30 20 30 6 z
rlabel alu1 30 6 30 6 6 vss
rlabel alu1 25 40 25 40 6 zn
rlabel alu1 40 30 40 30 6 c
rlabel alu1 40 50 40 50 6 b
rlabel alu1 30 60 30 60 6 a
rlabel alu1 40 70 40 70 6 a
rlabel ntiect1 30 94 30 94 6 vdd
rlabel alu1 41 20 41 20 6 zn
rlabel alu1 50 40 50 40 6 c
rlabel alu1 50 70 50 70 6 a
rlabel alu1 50 60 50 60 6 b
rlabel alu1 37 80 37 80 6 zn
<< end >>
