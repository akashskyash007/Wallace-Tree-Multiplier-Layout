magic
tech scmos
timestamp 1199203267
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 9 70 11 74
rect 29 72 55 74
rect 22 64 24 69
rect 29 64 31 72
rect 36 64 38 68
rect 46 61 48 66
rect 53 61 55 72
rect 60 61 62 65
rect 9 39 11 42
rect 22 39 24 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 9 30 11 33
rect 20 22 22 33
rect 29 31 31 42
rect 36 39 38 42
rect 46 39 48 42
rect 36 37 48 39
rect 53 37 55 42
rect 60 39 62 42
rect 60 37 67 39
rect 44 31 48 37
rect 60 35 63 37
rect 65 35 67 37
rect 60 33 67 35
rect 29 29 39 31
rect 29 27 35 29
rect 37 27 39 29
rect 29 25 39 27
rect 44 29 50 31
rect 44 27 46 29
rect 48 27 50 29
rect 44 25 50 27
rect 30 22 32 25
rect 44 22 46 25
rect 9 11 11 16
rect 20 9 22 14
rect 30 9 32 14
rect 44 9 46 14
<< ndif >>
rect 2 28 9 30
rect 2 26 4 28
rect 6 26 9 28
rect 2 21 9 26
rect 2 19 4 21
rect 6 19 9 21
rect 2 16 9 19
rect 11 22 18 30
rect 11 19 20 22
rect 11 17 15 19
rect 17 17 20 19
rect 11 16 20 17
rect 13 14 20 16
rect 22 20 30 22
rect 22 18 25 20
rect 27 18 30 20
rect 22 14 30 18
rect 32 14 44 22
rect 46 20 53 22
rect 46 18 49 20
rect 51 18 53 20
rect 46 16 53 18
rect 46 14 51 16
rect 34 11 42 14
rect 34 9 37 11
rect 39 9 42 11
rect 34 7 42 9
<< pdif >>
rect 4 55 9 70
rect 2 53 9 55
rect 2 51 4 53
rect 6 51 9 53
rect 2 46 9 51
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 68 20 70
rect 11 66 16 68
rect 18 66 20 68
rect 11 64 20 66
rect 11 61 22 64
rect 11 59 16 61
rect 18 59 22 61
rect 11 42 22 59
rect 24 42 29 64
rect 31 42 36 64
rect 38 61 43 64
rect 38 59 46 61
rect 38 57 41 59
rect 43 57 46 59
rect 38 52 46 57
rect 38 50 41 52
rect 43 50 46 52
rect 38 42 46 50
rect 48 42 53 61
rect 55 42 60 61
rect 62 59 70 61
rect 62 57 65 59
rect 67 57 70 59
rect 62 52 70 57
rect 62 50 65 52
rect 67 50 70 52
rect 62 42 70 50
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 53 14 55
rect 2 51 4 53
rect 6 51 14 53
rect 2 49 14 51
rect 2 46 6 49
rect 2 44 4 46
rect 2 30 6 44
rect 26 42 63 46
rect 26 39 30 42
rect 2 28 7 30
rect 2 26 4 28
rect 6 26 7 28
rect 2 21 7 26
rect 20 37 30 39
rect 57 38 63 42
rect 20 35 21 37
rect 23 35 30 37
rect 20 33 30 35
rect 34 34 47 38
rect 57 37 67 38
rect 57 35 63 37
rect 65 35 67 37
rect 57 34 67 35
rect 34 29 38 34
rect 34 27 35 29
rect 37 27 38 29
rect 34 25 38 27
rect 44 29 63 30
rect 44 27 46 29
rect 48 27 63 29
rect 44 26 63 27
rect 2 19 4 21
rect 6 19 7 21
rect 2 17 7 19
rect 57 18 63 26
rect -2 11 74 12
rect -2 9 37 11
rect 39 9 74 11
rect -2 1 74 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 9 16 11 30
rect 20 14 22 22
rect 30 14 32 22
rect 44 14 46 22
<< pmos >>
rect 9 42 11 70
rect 22 42 24 64
rect 29 42 31 64
rect 36 42 38 64
rect 46 42 48 61
rect 53 42 55 61
rect 60 42 62 61
<< polyct0 >>
rect 11 35 13 37
<< polyct1 >>
rect 21 35 23 37
rect 63 35 65 37
rect 35 27 37 29
rect 46 27 48 29
<< ndifct0 >>
rect 15 17 17 19
rect 25 18 27 20
rect 49 18 51 20
<< ndifct1 >>
rect 4 26 6 28
rect 4 19 6 21
rect 37 9 39 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 16 66 18 68
rect 16 59 18 61
rect 41 57 43 59
rect 41 50 43 52
rect 65 57 67 59
rect 65 50 67 52
<< pdifct1 >>
rect 4 51 6 53
rect 4 44 6 46
<< alu0 >>
rect 14 66 16 68
rect 18 66 20 68
rect 14 61 20 66
rect 14 59 16 61
rect 18 59 20 61
rect 14 58 20 59
rect 39 59 45 60
rect 39 57 41 59
rect 43 57 45 59
rect 39 53 45 57
rect 18 52 45 53
rect 18 50 41 52
rect 43 50 45 52
rect 18 49 45 50
rect 63 59 69 68
rect 63 57 65 59
rect 67 57 69 59
rect 63 52 69 57
rect 63 50 65 52
rect 67 50 69 52
rect 63 49 69 50
rect 6 42 7 49
rect 18 46 22 49
rect 10 42 22 46
rect 10 37 14 42
rect 10 35 11 37
rect 13 35 14 37
rect 10 29 14 35
rect 10 25 27 29
rect 23 21 27 25
rect 23 20 53 21
rect 13 19 19 20
rect 13 17 15 19
rect 17 17 19 19
rect 23 18 25 20
rect 27 18 49 20
rect 51 18 53 20
rect 23 17 53 18
rect 13 12 19 17
<< labels >>
rlabel alu0 12 35 12 35 6 zn
rlabel alu0 38 19 38 19 6 zn
rlabel alu0 31 51 31 51 6 zn
rlabel alu0 42 54 42 54 6 zn
rlabel alu1 4 36 4 36 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 28 36 28 36 6 a
rlabel alu1 36 6 36 6 6 vss
rlabel polyct1 36 28 36 28 6 b
rlabel alu1 44 36 44 36 6 b
rlabel alu1 52 28 52 28 6 c
rlabel alu1 44 44 44 44 6 a
rlabel alu1 52 44 52 44 6 a
rlabel alu1 36 44 36 44 6 a
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 60 24 60 24 6 c
rlabel alu1 60 40 60 40 6 a
<< end >>
