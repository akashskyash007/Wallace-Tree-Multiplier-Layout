magic
tech scmos
timestamp 1199202582
<< ab >>
rect 0 0 112 80
<< nwell >>
rect -5 36 117 88
<< pwell >>
rect -5 -8 117 36
<< poly >>
rect 9 68 11 73
rect 19 68 21 73
rect 29 68 31 73
rect 39 68 41 73
rect 49 68 51 73
rect 59 68 61 73
rect 69 60 71 65
rect 79 60 81 65
rect 91 64 93 69
rect 101 64 103 69
rect 9 39 11 42
rect 19 39 21 42
rect 29 39 31 42
rect 39 39 41 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 31 39
rect 19 35 27 37
rect 29 35 31 37
rect 19 33 31 35
rect 35 37 41 39
rect 35 35 37 37
rect 39 35 41 37
rect 49 35 51 42
rect 59 39 61 42
rect 69 39 71 42
rect 59 37 71 39
rect 59 35 61 37
rect 63 35 71 37
rect 79 39 81 42
rect 91 39 93 42
rect 101 39 103 42
rect 79 37 87 39
rect 79 35 83 37
rect 85 35 87 37
rect 35 33 54 35
rect 12 30 14 33
rect 19 30 21 33
rect 29 30 31 33
rect 36 30 38 33
rect 52 30 54 33
rect 59 33 71 35
rect 59 30 61 33
rect 69 30 71 33
rect 76 33 87 35
rect 91 37 103 39
rect 91 35 99 37
rect 101 35 103 37
rect 91 33 103 35
rect 76 30 78 33
rect 91 30 93 33
rect 101 30 103 33
rect 91 14 93 19
rect 101 15 103 19
rect 12 6 14 10
rect 19 6 21 10
rect 29 6 31 10
rect 36 6 38 10
rect 52 6 54 10
rect 59 6 61 10
rect 69 6 71 10
rect 76 6 78 10
<< ndif >>
rect 4 14 12 30
rect 4 12 7 14
rect 9 12 12 14
rect 4 10 12 12
rect 14 10 19 30
rect 21 21 29 30
rect 21 19 24 21
rect 26 19 29 21
rect 21 10 29 19
rect 31 10 36 30
rect 38 14 52 30
rect 38 12 44 14
rect 46 12 52 14
rect 38 10 52 12
rect 54 10 59 30
rect 61 21 69 30
rect 61 19 64 21
rect 66 19 69 21
rect 61 10 69 19
rect 71 10 76 30
rect 78 21 91 30
rect 78 19 83 21
rect 85 19 91 21
rect 93 28 101 30
rect 93 26 96 28
rect 98 26 101 28
rect 93 19 101 26
rect 103 23 110 30
rect 103 21 106 23
rect 108 21 110 23
rect 103 19 110 21
rect 78 14 89 19
rect 78 12 83 14
rect 85 12 89 14
rect 78 10 89 12
<< pdif >>
rect 2 66 9 68
rect 2 64 4 66
rect 6 64 9 66
rect 2 42 9 64
rect 11 60 19 68
rect 11 58 14 60
rect 16 58 19 60
rect 11 53 19 58
rect 11 51 14 53
rect 16 51 19 53
rect 11 42 19 51
rect 21 66 29 68
rect 21 64 24 66
rect 26 64 29 66
rect 21 42 29 64
rect 31 61 39 68
rect 31 59 34 61
rect 36 59 39 61
rect 31 53 39 59
rect 31 51 34 53
rect 36 51 39 53
rect 31 42 39 51
rect 41 66 49 68
rect 41 64 44 66
rect 46 64 49 66
rect 41 42 49 64
rect 51 53 59 68
rect 51 51 54 53
rect 56 51 59 53
rect 51 46 59 51
rect 51 44 54 46
rect 56 44 59 46
rect 51 42 59 44
rect 61 60 67 68
rect 83 60 91 64
rect 61 58 69 60
rect 61 56 64 58
rect 66 56 69 58
rect 61 42 69 56
rect 71 53 79 60
rect 71 51 74 53
rect 76 51 79 53
rect 71 46 79 51
rect 71 44 74 46
rect 76 44 79 46
rect 71 42 79 44
rect 81 58 91 60
rect 81 56 84 58
rect 86 56 91 58
rect 81 42 91 56
rect 93 53 101 64
rect 93 51 96 53
rect 98 51 101 53
rect 93 46 101 51
rect 93 44 96 46
rect 98 44 101 46
rect 93 42 101 44
rect 103 62 110 64
rect 103 60 106 62
rect 108 60 110 62
rect 103 42 110 60
<< alu1 >>
rect -2 81 114 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 114 81
rect -2 68 114 79
rect 2 54 15 55
rect 33 61 38 63
rect 33 59 34 61
rect 36 59 38 61
rect 33 54 38 59
rect 2 53 58 54
rect 2 51 14 53
rect 16 51 34 53
rect 36 51 54 53
rect 56 51 58 53
rect 2 50 58 51
rect 2 22 6 50
rect 53 46 58 50
rect 73 53 78 55
rect 73 51 74 53
rect 76 51 78 53
rect 73 46 78 51
rect 25 42 49 46
rect 53 44 54 46
rect 56 44 74 46
rect 76 44 78 46
rect 53 42 78 44
rect 25 37 31 42
rect 45 38 49 42
rect 25 35 27 37
rect 29 35 31 37
rect 25 34 31 35
rect 45 37 71 38
rect 45 35 61 37
rect 63 35 71 37
rect 45 34 71 35
rect 106 38 110 55
rect 97 37 110 38
rect 97 35 99 37
rect 101 35 110 37
rect 97 34 110 35
rect 2 21 71 22
rect 2 19 24 21
rect 26 19 64 21
rect 66 19 71 21
rect 2 18 71 19
rect -2 1 114 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 114 1
rect -2 -2 114 -1
<< ptie >>
rect 0 1 112 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 75 1
rect 77 -1 83 1
rect 85 -1 91 1
rect 93 -1 99 1
rect 101 -1 107 1
rect 109 -1 112 1
rect 0 -3 112 -1
<< ntie >>
rect 0 81 112 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 75 81
rect 77 79 83 81
rect 85 79 91 81
rect 93 79 99 81
rect 101 79 107 81
rect 109 79 112 81
rect 0 77 112 79
<< nmos >>
rect 12 10 14 30
rect 19 10 21 30
rect 29 10 31 30
rect 36 10 38 30
rect 52 10 54 30
rect 59 10 61 30
rect 69 10 71 30
rect 76 10 78 30
rect 91 19 93 30
rect 101 19 103 30
<< pmos >>
rect 9 42 11 68
rect 19 42 21 68
rect 29 42 31 68
rect 39 42 41 68
rect 49 42 51 68
rect 59 42 61 68
rect 69 42 71 60
rect 79 42 81 60
rect 91 42 93 64
rect 101 42 103 64
<< polyct0 >>
rect 11 35 13 37
rect 37 35 39 37
rect 83 35 85 37
<< polyct1 >>
rect 27 35 29 37
rect 61 35 63 37
rect 99 35 101 37
<< ndifct0 >>
rect 7 12 9 14
rect 44 12 46 14
rect 83 19 85 21
rect 96 26 98 28
rect 106 21 108 23
rect 83 12 85 14
<< ndifct1 >>
rect 24 19 26 21
rect 64 19 66 21
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
rect 75 79 77 81
rect 83 79 85 81
rect 91 79 93 81
rect 99 79 101 81
rect 107 79 109 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
rect 75 -1 77 1
rect 83 -1 85 1
rect 91 -1 93 1
rect 99 -1 101 1
rect 107 -1 109 1
<< pdifct0 >>
rect 4 64 6 66
rect 14 58 16 60
rect 24 64 26 66
rect 44 64 46 66
rect 64 56 66 58
rect 84 56 86 58
rect 96 51 98 53
rect 96 44 98 46
rect 106 60 108 62
<< pdifct1 >>
rect 14 51 16 53
rect 34 59 36 61
rect 34 51 36 53
rect 54 51 56 53
rect 54 44 56 46
rect 74 51 76 53
rect 74 44 76 46
<< alu0 >>
rect 3 66 7 68
rect 3 64 4 66
rect 6 64 7 66
rect 3 62 7 64
rect 23 66 27 68
rect 23 64 24 66
rect 26 64 27 66
rect 23 62 27 64
rect 43 66 47 68
rect 43 64 44 66
rect 46 64 47 66
rect 13 60 17 62
rect 13 58 14 60
rect 16 58 17 60
rect 13 55 17 58
rect 15 54 17 55
rect 43 62 47 64
rect 63 58 67 68
rect 63 56 64 58
rect 66 56 67 58
rect 63 54 67 56
rect 83 58 87 68
rect 104 62 110 68
rect 104 60 106 62
rect 108 60 110 62
rect 104 59 110 60
rect 83 56 84 58
rect 86 56 87 58
rect 83 54 87 56
rect 95 53 99 55
rect 95 51 96 53
rect 98 51 99 53
rect 95 46 99 51
rect 82 44 96 46
rect 98 44 99 46
rect 82 42 99 44
rect 10 37 14 39
rect 10 35 11 37
rect 13 35 14 37
rect 10 30 14 35
rect 35 37 41 38
rect 35 35 37 37
rect 39 35 41 37
rect 35 30 41 35
rect 82 37 86 42
rect 82 35 83 37
rect 85 35 86 37
rect 82 30 86 35
rect 10 28 100 30
rect 10 26 96 28
rect 98 26 100 28
rect 94 25 100 26
rect 105 23 109 25
rect 81 21 87 22
rect 81 19 83 21
rect 85 19 87 21
rect 5 14 11 15
rect 5 12 7 14
rect 9 12 11 14
rect 42 14 48 15
rect 42 12 44 14
rect 46 12 48 14
rect 81 14 87 19
rect 81 12 83 14
rect 85 12 87 14
rect 105 21 106 23
rect 108 21 109 23
rect 105 12 109 21
<< labels >>
rlabel alu0 12 32 12 32 6 an
rlabel alu0 38 32 38 32 6 an
rlabel ndifct0 97 27 97 27 6 an
rlabel alu0 97 48 97 48 6 an
rlabel polyct0 84 36 84 36 6 an
rlabel alu1 12 20 12 20 6 z
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 52 12 52 6 z
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 20 28 20 6 z
rlabel alu1 36 20 36 20 6 z
rlabel alu1 28 40 28 40 6 b
rlabel alu1 36 44 36 44 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 20 52 20 52 6 z
rlabel alu1 36 56 36 56 6 z
rlabel alu1 56 6 56 6 6 vss
rlabel alu1 44 20 44 20 6 z
rlabel alu1 52 20 52 20 6 z
rlabel alu1 60 20 60 20 6 z
rlabel alu1 44 44 44 44 6 b
rlabel alu1 52 36 52 36 6 b
rlabel alu1 60 36 60 36 6 b
rlabel alu1 60 44 60 44 6 z
rlabel alu1 52 52 52 52 6 z
rlabel alu1 44 52 44 52 6 z
rlabel alu1 56 74 56 74 6 vdd
rlabel alu1 68 20 68 20 6 z
rlabel alu1 68 36 68 36 6 b
rlabel alu1 68 44 68 44 6 z
rlabel alu1 76 52 76 52 6 z
rlabel polyct1 100 36 100 36 6 a
rlabel alu1 108 48 108 48 6 a
<< end >>
