magic
tech scmos
timestamp 1199203665
<< ab >>
rect 0 0 72 80
<< nwell >>
rect -5 36 77 88
<< pwell >>
rect -5 -8 77 36
<< poly >>
rect 20 69 22 74
rect 30 69 32 74
rect 40 69 42 74
rect 50 69 52 74
rect 2 60 8 62
rect 2 58 4 60
rect 6 58 8 60
rect 2 56 11 58
rect 9 53 11 56
rect 61 55 63 60
rect 9 39 11 42
rect 20 39 22 42
rect 30 39 32 42
rect 9 37 22 39
rect 26 37 32 39
rect 9 28 11 37
rect 26 35 28 37
rect 30 35 32 37
rect 26 33 32 35
rect 40 39 42 42
rect 50 39 52 42
rect 61 39 63 44
rect 40 37 46 39
rect 40 35 42 37
rect 44 35 46 37
rect 40 33 46 35
rect 50 37 70 39
rect 19 31 28 33
rect 19 28 21 31
rect 40 30 42 33
rect 50 30 52 37
rect 61 35 66 37
rect 68 35 70 37
rect 61 33 70 35
rect 61 30 63 33
rect 9 8 11 22
rect 29 23 31 27
rect 19 12 21 16
rect 61 19 63 24
rect 40 13 42 18
rect 50 13 52 18
rect 29 8 31 11
rect 9 6 31 8
<< ndif >>
rect 33 28 40 30
rect 2 26 9 28
rect 2 24 4 26
rect 6 24 9 26
rect 2 22 9 24
rect 11 26 19 28
rect 11 24 14 26
rect 16 24 19 26
rect 11 22 19 24
rect 13 16 19 22
rect 21 23 26 28
rect 33 26 35 28
rect 37 26 40 28
rect 33 23 40 26
rect 21 20 29 23
rect 21 18 24 20
rect 26 18 29 20
rect 21 16 29 18
rect 24 11 29 16
rect 31 18 40 23
rect 42 22 50 30
rect 42 20 45 22
rect 47 20 50 22
rect 42 18 50 20
rect 52 24 61 30
rect 63 28 70 30
rect 63 26 66 28
rect 68 26 70 28
rect 63 24 70 26
rect 52 22 59 24
rect 52 20 55 22
rect 57 20 59 22
rect 52 18 59 20
rect 31 11 36 18
<< pdif >>
rect 13 65 20 69
rect 13 63 15 65
rect 17 63 20 65
rect 13 53 20 63
rect 4 48 9 53
rect 2 46 9 48
rect 2 44 4 46
rect 6 44 9 46
rect 2 42 9 44
rect 11 42 20 53
rect 22 62 30 69
rect 22 60 25 62
rect 27 60 30 62
rect 22 42 30 60
rect 32 53 40 69
rect 32 51 35 53
rect 37 51 40 53
rect 32 46 40 51
rect 32 44 35 46
rect 37 44 40 46
rect 32 42 40 44
rect 42 62 50 69
rect 42 60 45 62
rect 47 60 50 62
rect 42 42 50 60
rect 52 61 59 69
rect 52 59 55 61
rect 57 59 59 61
rect 52 55 59 59
rect 52 44 61 55
rect 63 53 70 55
rect 63 51 66 53
rect 68 51 70 53
rect 63 49 70 51
rect 63 44 68 49
rect 52 42 59 44
<< alu1 >>
rect -2 81 74 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 74 81
rect -2 68 74 79
rect 2 60 7 63
rect 2 58 4 60
rect 6 58 7 60
rect 2 54 14 58
rect 10 49 14 54
rect 26 53 38 55
rect 26 51 35 53
rect 37 51 38 53
rect 26 49 38 51
rect 34 46 38 49
rect 34 44 35 46
rect 37 44 38 46
rect 34 28 38 44
rect 57 42 70 46
rect 65 37 70 42
rect 65 35 66 37
rect 68 35 70 37
rect 65 33 70 35
rect 34 26 35 28
rect 37 26 38 28
rect 34 24 38 26
rect -2 1 74 12
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 74 1
rect -2 -2 74 -1
<< ptie >>
rect 0 1 72 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 43 1
rect 45 -1 51 1
rect 53 -1 59 1
rect 61 -1 67 1
rect 69 -1 72 1
rect 0 -3 72 -1
<< ntie >>
rect 0 81 72 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 43 81
rect 45 79 51 81
rect 53 79 59 81
rect 61 79 67 81
rect 69 79 72 81
rect 0 77 72 79
<< nmos >>
rect 9 22 11 28
rect 19 16 21 28
rect 29 11 31 23
rect 40 18 42 30
rect 50 18 52 30
rect 61 24 63 30
<< pmos >>
rect 9 42 11 53
rect 20 42 22 69
rect 30 42 32 69
rect 40 42 42 69
rect 50 42 52 69
rect 61 44 63 55
<< polyct0 >>
rect 28 35 30 37
rect 42 35 44 37
<< polyct1 >>
rect 4 58 6 60
rect 66 35 68 37
<< ndifct0 >>
rect 4 24 6 26
rect 14 24 16 26
rect 24 18 26 20
rect 45 20 47 22
rect 66 26 68 28
rect 55 20 57 22
<< ndifct1 >>
rect 35 26 37 28
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
rect 43 79 45 81
rect 51 79 53 81
rect 59 79 61 81
rect 67 79 69 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
rect 43 -1 45 1
rect 51 -1 53 1
rect 59 -1 61 1
rect 67 -1 69 1
<< pdifct0 >>
rect 15 63 17 65
rect 4 44 6 46
rect 25 60 27 62
rect 45 60 47 62
rect 55 59 57 61
rect 66 51 68 53
<< pdifct1 >>
rect 35 51 37 53
rect 35 44 37 46
<< alu0 >>
rect 13 65 19 68
rect 13 63 15 65
rect 17 63 19 65
rect 13 62 19 63
rect 23 62 49 63
rect 23 60 25 62
rect 27 60 45 62
rect 47 60 49 62
rect 23 59 49 60
rect 53 61 59 68
rect 53 59 55 61
rect 57 59 59 61
rect 53 58 59 59
rect 3 46 7 48
rect 3 44 4 46
rect 6 44 7 46
rect 3 37 7 44
rect 27 37 31 39
rect 3 35 28 37
rect 30 35 31 37
rect 3 33 31 35
rect 3 26 7 33
rect 50 53 70 54
rect 50 51 66 53
rect 68 51 70 53
rect 50 50 70 51
rect 50 39 54 50
rect 41 37 54 39
rect 41 35 42 37
rect 44 35 54 37
rect 41 33 54 35
rect 3 24 4 26
rect 6 24 7 26
rect 3 22 7 24
rect 13 26 17 28
rect 13 24 14 26
rect 16 24 17 26
rect 50 30 54 33
rect 50 28 70 30
rect 50 26 66 28
rect 68 26 70 28
rect 64 25 70 26
rect 13 12 17 24
rect 43 22 49 23
rect 43 21 45 22
rect 22 20 45 21
rect 47 20 49 22
rect 22 18 24 20
rect 26 18 49 20
rect 22 17 49 18
rect 53 22 59 23
rect 53 20 55 22
rect 57 20 59 22
rect 53 12 59 20
<< labels >>
rlabel alu0 17 35 17 35 6 bn
rlabel alu0 35 19 35 19 6 n2
rlabel alu0 36 61 36 61 6 n1
rlabel alu0 47 36 47 36 6 an
rlabel ndifct0 67 27 67 27 6 an
rlabel alu0 60 52 60 52 6 an
rlabel alu1 12 52 12 52 6 b
rlabel alu1 4 60 4 60 6 b
rlabel alu1 28 52 28 52 6 z
rlabel alu1 36 6 36 6 6 vss
rlabel alu1 36 40 36 40 6 z
rlabel alu1 36 74 36 74 6 vdd
rlabel alu1 68 36 68 36 6 a
rlabel alu1 60 44 60 44 6 a
<< end >>
