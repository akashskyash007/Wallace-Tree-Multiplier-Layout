magic
tech scmos
timestamp 1199203705
<< ab >>
rect 0 0 128 72
<< nwell >>
rect -5 32 133 77
<< pwell >>
rect -5 -5 133 32
<< poly >>
rect 9 66 11 70
rect 19 66 21 70
rect 29 66 31 70
rect 39 66 41 70
rect 49 66 51 70
rect 69 66 71 70
rect 79 66 81 70
rect 89 66 91 70
rect 39 49 41 52
rect 49 49 51 52
rect 39 47 51 49
rect 45 45 47 47
rect 49 45 51 47
rect 45 43 51 45
rect 100 59 102 63
rect 110 59 112 63
rect 100 42 102 45
rect 110 42 112 45
rect 100 40 126 42
rect 9 35 11 38
rect 19 35 21 38
rect 29 35 31 38
rect 69 35 71 38
rect 79 35 81 38
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 29 33 65 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 10 20 12 29
rect 19 25 21 29
rect 37 25 39 33
rect 59 31 61 33
rect 63 31 65 33
rect 59 29 65 31
rect 69 33 75 35
rect 69 31 71 33
rect 73 31 75 33
rect 69 29 75 31
rect 79 33 85 35
rect 79 31 81 33
rect 83 31 85 33
rect 89 34 91 38
rect 89 32 103 34
rect 79 29 85 31
rect 97 30 99 32
rect 101 30 103 32
rect 49 27 55 29
rect 49 25 51 27
rect 53 25 55 27
rect 17 23 21 25
rect 17 20 19 23
rect 27 20 29 25
rect 49 23 55 25
rect 49 20 51 23
rect 72 20 74 29
rect 79 20 81 29
rect 97 28 103 30
rect 99 25 101 28
rect 110 26 112 40
rect 120 38 122 40
rect 124 38 126 40
rect 120 36 126 38
rect 89 20 91 25
rect 37 8 39 12
rect 10 2 12 7
rect 17 2 19 7
rect 27 4 29 7
rect 49 4 51 9
rect 27 2 51 4
rect 99 8 101 12
rect 72 2 74 7
rect 79 2 81 7
rect 89 4 91 7
rect 110 4 112 15
rect 89 2 112 4
<< ndif >>
rect 32 20 37 25
rect 2 7 10 20
rect 12 7 17 20
rect 19 17 27 20
rect 19 15 22 17
rect 24 15 27 17
rect 19 7 27 15
rect 29 18 37 20
rect 29 16 32 18
rect 34 16 37 18
rect 29 12 37 16
rect 39 20 47 25
rect 105 25 110 26
rect 94 20 99 25
rect 39 12 49 20
rect 29 7 34 12
rect 41 10 49 12
rect 41 8 43 10
rect 45 9 49 10
rect 51 18 58 20
rect 51 16 54 18
rect 56 16 58 18
rect 51 14 58 16
rect 51 9 56 14
rect 45 8 47 9
rect 2 5 4 7
rect 6 5 8 7
rect 2 3 8 5
rect 41 6 47 8
rect 64 7 72 20
rect 74 7 79 20
rect 81 17 89 20
rect 81 15 84 17
rect 86 15 89 17
rect 81 7 89 15
rect 91 18 99 20
rect 91 16 94 18
rect 96 16 99 18
rect 91 12 99 16
rect 101 16 110 25
rect 101 14 104 16
rect 106 15 110 16
rect 112 24 119 26
rect 112 22 115 24
rect 117 22 119 24
rect 112 20 119 22
rect 112 15 117 20
rect 106 14 108 15
rect 101 12 108 14
rect 91 7 96 12
rect 64 5 66 7
rect 68 5 70 7
rect 64 3 70 5
<< pdif >>
rect 4 59 9 66
rect 2 57 9 59
rect 2 55 4 57
rect 6 55 9 57
rect 2 53 9 55
rect 4 38 9 53
rect 11 49 19 66
rect 11 47 14 49
rect 16 47 19 49
rect 11 38 19 47
rect 21 49 29 66
rect 21 47 24 49
rect 26 47 29 49
rect 21 42 29 47
rect 21 40 24 42
rect 26 40 29 42
rect 21 38 29 40
rect 31 64 39 66
rect 31 62 34 64
rect 36 62 39 64
rect 31 52 39 62
rect 41 57 49 66
rect 41 55 44 57
rect 46 55 49 57
rect 41 52 49 55
rect 51 64 58 66
rect 51 62 54 64
rect 56 62 58 64
rect 51 57 58 62
rect 64 59 69 66
rect 51 55 54 57
rect 56 55 58 57
rect 51 52 58 55
rect 62 57 69 59
rect 62 55 64 57
rect 66 55 69 57
rect 62 53 69 55
rect 31 38 37 52
rect 64 38 69 53
rect 71 49 79 66
rect 71 47 74 49
rect 76 47 79 49
rect 71 38 79 47
rect 81 49 89 66
rect 81 47 84 49
rect 86 47 89 49
rect 81 42 89 47
rect 81 40 84 42
rect 86 40 89 42
rect 81 38 89 40
rect 91 64 98 66
rect 91 62 94 64
rect 96 62 98 64
rect 91 59 98 62
rect 91 45 100 59
rect 102 49 110 59
rect 102 47 105 49
rect 107 47 110 49
rect 102 45 110 47
rect 112 57 120 59
rect 112 55 115 57
rect 117 55 120 57
rect 112 45 120 55
rect 91 38 98 45
<< alu1 >>
rect -2 67 130 72
rect -2 65 121 67
rect 123 65 130 67
rect -2 64 130 65
rect 2 49 18 50
rect 2 47 14 49
rect 16 47 18 49
rect 2 46 18 47
rect 2 18 6 46
rect 41 47 54 50
rect 41 45 47 47
rect 49 45 54 47
rect 41 44 54 45
rect 2 17 26 18
rect 2 15 22 17
rect 24 15 26 17
rect 2 14 26 15
rect 50 27 54 44
rect 50 25 51 27
rect 53 25 54 27
rect 50 23 54 25
rect 113 46 126 51
rect 122 42 126 46
rect 98 32 111 35
rect 98 30 99 32
rect 101 30 111 32
rect 98 29 111 30
rect 105 22 111 29
rect 121 40 126 42
rect 121 38 122 40
rect 124 38 126 40
rect 121 36 126 38
rect 122 29 126 36
rect -2 7 130 8
rect -2 5 4 7
rect 6 5 66 7
rect 68 5 121 7
rect 123 5 130 7
rect -2 0 130 5
<< ptie >>
rect 119 7 125 9
rect 119 5 121 7
rect 123 5 125 7
rect 119 3 125 5
<< ntie >>
rect 119 67 125 69
rect 119 65 121 67
rect 123 65 125 67
rect 119 63 125 65
<< nmos >>
rect 10 7 12 20
rect 17 7 19 20
rect 27 7 29 20
rect 37 12 39 25
rect 49 9 51 20
rect 72 7 74 20
rect 79 7 81 20
rect 89 7 91 20
rect 99 12 101 25
rect 110 15 112 26
<< pmos >>
rect 9 38 11 66
rect 19 38 21 66
rect 29 38 31 66
rect 39 52 41 66
rect 49 52 51 66
rect 69 38 71 66
rect 79 38 81 66
rect 89 38 91 66
rect 100 45 102 59
rect 110 45 112 59
<< polyct0 >>
rect 11 31 13 33
rect 21 31 23 33
rect 61 31 63 33
rect 71 31 73 33
rect 81 31 83 33
<< polyct1 >>
rect 47 45 49 47
rect 99 30 101 32
rect 51 25 53 27
rect 122 38 124 40
<< ndifct0 >>
rect 32 16 34 18
rect 43 8 45 10
rect 54 16 56 18
rect 84 15 86 17
rect 94 16 96 18
rect 104 14 106 16
rect 115 22 117 24
<< ndifct1 >>
rect 22 15 24 17
rect 4 5 6 7
rect 66 5 68 7
<< ntiect1 >>
rect 121 65 123 67
<< ptiect1 >>
rect 121 5 123 7
<< pdifct0 >>
rect 4 55 6 57
rect 24 47 26 49
rect 24 40 26 42
rect 34 62 36 64
rect 44 55 46 57
rect 54 62 56 64
rect 54 55 56 57
rect 64 55 66 57
rect 74 47 76 49
rect 84 47 86 49
rect 84 40 86 42
rect 94 62 96 64
rect 105 47 107 49
rect 115 55 117 57
<< pdifct1 >>
rect 14 47 16 49
<< alu0 >>
rect 32 62 34 64
rect 36 62 38 64
rect 32 61 38 62
rect 52 62 54 64
rect 56 62 58 64
rect 2 57 48 58
rect 2 55 4 57
rect 6 55 44 57
rect 46 55 48 57
rect 2 54 48 55
rect 52 57 58 62
rect 92 62 94 64
rect 96 62 98 64
rect 92 61 98 62
rect 52 55 54 57
rect 56 55 58 57
rect 52 54 58 55
rect 62 57 94 58
rect 62 55 64 57
rect 66 55 94 57
rect 62 54 94 55
rect 113 57 119 64
rect 113 55 115 57
rect 117 55 119 57
rect 113 54 119 55
rect 22 49 28 50
rect 22 47 24 49
rect 26 47 28 49
rect 22 43 28 47
rect 10 42 28 43
rect 10 40 24 42
rect 26 40 28 42
rect 10 39 28 40
rect 10 33 14 39
rect 32 34 36 54
rect 90 51 94 54
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 19 33 45 34
rect 19 31 21 33
rect 23 31 45 33
rect 19 30 45 31
rect 10 22 35 26
rect 31 18 35 22
rect 31 16 32 18
rect 34 16 35 18
rect 31 14 35 16
rect 41 19 45 30
rect 62 49 78 50
rect 62 47 74 49
rect 76 47 78 49
rect 62 46 78 47
rect 83 49 87 51
rect 83 47 84 49
rect 86 47 87 49
rect 62 34 66 46
rect 83 42 87 47
rect 59 33 66 34
rect 59 31 61 33
rect 63 31 66 33
rect 59 30 66 31
rect 41 18 58 19
rect 41 16 54 18
rect 56 16 58 18
rect 41 15 58 16
rect 62 18 66 30
rect 70 40 84 42
rect 86 40 87 42
rect 70 38 87 40
rect 90 49 108 51
rect 90 47 105 49
rect 107 47 108 49
rect 70 33 74 38
rect 90 34 94 47
rect 104 42 108 47
rect 104 38 118 42
rect 70 31 71 33
rect 73 31 74 33
rect 70 26 74 31
rect 79 33 94 34
rect 79 31 81 33
rect 83 31 94 33
rect 79 30 94 31
rect 70 22 97 26
rect 114 24 118 38
rect 114 22 115 24
rect 117 22 118 24
rect 93 18 97 22
rect 114 20 118 22
rect 62 17 88 18
rect 62 15 84 17
rect 86 15 88 17
rect 62 14 88 15
rect 93 16 94 18
rect 96 16 97 18
rect 93 14 97 16
rect 103 16 107 18
rect 103 14 104 16
rect 106 14 107 16
rect 41 10 47 11
rect 41 8 43 10
rect 45 8 47 10
rect 103 8 107 14
<< labels >>
rlabel alu0 49 17 49 17 6 cn
rlabel alu0 25 56 25 56 6 cn
rlabel alu0 34 44 34 44 6 cn
rlabel alu0 85 44 85 44 6 an
rlabel polyct0 72 32 72 32 6 an
rlabel alu0 95 20 95 20 6 an
rlabel alu0 86 32 86 32 6 bn
rlabel alu0 106 44 106 44 6 bn
rlabel alu0 116 31 116 31 6 bn
rlabel alu0 78 56 78 56 6 bn
rlabel alu1 20 16 20 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 48 12 48 6 z
rlabel alu1 52 36 52 36 6 c
rlabel alu1 44 48 44 48 6 c
rlabel alu1 64 4 64 4 6 vss
rlabel alu1 64 68 64 68 6 vdd
rlabel alu1 100 32 100 32 6 a
rlabel alu1 108 28 108 28 6 a
rlabel alu1 124 40 124 40 6 b
rlabel alu1 116 48 116 48 6 b
<< end >>
