magic
tech scmos
timestamp 1199201717
<< ab >>
rect 0 0 56 72
<< nwell >>
rect -5 32 61 77
<< pwell >>
rect -5 -5 61 32
<< poly >>
rect 9 66 11 70
rect 19 63 21 68
rect 29 63 31 68
rect 41 63 43 68
rect 9 35 11 38
rect 19 35 21 46
rect 29 43 31 46
rect 29 41 35 43
rect 29 39 31 41
rect 33 39 35 41
rect 29 37 35 39
rect 9 33 15 35
rect 9 31 11 33
rect 13 31 15 33
rect 9 29 15 31
rect 19 33 25 35
rect 19 31 21 33
rect 23 31 25 33
rect 19 29 25 31
rect 9 25 11 29
rect 22 25 24 29
rect 29 25 31 37
rect 41 35 43 46
rect 41 33 47 35
rect 41 31 43 33
rect 45 31 47 33
rect 36 29 47 31
rect 36 25 38 29
rect 9 6 11 11
rect 22 3 24 8
rect 29 3 31 8
rect 36 3 38 8
<< ndif >>
rect 4 19 9 25
rect 2 17 9 19
rect 2 15 4 17
rect 6 15 9 17
rect 2 13 9 15
rect 4 11 9 13
rect 11 11 22 25
rect 13 8 22 11
rect 24 8 29 25
rect 31 8 36 25
rect 38 18 43 25
rect 38 16 45 18
rect 38 14 41 16
rect 43 14 45 16
rect 38 12 45 14
rect 38 8 43 12
rect 13 7 20 8
rect 13 5 16 7
rect 18 5 20 7
rect 13 3 20 5
<< pdif >>
rect 4 51 9 66
rect 2 49 9 51
rect 2 47 4 49
rect 6 47 9 49
rect 2 42 9 47
rect 2 40 4 42
rect 6 40 9 42
rect 2 38 9 40
rect 11 63 17 66
rect 33 67 39 69
rect 33 65 35 67
rect 37 65 39 67
rect 33 63 39 65
rect 11 61 19 63
rect 11 59 14 61
rect 16 59 19 61
rect 11 46 19 59
rect 21 57 29 63
rect 21 55 24 57
rect 26 55 29 57
rect 21 50 29 55
rect 21 48 24 50
rect 26 48 29 50
rect 21 46 29 48
rect 31 46 41 63
rect 43 60 48 63
rect 43 58 50 60
rect 43 56 46 58
rect 48 56 50 58
rect 43 54 50 56
rect 43 46 48 54
rect 11 38 17 46
<< alu1 >>
rect -2 67 58 72
rect -2 65 35 67
rect 37 65 58 67
rect -2 64 58 65
rect 2 49 7 51
rect 2 47 4 49
rect 6 47 7 49
rect 2 42 7 47
rect 2 40 4 42
rect 6 40 7 42
rect 2 38 7 40
rect 2 18 6 38
rect 18 34 22 43
rect 42 42 46 51
rect 29 41 46 42
rect 29 39 31 41
rect 33 39 46 41
rect 29 38 46 39
rect 18 33 31 34
rect 18 31 21 33
rect 23 31 31 33
rect 18 30 31 31
rect 41 33 47 34
rect 41 31 43 33
rect 45 31 47 33
rect 41 26 47 31
rect 33 22 47 26
rect 2 17 15 18
rect 2 15 4 17
rect 6 15 15 17
rect 2 13 15 15
rect -2 7 58 8
rect -2 5 16 7
rect 18 5 58 7
rect -2 0 58 5
<< nmos >>
rect 9 11 11 25
rect 22 8 24 25
rect 29 8 31 25
rect 36 8 38 25
<< pmos >>
rect 9 38 11 66
rect 19 46 21 63
rect 29 46 31 63
rect 41 46 43 63
<< polyct0 >>
rect 11 31 13 33
<< polyct1 >>
rect 31 39 33 41
rect 21 31 23 33
rect 43 31 45 33
<< ndifct0 >>
rect 41 14 43 16
<< ndifct1 >>
rect 4 15 6 17
rect 16 5 18 7
<< pdifct0 >>
rect 14 59 16 61
rect 24 55 26 57
rect 24 48 26 50
rect 46 56 48 58
<< pdifct1 >>
rect 4 47 6 49
rect 4 40 6 42
rect 35 65 37 67
<< alu0 >>
rect 13 61 17 64
rect 13 59 14 61
rect 16 59 17 61
rect 13 57 17 59
rect 23 58 50 59
rect 23 57 46 58
rect 23 55 24 57
rect 26 56 46 57
rect 48 56 50 58
rect 26 55 50 56
rect 23 51 28 55
rect 10 50 28 51
rect 10 48 24 50
rect 26 48 28 50
rect 10 47 28 48
rect 10 33 14 47
rect 10 31 11 33
rect 13 31 14 33
rect 10 26 14 31
rect 10 22 26 26
rect 22 17 26 22
rect 22 16 45 17
rect 22 14 41 16
rect 43 14 45 16
rect 22 13 45 14
<< labels >>
rlabel alu0 12 36 12 36 6 zn
rlabel alu0 25 53 25 53 6 zn
rlabel alu0 19 49 19 49 6 zn
rlabel alu0 33 15 33 15 6 zn
rlabel alu0 36 57 36 57 6 zn
rlabel alu1 4 32 4 32 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 40 20 40 6 a
rlabel alu1 28 4 28 4 6 vss
rlabel alu1 28 32 28 32 6 a
rlabel alu1 36 24 36 24 6 c
rlabel alu1 36 40 36 40 6 b
rlabel alu1 28 68 28 68 6 vdd
rlabel alu1 44 28 44 28 6 c
rlabel alu1 44 48 44 48 6 b
<< end >>
