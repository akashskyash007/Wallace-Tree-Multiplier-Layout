magic
tech scmos
timestamp 1199202847
<< ab >>
rect 0 0 80 72
<< nwell >>
rect -5 32 85 77
<< pwell >>
rect -5 -5 85 32
<< poly >>
rect 9 65 11 70
rect 19 65 21 70
rect 32 65 34 70
rect 42 65 44 70
rect 64 49 70 51
rect 64 47 66 49
rect 68 47 70 49
rect 64 45 70 47
rect 54 41 60 43
rect 9 31 11 40
rect 19 37 21 40
rect 32 37 34 40
rect 19 35 25 37
rect 19 33 21 35
rect 23 33 25 35
rect 32 35 38 37
rect 32 33 34 35
rect 36 33 38 35
rect 19 31 25 33
rect 29 31 38 33
rect 42 35 44 40
rect 54 39 56 41
rect 58 39 60 41
rect 54 37 60 39
rect 42 33 49 35
rect 42 31 45 33
rect 47 31 49 33
rect 9 29 15 31
rect 9 27 11 29
rect 13 27 15 29
rect 9 25 17 27
rect 15 22 17 25
rect 22 22 24 31
rect 29 22 31 31
rect 42 29 49 31
rect 42 27 48 29
rect 54 28 56 37
rect 64 33 66 45
rect 36 25 48 27
rect 36 22 38 25
rect 46 22 48 25
rect 53 25 56 28
rect 60 31 66 33
rect 53 22 55 25
rect 60 22 62 31
rect 72 29 78 31
rect 72 27 74 29
rect 76 27 78 29
rect 67 25 78 27
rect 67 22 69 25
rect 15 2 17 7
rect 22 2 24 7
rect 29 2 31 7
rect 36 2 38 7
rect 46 2 48 7
rect 53 2 55 7
rect 60 2 62 7
rect 67 2 69 7
<< ndif >>
rect 6 7 15 22
rect 17 7 22 22
rect 24 7 29 22
rect 31 7 36 22
rect 38 17 46 22
rect 38 15 41 17
rect 43 15 46 17
rect 38 7 46 15
rect 48 7 53 22
rect 55 7 60 22
rect 62 7 67 22
rect 69 11 77 22
rect 69 9 72 11
rect 74 9 77 11
rect 69 7 77 9
rect 6 5 9 7
rect 11 5 13 7
rect 6 3 13 5
<< pdif >>
rect 24 65 30 67
rect 2 63 9 65
rect 2 61 4 63
rect 6 61 9 63
rect 2 56 9 61
rect 2 54 4 56
rect 6 54 9 56
rect 2 40 9 54
rect 11 57 19 65
rect 11 55 14 57
rect 16 55 19 57
rect 11 49 19 55
rect 11 47 14 49
rect 16 47 19 49
rect 11 40 19 47
rect 21 64 32 65
rect 21 62 26 64
rect 28 62 32 64
rect 21 40 32 62
rect 34 57 42 65
rect 34 55 37 57
rect 39 55 42 57
rect 34 40 42 55
rect 44 63 52 65
rect 44 61 47 63
rect 49 61 52 63
rect 44 56 52 61
rect 44 54 47 56
rect 49 54 52 56
rect 44 40 52 54
<< alu1 >>
rect -2 67 82 72
rect -2 65 58 67
rect 60 65 73 67
rect 75 65 82 67
rect -2 64 82 65
rect 12 57 41 58
rect 12 55 14 57
rect 16 55 37 57
rect 39 55 41 57
rect 12 54 41 55
rect 12 50 18 54
rect 58 50 62 59
rect 2 49 18 50
rect 2 47 14 49
rect 16 47 18 49
rect 2 46 18 47
rect 24 49 71 50
rect 24 47 66 49
rect 68 47 71 49
rect 24 46 71 47
rect 2 18 6 46
rect 24 42 28 46
rect 17 38 28 42
rect 33 41 60 42
rect 33 39 56 41
rect 58 39 60 41
rect 33 38 60 39
rect 64 38 71 42
rect 20 35 24 38
rect 20 33 21 35
rect 23 33 24 35
rect 20 31 24 33
rect 33 35 39 38
rect 33 33 34 35
rect 36 33 39 35
rect 64 34 68 38
rect 10 29 14 31
rect 33 30 39 33
rect 43 33 68 34
rect 43 31 45 33
rect 47 31 68 33
rect 43 30 68 31
rect 10 27 11 29
rect 13 27 14 29
rect 10 26 14 27
rect 72 29 78 31
rect 72 27 74 29
rect 76 27 78 29
rect 72 26 78 27
rect 10 22 78 26
rect 58 21 78 22
rect 2 17 47 18
rect 2 15 41 17
rect 43 15 47 17
rect 2 14 47 15
rect 58 13 62 21
rect -2 7 82 8
rect -2 5 9 7
rect 11 5 82 7
rect -2 0 82 5
<< ntie >>
rect 56 67 77 69
rect 56 65 58 67
rect 60 65 73 67
rect 75 65 77 67
rect 56 63 77 65
<< nmos >>
rect 15 7 17 22
rect 22 7 24 22
rect 29 7 31 22
rect 36 7 38 22
rect 46 7 48 22
rect 53 7 55 22
rect 60 7 62 22
rect 67 7 69 22
<< pmos >>
rect 9 40 11 65
rect 19 40 21 65
rect 32 40 34 65
rect 42 40 44 65
<< polyct1 >>
rect 66 47 68 49
rect 21 33 23 35
rect 34 33 36 35
rect 56 39 58 41
rect 45 31 47 33
rect 11 27 13 29
rect 74 27 76 29
<< ndifct0 >>
rect 72 9 74 11
<< ndifct1 >>
rect 41 15 43 17
rect 9 5 11 7
<< ntiect1 >>
rect 58 65 60 67
rect 73 65 75 67
<< pdifct0 >>
rect 4 61 6 63
rect 4 54 6 56
rect 26 62 28 64
rect 47 61 49 63
rect 47 54 49 56
<< pdifct1 >>
rect 14 55 16 57
rect 14 47 16 49
rect 37 55 39 57
<< alu0 >>
rect 2 63 8 64
rect 2 61 4 63
rect 6 61 8 63
rect 24 62 26 64
rect 28 62 30 64
rect 24 61 30 62
rect 45 63 51 64
rect 45 61 47 63
rect 49 61 51 63
rect 2 56 8 61
rect 2 54 4 56
rect 6 54 8 56
rect 2 53 8 54
rect 45 56 51 61
rect 45 54 47 56
rect 49 54 51 56
rect 45 53 51 54
rect 71 11 75 13
rect 71 9 72 11
rect 74 9 75 11
rect 71 8 75 9
<< labels >>
rlabel alu1 4 32 4 32 6 z
rlabel alu1 20 16 20 16 6 z
rlabel alu1 28 16 28 16 6 z
rlabel alu1 12 16 12 16 6 z
rlabel alu1 20 24 20 24 6 a
rlabel alu1 28 24 28 24 6 a
rlabel alu1 20 40 20 40 6 b
rlabel alu1 12 48 12 48 6 z
rlabel alu1 28 48 28 48 6 b
rlabel alu1 20 56 20 56 6 z
rlabel alu1 28 56 28 56 6 z
rlabel alu1 40 4 40 4 6 vss
rlabel alu1 36 16 36 16 6 z
rlabel alu1 44 16 44 16 6 z
rlabel alu1 36 24 36 24 6 a
rlabel alu1 44 24 44 24 6 a
rlabel alu1 44 40 44 40 6 c
rlabel alu1 36 36 36 36 6 c
rlabel alu1 36 48 36 48 6 b
rlabel alu1 44 48 44 48 6 b
rlabel alu1 36 56 36 56 6 z
rlabel alu1 40 68 40 68 6 vdd
rlabel alu1 52 24 52 24 6 a
rlabel alu1 60 20 60 20 6 a
rlabel alu1 60 32 60 32 6 d
rlabel alu1 52 32 52 32 6 d
rlabel alu1 52 40 52 40 6 c
rlabel alu1 52 48 52 48 6 b
rlabel alu1 60 52 60 52 6 b
rlabel alu1 68 24 68 24 6 a
rlabel alu1 76 24 76 24 6 a
rlabel alu1 68 40 68 40 6 d
rlabel alu1 68 48 68 48 6 b
<< end >>
