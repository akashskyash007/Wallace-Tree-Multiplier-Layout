magic
tech scmos
timestamp 1199201847
<< ab >>
rect 0 0 40 80
<< nwell >>
rect -5 36 45 88
<< pwell >>
rect -5 -8 45 36
<< poly >>
rect 9 69 11 74
rect 19 69 21 74
rect 29 69 31 74
rect 9 39 11 42
rect 19 39 21 42
rect 9 37 15 39
rect 9 35 11 37
rect 13 35 15 37
rect 9 33 15 35
rect 19 37 25 39
rect 19 35 21 37
rect 23 35 25 37
rect 19 33 25 35
rect 10 22 12 33
rect 20 22 22 33
rect 29 31 31 42
rect 29 29 35 31
rect 29 28 31 29
rect 27 27 31 28
rect 33 27 35 29
rect 27 25 35 27
rect 27 22 29 25
rect 10 10 12 15
rect 20 6 22 10
rect 27 6 29 10
<< ndif >>
rect 2 15 10 22
rect 12 20 20 22
rect 12 18 15 20
rect 17 18 20 20
rect 12 15 20 18
rect 2 11 8 15
rect 2 9 4 11
rect 6 9 8 11
rect 15 10 20 15
rect 22 10 27 22
rect 29 11 38 22
rect 29 10 33 11
rect 2 7 8 9
rect 31 9 33 10
rect 35 9 38 11
rect 31 7 38 9
<< pdif >>
rect 4 63 9 69
rect 2 61 9 63
rect 2 59 4 61
rect 6 59 9 61
rect 2 54 9 59
rect 2 52 4 54
rect 6 52 9 54
rect 2 50 9 52
rect 4 42 9 50
rect 11 61 19 69
rect 11 59 14 61
rect 16 59 19 61
rect 11 54 19 59
rect 11 52 14 54
rect 16 52 19 54
rect 11 42 19 52
rect 21 67 29 69
rect 21 65 24 67
rect 26 65 29 67
rect 21 60 29 65
rect 21 58 24 60
rect 26 58 29 60
rect 21 42 29 58
rect 31 63 36 69
rect 31 61 38 63
rect 31 59 34 61
rect 36 59 38 61
rect 31 54 38 59
rect 31 52 34 54
rect 36 52 38 54
rect 31 50 38 52
rect 31 42 36 50
<< alu1 >>
rect -2 81 42 82
rect -2 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 42 81
rect -2 68 42 79
rect 2 61 8 63
rect 2 59 4 61
rect 6 59 8 61
rect 2 54 8 59
rect 2 52 4 54
rect 6 52 8 54
rect 2 51 8 52
rect 2 22 6 51
rect 10 42 23 47
rect 10 37 14 42
rect 34 38 38 47
rect 10 35 11 37
rect 13 35 14 37
rect 10 33 14 35
rect 19 37 38 38
rect 19 35 21 37
rect 23 35 38 37
rect 19 34 38 35
rect 25 29 38 30
rect 25 27 31 29
rect 33 27 38 29
rect 25 26 38 27
rect 2 20 23 22
rect 2 18 15 20
rect 17 18 23 20
rect 2 17 23 18
rect 34 17 38 26
rect -2 11 42 12
rect -2 9 4 11
rect 6 9 33 11
rect 35 9 42 11
rect -2 1 42 9
rect -2 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 42 1
rect -2 -2 42 -1
<< ptie >>
rect 0 1 40 3
rect 0 -1 3 1
rect 5 -1 11 1
rect 13 -1 19 1
rect 21 -1 27 1
rect 29 -1 35 1
rect 37 -1 40 1
rect 0 -3 40 -1
<< ntie >>
rect 0 81 40 83
rect 0 79 3 81
rect 5 79 11 81
rect 13 79 19 81
rect 21 79 27 81
rect 29 79 35 81
rect 37 79 40 81
rect 0 77 40 79
<< nmos >>
rect 10 15 12 22
rect 20 10 22 22
rect 27 10 29 22
<< pmos >>
rect 9 42 11 69
rect 19 42 21 69
rect 29 42 31 69
<< polyct1 >>
rect 11 35 13 37
rect 21 35 23 37
rect 31 27 33 29
<< ndifct1 >>
rect 15 18 17 20
rect 4 9 6 11
rect 33 9 35 11
<< ntiect1 >>
rect 3 79 5 81
rect 11 79 13 81
rect 19 79 21 81
rect 27 79 29 81
rect 35 79 37 81
<< ptiect1 >>
rect 3 -1 5 1
rect 11 -1 13 1
rect 19 -1 21 1
rect 27 -1 29 1
rect 35 -1 37 1
<< pdifct0 >>
rect 14 59 16 61
rect 14 52 16 54
rect 24 65 26 67
rect 24 58 26 60
rect 34 59 36 61
rect 34 52 36 54
<< pdifct1 >>
rect 4 59 6 61
rect 4 52 6 54
<< alu0 >>
rect 22 67 28 68
rect 22 65 24 67
rect 26 65 28 67
rect 13 61 17 63
rect 13 59 14 61
rect 16 59 17 61
rect 13 54 17 59
rect 22 60 28 65
rect 22 58 24 60
rect 26 58 28 60
rect 22 57 28 58
rect 33 61 37 63
rect 33 59 34 61
rect 36 59 37 61
rect 33 54 37 59
rect 13 52 14 54
rect 16 52 34 54
rect 36 52 37 54
rect 13 50 37 52
<< labels >>
rlabel alu0 15 56 15 56 6 n1
rlabel alu0 35 56 35 56 6 n1
rlabel alu1 4 40 4 40 6 z
rlabel alu1 12 20 12 20 6 z
rlabel alu1 12 40 12 40 6 b
rlabel alu1 20 6 20 6 6 vss
rlabel alu1 20 20 20 20 6 z
rlabel alu1 28 36 28 36 6 a2
rlabel alu1 28 28 28 28 6 a1
rlabel alu1 20 44 20 44 6 b
rlabel alu1 20 74 20 74 6 vdd
rlabel alu1 36 20 36 20 6 a1
rlabel alu1 36 44 36 44 6 a2
<< end >>
